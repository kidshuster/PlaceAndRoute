magic
tech scmos
timestamp 5.53202
<< polysilicon >>
rect 10 10 11 11 
rect 10 11 11 12 
rect 10 12 11 13 
rect 10 13 11 14 
rect 10 14 11 15 
rect 10 15 11 16 
rect 10 26 11 27 
rect 10 27 11 28 
rect 10 28 11 29 
rect 10 29 11 30 
rect 10 30 11 31 
rect 10 31 11 32 
rect 10 42 11 43 
rect 10 43 11 44 
rect 10 44 11 45 
rect 10 45 11 46 
rect 10 46 11 47 
rect 10 47 11 48 
rect 10 58 11 59 
rect 10 60 11 61 
rect 10 61 11 62 
rect 10 62 11 63 
rect 10 63 11 64 
rect 10 74 11 75 
rect 10 76 11 77 
rect 10 77 11 78 
rect 10 78 11 79 
rect 10 79 11 80 
rect 10 90 11 91 
rect 10 91 11 92 
rect 10 92 11 93 
rect 10 93 11 94 
rect 10 94 11 95 
rect 10 95 11 96 
rect 10 106 11 107 
rect 10 108 11 109 
rect 10 109 11 110 
rect 10 111 11 112 
rect 10 122 11 123 
rect 10 123 11 124 
rect 10 124 11 125 
rect 10 125 11 126 
rect 10 127 11 128 
rect 10 154 11 155 
rect 10 155 11 156 
rect 10 156 11 157 
rect 10 157 11 158 
rect 10 158 11 159 
rect 10 159 11 160 
rect 11 10 12 11 
rect 11 11 12 12 
rect 11 12 12 13 
rect 11 13 12 14 
rect 11 14 12 15 
rect 11 15 12 16 
rect 11 26 12 27 
rect 11 27 12 28 
rect 11 28 12 29 
rect 11 29 12 30 
rect 11 30 12 31 
rect 11 31 12 32 
rect 11 42 12 43 
rect 11 43 12 44 
rect 11 44 12 45 
rect 11 45 12 46 
rect 11 46 12 47 
rect 11 47 12 48 
rect 11 58 12 59 
rect 11 59 12 60 
rect 11 60 12 61 
rect 11 61 12 62 
rect 11 62 12 63 
rect 11 63 12 64 
rect 11 74 12 75 
rect 11 75 12 76 
rect 11 76 12 77 
rect 11 77 12 78 
rect 11 78 12 79 
rect 11 79 12 80 
rect 11 90 12 91 
rect 11 91 12 92 
rect 11 92 12 93 
rect 11 93 12 94 
rect 11 94 12 95 
rect 11 95 12 96 
rect 11 106 12 107 
rect 11 107 12 108 
rect 11 108 12 109 
rect 11 109 12 110 
rect 11 110 12 111 
rect 11 111 12 112 
rect 11 122 12 123 
rect 11 123 12 124 
rect 11 124 12 125 
rect 11 125 12 126 
rect 11 126 12 127 
rect 11 127 12 128 
rect 11 154 12 155 
rect 11 155 12 156 
rect 11 156 12 157 
rect 11 157 12 158 
rect 11 158 12 159 
rect 11 159 12 160 
rect 12 10 13 11 
rect 12 11 13 12 
rect 12 12 13 13 
rect 12 13 13 14 
rect 12 14 13 15 
rect 12 15 13 16 
rect 12 26 13 27 
rect 12 27 13 28 
rect 12 28 13 29 
rect 12 29 13 30 
rect 12 30 13 31 
rect 12 31 13 32 
rect 12 42 13 43 
rect 12 43 13 44 
rect 12 44 13 45 
rect 12 45 13 46 
rect 12 46 13 47 
rect 12 47 13 48 
rect 12 58 13 59 
rect 12 59 13 60 
rect 12 60 13 61 
rect 12 61 13 62 
rect 12 62 13 63 
rect 12 63 13 64 
rect 12 74 13 75 
rect 12 75 13 76 
rect 12 76 13 77 
rect 12 77 13 78 
rect 12 78 13 79 
rect 12 79 13 80 
rect 12 90 13 91 
rect 12 91 13 92 
rect 12 92 13 93 
rect 12 93 13 94 
rect 12 94 13 95 
rect 12 95 13 96 
rect 12 106 13 107 
rect 12 107 13 108 
rect 12 108 13 109 
rect 12 109 13 110 
rect 12 110 13 111 
rect 12 111 13 112 
rect 12 122 13 123 
rect 12 123 13 124 
rect 12 124 13 125 
rect 12 125 13 126 
rect 12 126 13 127 
rect 12 127 13 128 
rect 12 154 13 155 
rect 12 155 13 156 
rect 12 156 13 157 
rect 12 157 13 158 
rect 12 158 13 159 
rect 12 159 13 160 
rect 13 10 14 11 
rect 13 11 14 12 
rect 13 12 14 13 
rect 13 13 14 14 
rect 13 14 14 15 
rect 13 15 14 16 
rect 13 26 14 27 
rect 13 27 14 28 
rect 13 28 14 29 
rect 13 29 14 30 
rect 13 30 14 31 
rect 13 31 14 32 
rect 13 42 14 43 
rect 13 43 14 44 
rect 13 44 14 45 
rect 13 45 14 46 
rect 13 46 14 47 
rect 13 47 14 48 
rect 13 58 14 59 
rect 13 59 14 60 
rect 13 60 14 61 
rect 13 61 14 62 
rect 13 62 14 63 
rect 13 63 14 64 
rect 13 74 14 75 
rect 13 75 14 76 
rect 13 76 14 77 
rect 13 77 14 78 
rect 13 78 14 79 
rect 13 79 14 80 
rect 13 90 14 91 
rect 13 91 14 92 
rect 13 92 14 93 
rect 13 93 14 94 
rect 13 94 14 95 
rect 13 95 14 96 
rect 13 106 14 107 
rect 13 107 14 108 
rect 13 108 14 109 
rect 13 109 14 110 
rect 13 110 14 111 
rect 13 111 14 112 
rect 13 122 14 123 
rect 13 123 14 124 
rect 13 124 14 125 
rect 13 125 14 126 
rect 13 126 14 127 
rect 13 127 14 128 
rect 13 154 14 155 
rect 13 155 14 156 
rect 13 156 14 157 
rect 13 157 14 158 
rect 13 158 14 159 
rect 13 159 14 160 
rect 14 10 15 11 
rect 14 11 15 12 
rect 14 12 15 13 
rect 14 13 15 14 
rect 14 14 15 15 
rect 14 15 15 16 
rect 14 26 15 27 
rect 14 27 15 28 
rect 14 28 15 29 
rect 14 29 15 30 
rect 14 30 15 31 
rect 14 31 15 32 
rect 14 42 15 43 
rect 14 43 15 44 
rect 14 44 15 45 
rect 14 45 15 46 
rect 14 46 15 47 
rect 14 47 15 48 
rect 14 58 15 59 
rect 14 59 15 60 
rect 14 60 15 61 
rect 14 61 15 62 
rect 14 62 15 63 
rect 14 63 15 64 
rect 14 74 15 75 
rect 14 75 15 76 
rect 14 76 15 77 
rect 14 77 15 78 
rect 14 78 15 79 
rect 14 79 15 80 
rect 14 90 15 91 
rect 14 91 15 92 
rect 14 92 15 93 
rect 14 93 15 94 
rect 14 94 15 95 
rect 14 95 15 96 
rect 14 106 15 107 
rect 14 107 15 108 
rect 14 108 15 109 
rect 14 109 15 110 
rect 14 110 15 111 
rect 14 111 15 112 
rect 14 122 15 123 
rect 14 123 15 124 
rect 14 124 15 125 
rect 14 125 15 126 
rect 14 126 15 127 
rect 14 127 15 128 
rect 14 154 15 155 
rect 14 155 15 156 
rect 14 156 15 157 
rect 14 157 15 158 
rect 14 158 15 159 
rect 14 159 15 160 
rect 15 10 16 11 
rect 15 11 16 12 
rect 15 12 16 13 
rect 15 13 16 14 
rect 15 14 16 15 
rect 15 15 16 16 
rect 15 26 16 27 
rect 15 28 16 29 
rect 15 29 16 30 
rect 15 30 16 31 
rect 15 31 16 32 
rect 15 42 16 43 
rect 15 43 16 44 
rect 15 44 16 45 
rect 15 45 16 46 
rect 15 47 16 48 
rect 15 58 16 59 
rect 15 60 16 61 
rect 15 61 16 62 
rect 15 62 16 63 
rect 15 63 16 64 
rect 15 74 16 75 
rect 15 75 16 76 
rect 15 76 16 77 
rect 15 77 16 78 
rect 15 78 16 79 
rect 15 79 16 80 
rect 15 90 16 91 
rect 15 92 16 93 
rect 15 93 16 94 
rect 15 94 16 95 
rect 15 95 16 96 
rect 15 106 16 107 
rect 15 107 16 108 
rect 15 108 16 109 
rect 15 109 16 110 
rect 15 110 16 111 
rect 15 111 16 112 
rect 15 122 16 123 
rect 15 124 16 125 
rect 15 125 16 126 
rect 15 126 16 127 
rect 15 127 16 128 
rect 15 154 16 155 
rect 15 155 16 156 
rect 15 156 16 157 
rect 15 157 16 158 
rect 15 158 16 159 
rect 15 159 16 160 
rect 26 10 27 11 
rect 26 12 27 13 
rect 26 13 27 14 
rect 26 14 27 15 
rect 26 15 27 16 
rect 26 26 27 27 
rect 26 27 27 28 
rect 26 28 27 29 
rect 26 29 27 30 
rect 26 30 27 31 
rect 26 31 27 32 
rect 26 42 27 43 
rect 26 44 27 45 
rect 26 45 27 46 
rect 26 47 27 48 
rect 26 90 27 91 
rect 26 92 27 93 
rect 26 93 27 94 
rect 26 95 27 96 
rect 26 106 27 107 
rect 26 107 27 108 
rect 26 108 27 109 
rect 26 109 27 110 
rect 26 110 27 111 
rect 26 111 27 112 
rect 26 122 27 123 
rect 26 123 27 124 
rect 26 124 27 125 
rect 26 125 27 126 
rect 26 126 27 127 
rect 26 127 27 128 
rect 26 138 27 139 
rect 26 140 27 141 
rect 26 141 27 142 
rect 26 142 27 143 
rect 26 143 27 144 
rect 26 154 27 155 
rect 26 156 27 157 
rect 26 157 27 158 
rect 26 159 27 160 
rect 27 10 28 11 
rect 27 11 28 12 
rect 27 12 28 13 
rect 27 13 28 14 
rect 27 14 28 15 
rect 27 15 28 16 
rect 27 26 28 27 
rect 27 27 28 28 
rect 27 28 28 29 
rect 27 29 28 30 
rect 27 30 28 31 
rect 27 31 28 32 
rect 27 42 28 43 
rect 27 43 28 44 
rect 27 44 28 45 
rect 27 45 28 46 
rect 27 46 28 47 
rect 27 47 28 48 
rect 27 90 28 91 
rect 27 91 28 92 
rect 27 92 28 93 
rect 27 93 28 94 
rect 27 94 28 95 
rect 27 95 28 96 
rect 27 106 28 107 
rect 27 107 28 108 
rect 27 108 28 109 
rect 27 109 28 110 
rect 27 110 28 111 
rect 27 111 28 112 
rect 27 122 28 123 
rect 27 123 28 124 
rect 27 124 28 125 
rect 27 125 28 126 
rect 27 126 28 127 
rect 27 127 28 128 
rect 27 138 28 139 
rect 27 139 28 140 
rect 27 140 28 141 
rect 27 141 28 142 
rect 27 142 28 143 
rect 27 143 28 144 
rect 27 154 28 155 
rect 27 155 28 156 
rect 27 156 28 157 
rect 27 157 28 158 
rect 27 158 28 159 
rect 27 159 28 160 
rect 28 10 29 11 
rect 28 11 29 12 
rect 28 12 29 13 
rect 28 13 29 14 
rect 28 14 29 15 
rect 28 15 29 16 
rect 28 26 29 27 
rect 28 27 29 28 
rect 28 28 29 29 
rect 28 29 29 30 
rect 28 30 29 31 
rect 28 31 29 32 
rect 28 42 29 43 
rect 28 43 29 44 
rect 28 44 29 45 
rect 28 45 29 46 
rect 28 46 29 47 
rect 28 47 29 48 
rect 28 90 29 91 
rect 28 91 29 92 
rect 28 92 29 93 
rect 28 93 29 94 
rect 28 94 29 95 
rect 28 95 29 96 
rect 28 106 29 107 
rect 28 107 29 108 
rect 28 108 29 109 
rect 28 109 29 110 
rect 28 110 29 111 
rect 28 111 29 112 
rect 28 122 29 123 
rect 28 123 29 124 
rect 28 124 29 125 
rect 28 125 29 126 
rect 28 126 29 127 
rect 28 127 29 128 
rect 28 138 29 139 
rect 28 139 29 140 
rect 28 140 29 141 
rect 28 141 29 142 
rect 28 142 29 143 
rect 28 143 29 144 
rect 28 154 29 155 
rect 28 155 29 156 
rect 28 156 29 157 
rect 28 157 29 158 
rect 28 158 29 159 
rect 28 159 29 160 
rect 29 10 30 11 
rect 29 11 30 12 
rect 29 12 30 13 
rect 29 13 30 14 
rect 29 14 30 15 
rect 29 15 30 16 
rect 29 26 30 27 
rect 29 27 30 28 
rect 29 28 30 29 
rect 29 29 30 30 
rect 29 30 30 31 
rect 29 31 30 32 
rect 29 42 30 43 
rect 29 43 30 44 
rect 29 44 30 45 
rect 29 45 30 46 
rect 29 46 30 47 
rect 29 47 30 48 
rect 29 90 30 91 
rect 29 91 30 92 
rect 29 92 30 93 
rect 29 93 30 94 
rect 29 94 30 95 
rect 29 95 30 96 
rect 29 106 30 107 
rect 29 107 30 108 
rect 29 108 30 109 
rect 29 109 30 110 
rect 29 110 30 111 
rect 29 111 30 112 
rect 29 122 30 123 
rect 29 123 30 124 
rect 29 124 30 125 
rect 29 125 30 126 
rect 29 126 30 127 
rect 29 127 30 128 
rect 29 138 30 139 
rect 29 139 30 140 
rect 29 140 30 141 
rect 29 141 30 142 
rect 29 142 30 143 
rect 29 143 30 144 
rect 29 154 30 155 
rect 29 155 30 156 
rect 29 156 30 157 
rect 29 157 30 158 
rect 29 158 30 159 
rect 29 159 30 160 
rect 30 10 31 11 
rect 30 11 31 12 
rect 30 12 31 13 
rect 30 13 31 14 
rect 30 14 31 15 
rect 30 15 31 16 
rect 30 26 31 27 
rect 30 27 31 28 
rect 30 28 31 29 
rect 30 29 31 30 
rect 30 30 31 31 
rect 30 31 31 32 
rect 30 42 31 43 
rect 30 43 31 44 
rect 30 44 31 45 
rect 30 45 31 46 
rect 30 46 31 47 
rect 30 47 31 48 
rect 30 90 31 91 
rect 30 91 31 92 
rect 30 92 31 93 
rect 30 93 31 94 
rect 30 94 31 95 
rect 30 95 31 96 
rect 30 106 31 107 
rect 30 107 31 108 
rect 30 108 31 109 
rect 30 109 31 110 
rect 30 110 31 111 
rect 30 111 31 112 
rect 30 122 31 123 
rect 30 123 31 124 
rect 30 124 31 125 
rect 30 125 31 126 
rect 30 126 31 127 
rect 30 127 31 128 
rect 30 138 31 139 
rect 30 139 31 140 
rect 30 140 31 141 
rect 30 141 31 142 
rect 30 142 31 143 
rect 30 143 31 144 
rect 30 154 31 155 
rect 30 155 31 156 
rect 30 156 31 157 
rect 30 157 31 158 
rect 30 158 31 159 
rect 30 159 31 160 
rect 31 10 32 11 
rect 31 12 32 13 
rect 31 13 32 14 
rect 31 14 32 15 
rect 31 15 32 16 
rect 31 26 32 27 
rect 31 28 32 29 
rect 31 29 32 30 
rect 31 30 32 31 
rect 31 31 32 32 
rect 31 42 32 43 
rect 31 43 32 44 
rect 31 44 32 45 
rect 31 45 32 46 
rect 31 47 32 48 
rect 31 90 32 91 
rect 31 92 32 93 
rect 31 93 32 94 
rect 31 94 32 95 
rect 31 95 32 96 
rect 31 106 32 107 
rect 31 108 32 109 
rect 31 109 32 110 
rect 31 111 32 112 
rect 31 122 32 123 
rect 31 123 32 124 
rect 31 124 32 125 
rect 31 125 32 126 
rect 31 126 32 127 
rect 31 127 32 128 
rect 31 138 32 139 
rect 31 140 32 141 
rect 31 141 32 142 
rect 31 142 32 143 
rect 31 143 32 144 
rect 31 154 32 155 
rect 31 156 32 157 
rect 31 157 32 158 
rect 31 159 32 160 
rect 42 10 43 11 
rect 42 11 43 12 
rect 42 12 43 13 
rect 42 13 43 14 
rect 42 15 43 16 
rect 42 26 43 27 
rect 42 28 43 29 
rect 42 29 43 30 
rect 42 30 43 31 
rect 42 31 43 32 
rect 42 42 43 43 
rect 42 43 43 44 
rect 42 44 43 45 
rect 42 45 43 46 
rect 42 47 43 48 
rect 42 74 43 75 
rect 42 75 43 76 
rect 42 76 43 77 
rect 42 77 43 78 
rect 42 79 43 80 
rect 42 90 43 91 
rect 42 91 43 92 
rect 42 92 43 93 
rect 42 93 43 94 
rect 42 95 43 96 
rect 42 106 43 107 
rect 42 108 43 109 
rect 42 109 43 110 
rect 42 111 43 112 
rect 42 122 43 123 
rect 42 124 43 125 
rect 42 125 43 126 
rect 42 126 43 127 
rect 42 127 43 128 
rect 42 138 43 139 
rect 42 140 43 141 
rect 42 141 43 142 
rect 42 143 43 144 
rect 42 154 43 155 
rect 42 156 43 157 
rect 42 157 43 158 
rect 42 158 43 159 
rect 42 159 43 160 
rect 43 10 44 11 
rect 43 11 44 12 
rect 43 12 44 13 
rect 43 13 44 14 
rect 43 14 44 15 
rect 43 15 44 16 
rect 43 26 44 27 
rect 43 27 44 28 
rect 43 28 44 29 
rect 43 29 44 30 
rect 43 30 44 31 
rect 43 31 44 32 
rect 43 42 44 43 
rect 43 43 44 44 
rect 43 44 44 45 
rect 43 45 44 46 
rect 43 46 44 47 
rect 43 47 44 48 
rect 43 74 44 75 
rect 43 75 44 76 
rect 43 76 44 77 
rect 43 77 44 78 
rect 43 78 44 79 
rect 43 79 44 80 
rect 43 90 44 91 
rect 43 91 44 92 
rect 43 92 44 93 
rect 43 93 44 94 
rect 43 94 44 95 
rect 43 95 44 96 
rect 43 106 44 107 
rect 43 107 44 108 
rect 43 108 44 109 
rect 43 109 44 110 
rect 43 110 44 111 
rect 43 111 44 112 
rect 43 122 44 123 
rect 43 123 44 124 
rect 43 124 44 125 
rect 43 125 44 126 
rect 43 126 44 127 
rect 43 127 44 128 
rect 43 138 44 139 
rect 43 139 44 140 
rect 43 140 44 141 
rect 43 141 44 142 
rect 43 142 44 143 
rect 43 143 44 144 
rect 43 154 44 155 
rect 43 155 44 156 
rect 43 156 44 157 
rect 43 157 44 158 
rect 43 158 44 159 
rect 43 159 44 160 
rect 44 10 45 11 
rect 44 11 45 12 
rect 44 12 45 13 
rect 44 13 45 14 
rect 44 14 45 15 
rect 44 15 45 16 
rect 44 26 45 27 
rect 44 27 45 28 
rect 44 28 45 29 
rect 44 29 45 30 
rect 44 30 45 31 
rect 44 31 45 32 
rect 44 42 45 43 
rect 44 43 45 44 
rect 44 44 45 45 
rect 44 45 45 46 
rect 44 46 45 47 
rect 44 47 45 48 
rect 44 74 45 75 
rect 44 75 45 76 
rect 44 76 45 77 
rect 44 77 45 78 
rect 44 78 45 79 
rect 44 79 45 80 
rect 44 90 45 91 
rect 44 91 45 92 
rect 44 92 45 93 
rect 44 93 45 94 
rect 44 94 45 95 
rect 44 95 45 96 
rect 44 106 45 107 
rect 44 107 45 108 
rect 44 108 45 109 
rect 44 109 45 110 
rect 44 110 45 111 
rect 44 111 45 112 
rect 44 122 45 123 
rect 44 123 45 124 
rect 44 124 45 125 
rect 44 125 45 126 
rect 44 126 45 127 
rect 44 127 45 128 
rect 44 138 45 139 
rect 44 139 45 140 
rect 44 140 45 141 
rect 44 141 45 142 
rect 44 142 45 143 
rect 44 143 45 144 
rect 44 154 45 155 
rect 44 155 45 156 
rect 44 156 45 157 
rect 44 157 45 158 
rect 44 158 45 159 
rect 44 159 45 160 
rect 45 10 46 11 
rect 45 11 46 12 
rect 45 12 46 13 
rect 45 13 46 14 
rect 45 14 46 15 
rect 45 15 46 16 
rect 45 26 46 27 
rect 45 27 46 28 
rect 45 28 46 29 
rect 45 29 46 30 
rect 45 30 46 31 
rect 45 31 46 32 
rect 45 42 46 43 
rect 45 43 46 44 
rect 45 44 46 45 
rect 45 45 46 46 
rect 45 46 46 47 
rect 45 47 46 48 
rect 45 74 46 75 
rect 45 75 46 76 
rect 45 76 46 77 
rect 45 77 46 78 
rect 45 78 46 79 
rect 45 79 46 80 
rect 45 90 46 91 
rect 45 91 46 92 
rect 45 92 46 93 
rect 45 93 46 94 
rect 45 94 46 95 
rect 45 95 46 96 
rect 45 106 46 107 
rect 45 107 46 108 
rect 45 108 46 109 
rect 45 109 46 110 
rect 45 110 46 111 
rect 45 111 46 112 
rect 45 122 46 123 
rect 45 123 46 124 
rect 45 124 46 125 
rect 45 125 46 126 
rect 45 126 46 127 
rect 45 127 46 128 
rect 45 138 46 139 
rect 45 139 46 140 
rect 45 140 46 141 
rect 45 141 46 142 
rect 45 142 46 143 
rect 45 143 46 144 
rect 45 154 46 155 
rect 45 155 46 156 
rect 45 156 46 157 
rect 45 157 46 158 
rect 45 158 46 159 
rect 45 159 46 160 
rect 46 10 47 11 
rect 46 11 47 12 
rect 46 12 47 13 
rect 46 13 47 14 
rect 46 14 47 15 
rect 46 15 47 16 
rect 46 26 47 27 
rect 46 27 47 28 
rect 46 28 47 29 
rect 46 29 47 30 
rect 46 30 47 31 
rect 46 31 47 32 
rect 46 42 47 43 
rect 46 43 47 44 
rect 46 44 47 45 
rect 46 45 47 46 
rect 46 46 47 47 
rect 46 47 47 48 
rect 46 74 47 75 
rect 46 75 47 76 
rect 46 76 47 77 
rect 46 77 47 78 
rect 46 78 47 79 
rect 46 79 47 80 
rect 46 90 47 91 
rect 46 91 47 92 
rect 46 92 47 93 
rect 46 93 47 94 
rect 46 94 47 95 
rect 46 95 47 96 
rect 46 106 47 107 
rect 46 107 47 108 
rect 46 108 47 109 
rect 46 109 47 110 
rect 46 110 47 111 
rect 46 111 47 112 
rect 46 122 47 123 
rect 46 123 47 124 
rect 46 124 47 125 
rect 46 125 47 126 
rect 46 126 47 127 
rect 46 127 47 128 
rect 46 138 47 139 
rect 46 139 47 140 
rect 46 140 47 141 
rect 46 141 47 142 
rect 46 142 47 143 
rect 46 143 47 144 
rect 46 154 47 155 
rect 46 155 47 156 
rect 46 156 47 157 
rect 46 157 47 158 
rect 46 158 47 159 
rect 46 159 47 160 
rect 47 10 48 11 
rect 47 11 48 12 
rect 47 12 48 13 
rect 47 13 48 14 
rect 47 14 48 15 
rect 47 15 48 16 
rect 47 26 48 27 
rect 47 28 48 29 
rect 47 29 48 30 
rect 47 30 48 31 
rect 47 31 48 32 
rect 47 42 48 43 
rect 47 44 48 45 
rect 47 45 48 46 
rect 47 46 48 47 
rect 47 47 48 48 
rect 47 74 48 75 
rect 47 76 48 77 
rect 47 77 48 78 
rect 47 79 48 80 
rect 47 90 48 91 
rect 47 92 48 93 
rect 47 93 48 94 
rect 47 95 48 96 
rect 47 106 48 107 
rect 47 108 48 109 
rect 47 109 48 110 
rect 47 111 48 112 
rect 47 122 48 123 
rect 47 123 48 124 
rect 47 124 48 125 
rect 47 125 48 126 
rect 47 126 48 127 
rect 47 127 48 128 
rect 47 138 48 139 
rect 47 140 48 141 
rect 47 141 48 142 
rect 47 143 48 144 
rect 47 154 48 155 
rect 47 156 48 157 
rect 47 157 48 158 
rect 47 158 48 159 
rect 47 159 48 160 
rect 58 10 59 11 
rect 58 12 59 13 
rect 58 13 59 14 
rect 58 15 59 16 
rect 58 26 59 27 
rect 58 28 59 29 
rect 58 29 59 30 
rect 58 31 59 32 
rect 58 42 59 43 
rect 58 44 59 45 
rect 58 45 59 46 
rect 58 47 59 48 
rect 58 58 59 59 
rect 58 60 59 61 
rect 58 61 59 62 
rect 58 63 59 64 
rect 58 74 59 75 
rect 58 75 59 76 
rect 58 76 59 77 
rect 58 77 59 78 
rect 58 78 59 79 
rect 58 79 59 80 
rect 58 106 59 107 
rect 58 108 59 109 
rect 58 109 59 110 
rect 58 111 59 112 
rect 58 138 59 139 
rect 58 140 59 141 
rect 58 141 59 142 
rect 58 143 59 144 
rect 58 154 59 155 
rect 58 156 59 157 
rect 58 157 59 158 
rect 58 158 59 159 
rect 58 159 59 160 
rect 59 10 60 11 
rect 59 11 60 12 
rect 59 12 60 13 
rect 59 13 60 14 
rect 59 14 60 15 
rect 59 15 60 16 
rect 59 26 60 27 
rect 59 27 60 28 
rect 59 28 60 29 
rect 59 29 60 30 
rect 59 30 60 31 
rect 59 31 60 32 
rect 59 42 60 43 
rect 59 43 60 44 
rect 59 44 60 45 
rect 59 45 60 46 
rect 59 46 60 47 
rect 59 47 60 48 
rect 59 58 60 59 
rect 59 59 60 60 
rect 59 60 60 61 
rect 59 61 60 62 
rect 59 62 60 63 
rect 59 63 60 64 
rect 59 74 60 75 
rect 59 75 60 76 
rect 59 76 60 77 
rect 59 77 60 78 
rect 59 78 60 79 
rect 59 79 60 80 
rect 59 106 60 107 
rect 59 107 60 108 
rect 59 108 60 109 
rect 59 109 60 110 
rect 59 110 60 111 
rect 59 111 60 112 
rect 59 138 60 139 
rect 59 139 60 140 
rect 59 140 60 141 
rect 59 141 60 142 
rect 59 142 60 143 
rect 59 143 60 144 
rect 59 154 60 155 
rect 59 155 60 156 
rect 59 156 60 157 
rect 59 157 60 158 
rect 59 158 60 159 
rect 59 159 60 160 
rect 60 10 61 11 
rect 60 11 61 12 
rect 60 12 61 13 
rect 60 13 61 14 
rect 60 14 61 15 
rect 60 15 61 16 
rect 60 26 61 27 
rect 60 27 61 28 
rect 60 28 61 29 
rect 60 29 61 30 
rect 60 30 61 31 
rect 60 31 61 32 
rect 60 42 61 43 
rect 60 43 61 44 
rect 60 44 61 45 
rect 60 45 61 46 
rect 60 46 61 47 
rect 60 47 61 48 
rect 60 58 61 59 
rect 60 59 61 60 
rect 60 60 61 61 
rect 60 61 61 62 
rect 60 62 61 63 
rect 60 63 61 64 
rect 60 74 61 75 
rect 60 75 61 76 
rect 60 76 61 77 
rect 60 77 61 78 
rect 60 78 61 79 
rect 60 79 61 80 
rect 60 106 61 107 
rect 60 107 61 108 
rect 60 108 61 109 
rect 60 109 61 110 
rect 60 110 61 111 
rect 60 111 61 112 
rect 60 138 61 139 
rect 60 139 61 140 
rect 60 140 61 141 
rect 60 141 61 142 
rect 60 142 61 143 
rect 60 143 61 144 
rect 60 154 61 155 
rect 60 155 61 156 
rect 60 156 61 157 
rect 60 157 61 158 
rect 60 158 61 159 
rect 60 159 61 160 
rect 61 10 62 11 
rect 61 11 62 12 
rect 61 12 62 13 
rect 61 13 62 14 
rect 61 14 62 15 
rect 61 15 62 16 
rect 61 26 62 27 
rect 61 27 62 28 
rect 61 28 62 29 
rect 61 29 62 30 
rect 61 30 62 31 
rect 61 31 62 32 
rect 61 42 62 43 
rect 61 43 62 44 
rect 61 44 62 45 
rect 61 45 62 46 
rect 61 46 62 47 
rect 61 47 62 48 
rect 61 58 62 59 
rect 61 59 62 60 
rect 61 60 62 61 
rect 61 61 62 62 
rect 61 62 62 63 
rect 61 63 62 64 
rect 61 74 62 75 
rect 61 75 62 76 
rect 61 76 62 77 
rect 61 77 62 78 
rect 61 78 62 79 
rect 61 79 62 80 
rect 61 106 62 107 
rect 61 107 62 108 
rect 61 108 62 109 
rect 61 109 62 110 
rect 61 110 62 111 
rect 61 111 62 112 
rect 61 138 62 139 
rect 61 139 62 140 
rect 61 140 62 141 
rect 61 141 62 142 
rect 61 142 62 143 
rect 61 143 62 144 
rect 61 154 62 155 
rect 61 155 62 156 
rect 61 156 62 157 
rect 61 157 62 158 
rect 61 158 62 159 
rect 61 159 62 160 
rect 62 10 63 11 
rect 62 11 63 12 
rect 62 12 63 13 
rect 62 13 63 14 
rect 62 14 63 15 
rect 62 15 63 16 
rect 62 26 63 27 
rect 62 27 63 28 
rect 62 28 63 29 
rect 62 29 63 30 
rect 62 30 63 31 
rect 62 31 63 32 
rect 62 42 63 43 
rect 62 43 63 44 
rect 62 44 63 45 
rect 62 45 63 46 
rect 62 46 63 47 
rect 62 47 63 48 
rect 62 58 63 59 
rect 62 59 63 60 
rect 62 60 63 61 
rect 62 61 63 62 
rect 62 62 63 63 
rect 62 63 63 64 
rect 62 74 63 75 
rect 62 75 63 76 
rect 62 76 63 77 
rect 62 77 63 78 
rect 62 78 63 79 
rect 62 79 63 80 
rect 62 106 63 107 
rect 62 107 63 108 
rect 62 108 63 109 
rect 62 109 63 110 
rect 62 110 63 111 
rect 62 111 63 112 
rect 62 138 63 139 
rect 62 139 63 140 
rect 62 140 63 141 
rect 62 141 63 142 
rect 62 142 63 143 
rect 62 143 63 144 
rect 62 154 63 155 
rect 62 155 63 156 
rect 62 156 63 157 
rect 62 157 63 158 
rect 62 158 63 159 
rect 62 159 63 160 
rect 63 10 64 11 
rect 63 12 64 13 
rect 63 13 64 14 
rect 63 14 64 15 
rect 63 15 64 16 
rect 63 26 64 27 
rect 63 28 64 29 
rect 63 29 64 30 
rect 63 31 64 32 
rect 63 42 64 43 
rect 63 44 64 45 
rect 63 45 64 46 
rect 63 46 64 47 
rect 63 47 64 48 
rect 63 58 64 59 
rect 63 60 64 61 
rect 63 61 64 62 
rect 63 63 64 64 
rect 63 74 64 75 
rect 63 75 64 76 
rect 63 76 64 77 
rect 63 77 64 78 
rect 63 79 64 80 
rect 63 106 64 107 
rect 63 108 64 109 
rect 63 109 64 110 
rect 63 110 64 111 
rect 63 111 64 112 
rect 63 138 64 139 
rect 63 139 64 140 
rect 63 140 64 141 
rect 63 141 64 142 
rect 63 143 64 144 
rect 63 154 64 155 
rect 63 155 64 156 
rect 63 156 64 157 
rect 63 157 64 158 
rect 63 159 64 160 
rect 74 10 75 11 
rect 74 12 75 13 
rect 74 13 75 14 
rect 74 15 75 16 
rect 74 42 75 43 
rect 74 43 75 44 
rect 74 44 75 45 
rect 74 45 75 46 
rect 74 47 75 48 
rect 74 58 75 59 
rect 74 59 75 60 
rect 74 60 75 61 
rect 74 61 75 62 
rect 74 63 75 64 
rect 74 74 75 75 
rect 74 76 75 77 
rect 74 77 75 78 
rect 74 79 75 80 
rect 74 90 75 91 
rect 74 92 75 93 
rect 74 93 75 94 
rect 74 95 75 96 
rect 74 106 75 107 
rect 74 107 75 108 
rect 74 108 75 109 
rect 74 109 75 110 
rect 74 110 75 111 
rect 74 111 75 112 
rect 74 138 75 139 
rect 74 139 75 140 
rect 74 140 75 141 
rect 74 141 75 142 
rect 74 143 75 144 
rect 75 10 76 11 
rect 75 11 76 12 
rect 75 12 76 13 
rect 75 13 76 14 
rect 75 14 76 15 
rect 75 15 76 16 
rect 75 42 76 43 
rect 75 43 76 44 
rect 75 44 76 45 
rect 75 45 76 46 
rect 75 46 76 47 
rect 75 47 76 48 
rect 75 58 76 59 
rect 75 59 76 60 
rect 75 60 76 61 
rect 75 61 76 62 
rect 75 62 76 63 
rect 75 63 76 64 
rect 75 74 76 75 
rect 75 75 76 76 
rect 75 76 76 77 
rect 75 77 76 78 
rect 75 78 76 79 
rect 75 79 76 80 
rect 75 90 76 91 
rect 75 91 76 92 
rect 75 92 76 93 
rect 75 93 76 94 
rect 75 94 76 95 
rect 75 95 76 96 
rect 75 106 76 107 
rect 75 107 76 108 
rect 75 108 76 109 
rect 75 109 76 110 
rect 75 110 76 111 
rect 75 111 76 112 
rect 75 138 76 139 
rect 75 139 76 140 
rect 75 140 76 141 
rect 75 141 76 142 
rect 75 142 76 143 
rect 75 143 76 144 
rect 76 10 77 11 
rect 76 11 77 12 
rect 76 12 77 13 
rect 76 13 77 14 
rect 76 14 77 15 
rect 76 15 77 16 
rect 76 42 77 43 
rect 76 43 77 44 
rect 76 44 77 45 
rect 76 45 77 46 
rect 76 46 77 47 
rect 76 47 77 48 
rect 76 58 77 59 
rect 76 59 77 60 
rect 76 60 77 61 
rect 76 61 77 62 
rect 76 62 77 63 
rect 76 63 77 64 
rect 76 74 77 75 
rect 76 75 77 76 
rect 76 76 77 77 
rect 76 77 77 78 
rect 76 78 77 79 
rect 76 79 77 80 
rect 76 90 77 91 
rect 76 91 77 92 
rect 76 92 77 93 
rect 76 93 77 94 
rect 76 94 77 95 
rect 76 95 77 96 
rect 76 106 77 107 
rect 76 107 77 108 
rect 76 108 77 109 
rect 76 109 77 110 
rect 76 110 77 111 
rect 76 111 77 112 
rect 76 138 77 139 
rect 76 139 77 140 
rect 76 140 77 141 
rect 76 141 77 142 
rect 76 142 77 143 
rect 76 143 77 144 
rect 77 10 78 11 
rect 77 11 78 12 
rect 77 12 78 13 
rect 77 13 78 14 
rect 77 14 78 15 
rect 77 15 78 16 
rect 77 42 78 43 
rect 77 43 78 44 
rect 77 44 78 45 
rect 77 45 78 46 
rect 77 46 78 47 
rect 77 47 78 48 
rect 77 58 78 59 
rect 77 59 78 60 
rect 77 60 78 61 
rect 77 61 78 62 
rect 77 62 78 63 
rect 77 63 78 64 
rect 77 74 78 75 
rect 77 75 78 76 
rect 77 76 78 77 
rect 77 77 78 78 
rect 77 78 78 79 
rect 77 79 78 80 
rect 77 90 78 91 
rect 77 91 78 92 
rect 77 92 78 93 
rect 77 93 78 94 
rect 77 94 78 95 
rect 77 95 78 96 
rect 77 106 78 107 
rect 77 107 78 108 
rect 77 108 78 109 
rect 77 109 78 110 
rect 77 110 78 111 
rect 77 111 78 112 
rect 77 138 78 139 
rect 77 139 78 140 
rect 77 140 78 141 
rect 77 141 78 142 
rect 77 142 78 143 
rect 77 143 78 144 
rect 78 10 79 11 
rect 78 11 79 12 
rect 78 12 79 13 
rect 78 13 79 14 
rect 78 14 79 15 
rect 78 15 79 16 
rect 78 42 79 43 
rect 78 43 79 44 
rect 78 44 79 45 
rect 78 45 79 46 
rect 78 46 79 47 
rect 78 47 79 48 
rect 78 58 79 59 
rect 78 59 79 60 
rect 78 60 79 61 
rect 78 61 79 62 
rect 78 62 79 63 
rect 78 63 79 64 
rect 78 74 79 75 
rect 78 75 79 76 
rect 78 76 79 77 
rect 78 77 79 78 
rect 78 78 79 79 
rect 78 79 79 80 
rect 78 90 79 91 
rect 78 91 79 92 
rect 78 92 79 93 
rect 78 93 79 94 
rect 78 94 79 95 
rect 78 95 79 96 
rect 78 106 79 107 
rect 78 107 79 108 
rect 78 108 79 109 
rect 78 109 79 110 
rect 78 110 79 111 
rect 78 111 79 112 
rect 78 138 79 139 
rect 78 139 79 140 
rect 78 140 79 141 
rect 78 141 79 142 
rect 78 142 79 143 
rect 78 143 79 144 
rect 79 10 80 11 
rect 79 11 80 12 
rect 79 12 80 13 
rect 79 13 80 14 
rect 79 14 80 15 
rect 79 15 80 16 
rect 79 42 80 43 
rect 79 44 80 45 
rect 79 45 80 46 
rect 79 46 80 47 
rect 79 47 80 48 
rect 79 58 80 59 
rect 79 59 80 60 
rect 79 60 80 61 
rect 79 61 80 62 
rect 79 62 80 63 
rect 79 63 80 64 
rect 79 74 80 75 
rect 79 76 80 77 
rect 79 77 80 78 
rect 79 79 80 80 
rect 79 90 80 91 
rect 79 91 80 92 
rect 79 92 80 93 
rect 79 93 80 94 
rect 79 95 80 96 
rect 79 106 80 107 
rect 79 107 80 108 
rect 79 108 80 109 
rect 79 109 80 110 
rect 79 111 80 112 
rect 79 138 80 139 
rect 79 140 80 141 
rect 79 141 80 142 
rect 79 142 80 143 
rect 79 143 80 144 
rect 90 10 91 11 
rect 90 11 91 12 
rect 90 12 91 13 
rect 90 13 91 14 
rect 90 14 91 15 
rect 90 15 91 16 
rect 90 26 91 27 
rect 90 28 91 29 
rect 90 29 91 30 
rect 90 30 91 31 
rect 90 31 91 32 
rect 90 42 91 43 
rect 90 43 91 44 
rect 90 44 91 45 
rect 90 45 91 46 
rect 90 47 91 48 
rect 90 58 91 59 
rect 90 60 91 61 
rect 90 61 91 62 
rect 90 62 91 63 
rect 90 63 91 64 
rect 90 90 91 91 
rect 90 91 91 92 
rect 90 92 91 93 
rect 90 93 91 94 
rect 90 94 91 95 
rect 90 95 91 96 
rect 90 122 91 123 
rect 90 124 91 125 
rect 90 125 91 126 
rect 90 127 91 128 
rect 90 138 91 139 
rect 90 140 91 141 
rect 90 141 91 142 
rect 90 143 91 144 
rect 90 154 91 155 
rect 90 156 91 157 
rect 90 157 91 158 
rect 90 159 91 160 
rect 91 10 92 11 
rect 91 11 92 12 
rect 91 12 92 13 
rect 91 13 92 14 
rect 91 14 92 15 
rect 91 15 92 16 
rect 91 26 92 27 
rect 91 27 92 28 
rect 91 28 92 29 
rect 91 29 92 30 
rect 91 30 92 31 
rect 91 31 92 32 
rect 91 42 92 43 
rect 91 43 92 44 
rect 91 44 92 45 
rect 91 45 92 46 
rect 91 46 92 47 
rect 91 47 92 48 
rect 91 58 92 59 
rect 91 59 92 60 
rect 91 60 92 61 
rect 91 61 92 62 
rect 91 62 92 63 
rect 91 63 92 64 
rect 91 90 92 91 
rect 91 91 92 92 
rect 91 92 92 93 
rect 91 93 92 94 
rect 91 94 92 95 
rect 91 95 92 96 
rect 91 122 92 123 
rect 91 123 92 124 
rect 91 124 92 125 
rect 91 125 92 126 
rect 91 126 92 127 
rect 91 127 92 128 
rect 91 138 92 139 
rect 91 139 92 140 
rect 91 140 92 141 
rect 91 141 92 142 
rect 91 142 92 143 
rect 91 143 92 144 
rect 91 154 92 155 
rect 91 155 92 156 
rect 91 156 92 157 
rect 91 157 92 158 
rect 91 158 92 159 
rect 91 159 92 160 
rect 92 10 93 11 
rect 92 11 93 12 
rect 92 12 93 13 
rect 92 13 93 14 
rect 92 14 93 15 
rect 92 15 93 16 
rect 92 26 93 27 
rect 92 27 93 28 
rect 92 28 93 29 
rect 92 29 93 30 
rect 92 30 93 31 
rect 92 31 93 32 
rect 92 42 93 43 
rect 92 43 93 44 
rect 92 44 93 45 
rect 92 45 93 46 
rect 92 46 93 47 
rect 92 47 93 48 
rect 92 58 93 59 
rect 92 59 93 60 
rect 92 60 93 61 
rect 92 61 93 62 
rect 92 62 93 63 
rect 92 63 93 64 
rect 92 90 93 91 
rect 92 91 93 92 
rect 92 92 93 93 
rect 92 93 93 94 
rect 92 94 93 95 
rect 92 95 93 96 
rect 92 122 93 123 
rect 92 123 93 124 
rect 92 124 93 125 
rect 92 125 93 126 
rect 92 126 93 127 
rect 92 127 93 128 
rect 92 138 93 139 
rect 92 139 93 140 
rect 92 140 93 141 
rect 92 141 93 142 
rect 92 142 93 143 
rect 92 143 93 144 
rect 92 154 93 155 
rect 92 155 93 156 
rect 92 156 93 157 
rect 92 157 93 158 
rect 92 158 93 159 
rect 92 159 93 160 
rect 93 10 94 11 
rect 93 11 94 12 
rect 93 12 94 13 
rect 93 13 94 14 
rect 93 14 94 15 
rect 93 15 94 16 
rect 93 26 94 27 
rect 93 27 94 28 
rect 93 28 94 29 
rect 93 29 94 30 
rect 93 30 94 31 
rect 93 31 94 32 
rect 93 42 94 43 
rect 93 43 94 44 
rect 93 44 94 45 
rect 93 45 94 46 
rect 93 46 94 47 
rect 93 47 94 48 
rect 93 58 94 59 
rect 93 59 94 60 
rect 93 60 94 61 
rect 93 61 94 62 
rect 93 62 94 63 
rect 93 63 94 64 
rect 93 90 94 91 
rect 93 91 94 92 
rect 93 92 94 93 
rect 93 93 94 94 
rect 93 94 94 95 
rect 93 95 94 96 
rect 93 122 94 123 
rect 93 123 94 124 
rect 93 124 94 125 
rect 93 125 94 126 
rect 93 126 94 127 
rect 93 127 94 128 
rect 93 138 94 139 
rect 93 139 94 140 
rect 93 140 94 141 
rect 93 141 94 142 
rect 93 142 94 143 
rect 93 143 94 144 
rect 93 154 94 155 
rect 93 155 94 156 
rect 93 156 94 157 
rect 93 157 94 158 
rect 93 158 94 159 
rect 93 159 94 160 
rect 94 10 95 11 
rect 94 11 95 12 
rect 94 12 95 13 
rect 94 13 95 14 
rect 94 14 95 15 
rect 94 15 95 16 
rect 94 26 95 27 
rect 94 27 95 28 
rect 94 28 95 29 
rect 94 29 95 30 
rect 94 30 95 31 
rect 94 31 95 32 
rect 94 42 95 43 
rect 94 43 95 44 
rect 94 44 95 45 
rect 94 45 95 46 
rect 94 46 95 47 
rect 94 47 95 48 
rect 94 58 95 59 
rect 94 59 95 60 
rect 94 60 95 61 
rect 94 61 95 62 
rect 94 62 95 63 
rect 94 63 95 64 
rect 94 90 95 91 
rect 94 91 95 92 
rect 94 92 95 93 
rect 94 93 95 94 
rect 94 94 95 95 
rect 94 95 95 96 
rect 94 122 95 123 
rect 94 123 95 124 
rect 94 124 95 125 
rect 94 125 95 126 
rect 94 126 95 127 
rect 94 127 95 128 
rect 94 138 95 139 
rect 94 139 95 140 
rect 94 140 95 141 
rect 94 141 95 142 
rect 94 142 95 143 
rect 94 143 95 144 
rect 94 154 95 155 
rect 94 155 95 156 
rect 94 156 95 157 
rect 94 157 95 158 
rect 94 158 95 159 
rect 94 159 95 160 
rect 95 10 96 11 
rect 95 11 96 12 
rect 95 12 96 13 
rect 95 13 96 14 
rect 95 14 96 15 
rect 95 15 96 16 
rect 95 26 96 27 
rect 95 28 96 29 
rect 95 29 96 30 
rect 95 31 96 32 
rect 95 42 96 43 
rect 95 43 96 44 
rect 95 44 96 45 
rect 95 45 96 46 
rect 95 47 96 48 
rect 95 58 96 59 
rect 95 59 96 60 
rect 95 60 96 61 
rect 95 61 96 62 
rect 95 63 96 64 
rect 95 90 96 91 
rect 95 91 96 92 
rect 95 92 96 93 
rect 95 93 96 94 
rect 95 94 96 95 
rect 95 95 96 96 
rect 95 122 96 123 
rect 95 123 96 124 
rect 95 124 96 125 
rect 95 125 96 126 
rect 95 126 96 127 
rect 95 127 96 128 
rect 95 138 96 139 
rect 95 139 96 140 
rect 95 140 96 141 
rect 95 141 96 142 
rect 95 143 96 144 
rect 95 154 96 155 
rect 95 156 96 157 
rect 95 157 96 158 
rect 95 158 96 159 
rect 95 159 96 160 
rect 106 10 107 11 
rect 106 11 107 12 
rect 106 12 107 13 
rect 106 13 107 14 
rect 106 14 107 15 
rect 106 15 107 16 
rect 106 58 107 59 
rect 106 59 107 60 
rect 106 60 107 61 
rect 106 61 107 62 
rect 106 63 107 64 
rect 106 74 107 75 
rect 106 75 107 76 
rect 106 76 107 77 
rect 106 77 107 78 
rect 106 79 107 80 
rect 106 90 107 91 
rect 106 91 107 92 
rect 106 92 107 93 
rect 106 93 107 94 
rect 106 94 107 95 
rect 106 95 107 96 
rect 106 106 107 107 
rect 106 107 107 108 
rect 106 108 107 109 
rect 106 109 107 110 
rect 106 111 107 112 
rect 106 122 107 123 
rect 106 124 107 125 
rect 106 125 107 126 
rect 106 127 107 128 
rect 106 138 107 139 
rect 106 140 107 141 
rect 106 141 107 142 
rect 106 142 107 143 
rect 106 143 107 144 
rect 107 10 108 11 
rect 107 11 108 12 
rect 107 12 108 13 
rect 107 13 108 14 
rect 107 14 108 15 
rect 107 15 108 16 
rect 107 58 108 59 
rect 107 59 108 60 
rect 107 60 108 61 
rect 107 61 108 62 
rect 107 62 108 63 
rect 107 63 108 64 
rect 107 74 108 75 
rect 107 75 108 76 
rect 107 76 108 77 
rect 107 77 108 78 
rect 107 78 108 79 
rect 107 79 108 80 
rect 107 90 108 91 
rect 107 91 108 92 
rect 107 92 108 93 
rect 107 93 108 94 
rect 107 94 108 95 
rect 107 95 108 96 
rect 107 106 108 107 
rect 107 107 108 108 
rect 107 108 108 109 
rect 107 109 108 110 
rect 107 110 108 111 
rect 107 111 108 112 
rect 107 122 108 123 
rect 107 123 108 124 
rect 107 124 108 125 
rect 107 125 108 126 
rect 107 126 108 127 
rect 107 127 108 128 
rect 107 138 108 139 
rect 107 139 108 140 
rect 107 140 108 141 
rect 107 141 108 142 
rect 107 142 108 143 
rect 107 143 108 144 
rect 108 10 109 11 
rect 108 11 109 12 
rect 108 12 109 13 
rect 108 13 109 14 
rect 108 14 109 15 
rect 108 15 109 16 
rect 108 58 109 59 
rect 108 59 109 60 
rect 108 60 109 61 
rect 108 61 109 62 
rect 108 62 109 63 
rect 108 63 109 64 
rect 108 74 109 75 
rect 108 75 109 76 
rect 108 76 109 77 
rect 108 77 109 78 
rect 108 78 109 79 
rect 108 79 109 80 
rect 108 90 109 91 
rect 108 91 109 92 
rect 108 92 109 93 
rect 108 93 109 94 
rect 108 94 109 95 
rect 108 95 109 96 
rect 108 106 109 107 
rect 108 107 109 108 
rect 108 108 109 109 
rect 108 109 109 110 
rect 108 110 109 111 
rect 108 111 109 112 
rect 108 122 109 123 
rect 108 123 109 124 
rect 108 124 109 125 
rect 108 125 109 126 
rect 108 126 109 127 
rect 108 127 109 128 
rect 108 138 109 139 
rect 108 139 109 140 
rect 108 140 109 141 
rect 108 141 109 142 
rect 108 142 109 143 
rect 108 143 109 144 
rect 109 10 110 11 
rect 109 11 110 12 
rect 109 12 110 13 
rect 109 13 110 14 
rect 109 14 110 15 
rect 109 15 110 16 
rect 109 58 110 59 
rect 109 59 110 60 
rect 109 60 110 61 
rect 109 61 110 62 
rect 109 62 110 63 
rect 109 63 110 64 
rect 109 74 110 75 
rect 109 75 110 76 
rect 109 76 110 77 
rect 109 77 110 78 
rect 109 78 110 79 
rect 109 79 110 80 
rect 109 90 110 91 
rect 109 91 110 92 
rect 109 92 110 93 
rect 109 93 110 94 
rect 109 94 110 95 
rect 109 95 110 96 
rect 109 106 110 107 
rect 109 107 110 108 
rect 109 108 110 109 
rect 109 109 110 110 
rect 109 110 110 111 
rect 109 111 110 112 
rect 109 122 110 123 
rect 109 123 110 124 
rect 109 124 110 125 
rect 109 125 110 126 
rect 109 126 110 127 
rect 109 127 110 128 
rect 109 138 110 139 
rect 109 139 110 140 
rect 109 140 110 141 
rect 109 141 110 142 
rect 109 142 110 143 
rect 109 143 110 144 
rect 110 10 111 11 
rect 110 11 111 12 
rect 110 12 111 13 
rect 110 13 111 14 
rect 110 14 111 15 
rect 110 15 111 16 
rect 110 58 111 59 
rect 110 59 111 60 
rect 110 60 111 61 
rect 110 61 111 62 
rect 110 62 111 63 
rect 110 63 111 64 
rect 110 74 111 75 
rect 110 75 111 76 
rect 110 76 111 77 
rect 110 77 111 78 
rect 110 78 111 79 
rect 110 79 111 80 
rect 110 90 111 91 
rect 110 91 111 92 
rect 110 92 111 93 
rect 110 93 111 94 
rect 110 94 111 95 
rect 110 95 111 96 
rect 110 106 111 107 
rect 110 107 111 108 
rect 110 108 111 109 
rect 110 109 111 110 
rect 110 110 111 111 
rect 110 111 111 112 
rect 110 122 111 123 
rect 110 123 111 124 
rect 110 124 111 125 
rect 110 125 111 126 
rect 110 126 111 127 
rect 110 127 111 128 
rect 110 138 111 139 
rect 110 139 111 140 
rect 110 140 111 141 
rect 110 141 111 142 
rect 110 142 111 143 
rect 110 143 111 144 
rect 111 10 112 11 
rect 111 12 112 13 
rect 111 13 112 14 
rect 111 14 112 15 
rect 111 15 112 16 
rect 111 58 112 59 
rect 111 59 112 60 
rect 111 60 112 61 
rect 111 61 112 62 
rect 111 62 112 63 
rect 111 63 112 64 
rect 111 74 112 75 
rect 111 75 112 76 
rect 111 76 112 77 
rect 111 77 112 78 
rect 111 78 112 79 
rect 111 79 112 80 
rect 111 90 112 91 
rect 111 91 112 92 
rect 111 92 112 93 
rect 111 93 112 94 
rect 111 94 112 95 
rect 111 95 112 96 
rect 111 106 112 107 
rect 111 108 112 109 
rect 111 109 112 110 
rect 111 110 112 111 
rect 111 111 112 112 
rect 111 122 112 123 
rect 111 124 112 125 
rect 111 125 112 126 
rect 111 127 112 128 
rect 111 138 112 139 
rect 111 139 112 140 
rect 111 140 112 141 
rect 111 141 112 142 
rect 111 142 112 143 
rect 111 143 112 144 
rect 122 10 123 11 
rect 122 11 123 12 
rect 122 12 123 13 
rect 122 13 123 14 
rect 122 14 123 15 
rect 122 15 123 16 
rect 122 26 123 27 
rect 122 27 123 28 
rect 122 28 123 29 
rect 122 29 123 30 
rect 122 31 123 32 
rect 122 42 123 43 
rect 122 43 123 44 
rect 122 44 123 45 
rect 122 45 123 46 
rect 122 46 123 47 
rect 122 47 123 48 
rect 122 58 123 59 
rect 122 60 123 61 
rect 122 61 123 62 
rect 122 63 123 64 
rect 122 74 123 75 
rect 122 75 123 76 
rect 122 76 123 77 
rect 122 77 123 78 
rect 122 79 123 80 
rect 122 90 123 91 
rect 122 92 123 93 
rect 122 93 123 94 
rect 122 94 123 95 
rect 122 95 123 96 
rect 122 122 123 123 
rect 122 124 123 125 
rect 122 125 123 126 
rect 122 126 123 127 
rect 122 127 123 128 
rect 122 154 123 155 
rect 122 156 123 157 
rect 122 157 123 158 
rect 122 158 123 159 
rect 122 159 123 160 
rect 123 10 124 11 
rect 123 11 124 12 
rect 123 12 124 13 
rect 123 13 124 14 
rect 123 14 124 15 
rect 123 15 124 16 
rect 123 26 124 27 
rect 123 27 124 28 
rect 123 28 124 29 
rect 123 29 124 30 
rect 123 30 124 31 
rect 123 31 124 32 
rect 123 42 124 43 
rect 123 43 124 44 
rect 123 44 124 45 
rect 123 45 124 46 
rect 123 46 124 47 
rect 123 47 124 48 
rect 123 58 124 59 
rect 123 59 124 60 
rect 123 60 124 61 
rect 123 61 124 62 
rect 123 62 124 63 
rect 123 63 124 64 
rect 123 74 124 75 
rect 123 75 124 76 
rect 123 76 124 77 
rect 123 77 124 78 
rect 123 78 124 79 
rect 123 79 124 80 
rect 123 90 124 91 
rect 123 91 124 92 
rect 123 92 124 93 
rect 123 93 124 94 
rect 123 94 124 95 
rect 123 95 124 96 
rect 123 122 124 123 
rect 123 123 124 124 
rect 123 124 124 125 
rect 123 125 124 126 
rect 123 126 124 127 
rect 123 127 124 128 
rect 123 154 124 155 
rect 123 155 124 156 
rect 123 156 124 157 
rect 123 157 124 158 
rect 123 158 124 159 
rect 123 159 124 160 
rect 124 10 125 11 
rect 124 11 125 12 
rect 124 12 125 13 
rect 124 13 125 14 
rect 124 14 125 15 
rect 124 15 125 16 
rect 124 26 125 27 
rect 124 27 125 28 
rect 124 28 125 29 
rect 124 29 125 30 
rect 124 30 125 31 
rect 124 31 125 32 
rect 124 42 125 43 
rect 124 43 125 44 
rect 124 44 125 45 
rect 124 45 125 46 
rect 124 46 125 47 
rect 124 47 125 48 
rect 124 58 125 59 
rect 124 59 125 60 
rect 124 60 125 61 
rect 124 61 125 62 
rect 124 62 125 63 
rect 124 63 125 64 
rect 124 74 125 75 
rect 124 75 125 76 
rect 124 76 125 77 
rect 124 77 125 78 
rect 124 78 125 79 
rect 124 79 125 80 
rect 124 90 125 91 
rect 124 91 125 92 
rect 124 92 125 93 
rect 124 93 125 94 
rect 124 94 125 95 
rect 124 95 125 96 
rect 124 122 125 123 
rect 124 123 125 124 
rect 124 124 125 125 
rect 124 125 125 126 
rect 124 126 125 127 
rect 124 127 125 128 
rect 124 154 125 155 
rect 124 155 125 156 
rect 124 156 125 157 
rect 124 157 125 158 
rect 124 158 125 159 
rect 124 159 125 160 
rect 125 10 126 11 
rect 125 11 126 12 
rect 125 12 126 13 
rect 125 13 126 14 
rect 125 14 126 15 
rect 125 15 126 16 
rect 125 26 126 27 
rect 125 27 126 28 
rect 125 28 126 29 
rect 125 29 126 30 
rect 125 30 126 31 
rect 125 31 126 32 
rect 125 42 126 43 
rect 125 43 126 44 
rect 125 44 126 45 
rect 125 45 126 46 
rect 125 46 126 47 
rect 125 47 126 48 
rect 125 58 126 59 
rect 125 59 126 60 
rect 125 60 126 61 
rect 125 61 126 62 
rect 125 62 126 63 
rect 125 63 126 64 
rect 125 74 126 75 
rect 125 75 126 76 
rect 125 76 126 77 
rect 125 77 126 78 
rect 125 78 126 79 
rect 125 79 126 80 
rect 125 90 126 91 
rect 125 91 126 92 
rect 125 92 126 93 
rect 125 93 126 94 
rect 125 94 126 95 
rect 125 95 126 96 
rect 125 122 126 123 
rect 125 123 126 124 
rect 125 124 126 125 
rect 125 125 126 126 
rect 125 126 126 127 
rect 125 127 126 128 
rect 125 154 126 155 
rect 125 155 126 156 
rect 125 156 126 157 
rect 125 157 126 158 
rect 125 158 126 159 
rect 125 159 126 160 
rect 126 10 127 11 
rect 126 11 127 12 
rect 126 12 127 13 
rect 126 13 127 14 
rect 126 14 127 15 
rect 126 15 127 16 
rect 126 26 127 27 
rect 126 27 127 28 
rect 126 28 127 29 
rect 126 29 127 30 
rect 126 30 127 31 
rect 126 31 127 32 
rect 126 42 127 43 
rect 126 43 127 44 
rect 126 44 127 45 
rect 126 45 127 46 
rect 126 46 127 47 
rect 126 47 127 48 
rect 126 58 127 59 
rect 126 59 127 60 
rect 126 60 127 61 
rect 126 61 127 62 
rect 126 62 127 63 
rect 126 63 127 64 
rect 126 74 127 75 
rect 126 75 127 76 
rect 126 76 127 77 
rect 126 77 127 78 
rect 126 78 127 79 
rect 126 79 127 80 
rect 126 90 127 91 
rect 126 91 127 92 
rect 126 92 127 93 
rect 126 93 127 94 
rect 126 94 127 95 
rect 126 95 127 96 
rect 126 122 127 123 
rect 126 123 127 124 
rect 126 124 127 125 
rect 126 125 127 126 
rect 126 126 127 127 
rect 126 127 127 128 
rect 126 154 127 155 
rect 126 155 127 156 
rect 126 156 127 157 
rect 126 157 127 158 
rect 126 158 127 159 
rect 126 159 127 160 
rect 127 10 128 11 
rect 127 12 128 13 
rect 127 13 128 14 
rect 127 14 128 15 
rect 127 15 128 16 
rect 127 26 128 27 
rect 127 27 128 28 
rect 127 28 128 29 
rect 127 29 128 30 
rect 127 30 128 31 
rect 127 31 128 32 
rect 127 42 128 43 
rect 127 44 128 45 
rect 127 45 128 46 
rect 127 46 128 47 
rect 127 47 128 48 
rect 127 58 128 59 
rect 127 59 128 60 
rect 127 60 128 61 
rect 127 61 128 62 
rect 127 63 128 64 
rect 127 74 128 75 
rect 127 76 128 77 
rect 127 77 128 78 
rect 127 79 128 80 
rect 127 90 128 91 
rect 127 92 128 93 
rect 127 93 128 94 
rect 127 95 128 96 
rect 127 122 128 123 
rect 127 123 128 124 
rect 127 124 128 125 
rect 127 125 128 126 
rect 127 127 128 128 
rect 127 154 128 155 
rect 127 155 128 156 
rect 127 156 128 157 
rect 127 157 128 158 
rect 127 158 128 159 
rect 127 159 128 160 
rect 138 10 139 11 
rect 138 11 139 12 
rect 138 12 139 13 
rect 138 13 139 14 
rect 138 14 139 15 
rect 138 15 139 16 
rect 138 42 139 43 
rect 138 43 139 44 
rect 138 44 139 45 
rect 138 45 139 46 
rect 138 47 139 48 
rect 138 90 139 91 
rect 138 92 139 93 
rect 138 93 139 94 
rect 138 94 139 95 
rect 138 95 139 96 
rect 138 106 139 107 
rect 138 107 139 108 
rect 138 108 139 109 
rect 138 109 139 110 
rect 138 111 139 112 
rect 138 122 139 123 
rect 138 124 139 125 
rect 138 125 139 126 
rect 138 126 139 127 
rect 138 127 139 128 
rect 138 138 139 139 
rect 138 140 139 141 
rect 138 141 139 142 
rect 138 143 139 144 
rect 139 10 140 11 
rect 139 11 140 12 
rect 139 12 140 13 
rect 139 13 140 14 
rect 139 14 140 15 
rect 139 15 140 16 
rect 139 42 140 43 
rect 139 43 140 44 
rect 139 44 140 45 
rect 139 45 140 46 
rect 139 46 140 47 
rect 139 47 140 48 
rect 139 90 140 91 
rect 139 91 140 92 
rect 139 92 140 93 
rect 139 93 140 94 
rect 139 94 140 95 
rect 139 95 140 96 
rect 139 106 140 107 
rect 139 107 140 108 
rect 139 108 140 109 
rect 139 109 140 110 
rect 139 110 140 111 
rect 139 111 140 112 
rect 139 122 140 123 
rect 139 123 140 124 
rect 139 124 140 125 
rect 139 125 140 126 
rect 139 126 140 127 
rect 139 127 140 128 
rect 139 138 140 139 
rect 139 139 140 140 
rect 139 140 140 141 
rect 139 141 140 142 
rect 139 142 140 143 
rect 139 143 140 144 
rect 140 10 141 11 
rect 140 11 141 12 
rect 140 12 141 13 
rect 140 13 141 14 
rect 140 14 141 15 
rect 140 15 141 16 
rect 140 42 141 43 
rect 140 43 141 44 
rect 140 44 141 45 
rect 140 45 141 46 
rect 140 46 141 47 
rect 140 47 141 48 
rect 140 90 141 91 
rect 140 91 141 92 
rect 140 92 141 93 
rect 140 93 141 94 
rect 140 94 141 95 
rect 140 95 141 96 
rect 140 106 141 107 
rect 140 107 141 108 
rect 140 108 141 109 
rect 140 109 141 110 
rect 140 110 141 111 
rect 140 111 141 112 
rect 140 122 141 123 
rect 140 123 141 124 
rect 140 124 141 125 
rect 140 125 141 126 
rect 140 126 141 127 
rect 140 127 141 128 
rect 140 138 141 139 
rect 140 139 141 140 
rect 140 140 141 141 
rect 140 141 141 142 
rect 140 142 141 143 
rect 140 143 141 144 
rect 141 10 142 11 
rect 141 11 142 12 
rect 141 12 142 13 
rect 141 13 142 14 
rect 141 14 142 15 
rect 141 15 142 16 
rect 141 42 142 43 
rect 141 43 142 44 
rect 141 44 142 45 
rect 141 45 142 46 
rect 141 46 142 47 
rect 141 47 142 48 
rect 141 90 142 91 
rect 141 91 142 92 
rect 141 92 142 93 
rect 141 93 142 94 
rect 141 94 142 95 
rect 141 95 142 96 
rect 141 106 142 107 
rect 141 107 142 108 
rect 141 108 142 109 
rect 141 109 142 110 
rect 141 110 142 111 
rect 141 111 142 112 
rect 141 122 142 123 
rect 141 123 142 124 
rect 141 124 142 125 
rect 141 125 142 126 
rect 141 126 142 127 
rect 141 127 142 128 
rect 141 138 142 139 
rect 141 139 142 140 
rect 141 140 142 141 
rect 141 141 142 142 
rect 141 142 142 143 
rect 141 143 142 144 
rect 142 10 143 11 
rect 142 11 143 12 
rect 142 12 143 13 
rect 142 13 143 14 
rect 142 14 143 15 
rect 142 15 143 16 
rect 142 42 143 43 
rect 142 43 143 44 
rect 142 44 143 45 
rect 142 45 143 46 
rect 142 46 143 47 
rect 142 47 143 48 
rect 142 90 143 91 
rect 142 91 143 92 
rect 142 92 143 93 
rect 142 93 143 94 
rect 142 94 143 95 
rect 142 95 143 96 
rect 142 106 143 107 
rect 142 107 143 108 
rect 142 108 143 109 
rect 142 109 143 110 
rect 142 110 143 111 
rect 142 111 143 112 
rect 142 122 143 123 
rect 142 123 143 124 
rect 142 124 143 125 
rect 142 125 143 126 
rect 142 126 143 127 
rect 142 127 143 128 
rect 142 138 143 139 
rect 142 139 143 140 
rect 142 140 143 141 
rect 142 141 143 142 
rect 142 142 143 143 
rect 142 143 143 144 
rect 143 10 144 11 
rect 143 11 144 12 
rect 143 12 144 13 
rect 143 13 144 14 
rect 143 15 144 16 
rect 143 42 144 43 
rect 143 44 144 45 
rect 143 45 144 46 
rect 143 47 144 48 
rect 143 90 144 91 
rect 143 92 144 93 
rect 143 93 144 94 
rect 143 94 144 95 
rect 143 95 144 96 
rect 143 106 144 107 
rect 143 108 144 109 
rect 143 109 144 110 
rect 143 111 144 112 
rect 143 122 144 123 
rect 143 123 144 124 
rect 143 124 144 125 
rect 143 125 144 126 
rect 143 126 144 127 
rect 143 127 144 128 
rect 143 138 144 139 
rect 143 139 144 140 
rect 143 140 144 141 
rect 143 141 144 142 
rect 143 143 144 144 
rect 154 74 155 75 
rect 154 75 155 76 
rect 154 76 155 77 
rect 154 77 155 78 
rect 154 78 155 79 
rect 154 79 155 80 
rect 154 90 155 91 
rect 154 91 155 92 
rect 154 92 155 93 
rect 154 93 155 94 
rect 154 95 155 96 
rect 154 106 155 107 
rect 154 107 155 108 
rect 154 108 155 109 
rect 154 109 155 110 
rect 154 111 155 112 
rect 154 122 155 123 
rect 154 124 155 125 
rect 154 125 155 126 
rect 154 127 155 128 
rect 154 138 155 139 
rect 154 139 155 140 
rect 154 140 155 141 
rect 154 141 155 142 
rect 154 143 155 144 
rect 155 74 156 75 
rect 155 75 156 76 
rect 155 76 156 77 
rect 155 77 156 78 
rect 155 78 156 79 
rect 155 79 156 80 
rect 155 90 156 91 
rect 155 91 156 92 
rect 155 92 156 93 
rect 155 93 156 94 
rect 155 94 156 95 
rect 155 95 156 96 
rect 155 106 156 107 
rect 155 107 156 108 
rect 155 108 156 109 
rect 155 109 156 110 
rect 155 110 156 111 
rect 155 111 156 112 
rect 155 122 156 123 
rect 155 123 156 124 
rect 155 124 156 125 
rect 155 125 156 126 
rect 155 126 156 127 
rect 155 127 156 128 
rect 155 138 156 139 
rect 155 139 156 140 
rect 155 140 156 141 
rect 155 141 156 142 
rect 155 142 156 143 
rect 155 143 156 144 
rect 156 74 157 75 
rect 156 75 157 76 
rect 156 76 157 77 
rect 156 77 157 78 
rect 156 78 157 79 
rect 156 79 157 80 
rect 156 90 157 91 
rect 156 91 157 92 
rect 156 92 157 93 
rect 156 93 157 94 
rect 156 94 157 95 
rect 156 95 157 96 
rect 156 106 157 107 
rect 156 107 157 108 
rect 156 108 157 109 
rect 156 109 157 110 
rect 156 110 157 111 
rect 156 111 157 112 
rect 156 122 157 123 
rect 156 123 157 124 
rect 156 124 157 125 
rect 156 125 157 126 
rect 156 126 157 127 
rect 156 127 157 128 
rect 156 138 157 139 
rect 156 139 157 140 
rect 156 140 157 141 
rect 156 141 157 142 
rect 156 142 157 143 
rect 156 143 157 144 
rect 157 74 158 75 
rect 157 75 158 76 
rect 157 76 158 77 
rect 157 77 158 78 
rect 157 78 158 79 
rect 157 79 158 80 
rect 157 90 158 91 
rect 157 91 158 92 
rect 157 92 158 93 
rect 157 93 158 94 
rect 157 94 158 95 
rect 157 95 158 96 
rect 157 106 158 107 
rect 157 107 158 108 
rect 157 108 158 109 
rect 157 109 158 110 
rect 157 110 158 111 
rect 157 111 158 112 
rect 157 122 158 123 
rect 157 123 158 124 
rect 157 124 158 125 
rect 157 125 158 126 
rect 157 126 158 127 
rect 157 127 158 128 
rect 157 138 158 139 
rect 157 139 158 140 
rect 157 140 158 141 
rect 157 141 158 142 
rect 157 142 158 143 
rect 157 143 158 144 
rect 158 74 159 75 
rect 158 75 159 76 
rect 158 76 159 77 
rect 158 77 159 78 
rect 158 78 159 79 
rect 158 79 159 80 
rect 158 90 159 91 
rect 158 91 159 92 
rect 158 92 159 93 
rect 158 93 159 94 
rect 158 94 159 95 
rect 158 95 159 96 
rect 158 106 159 107 
rect 158 107 159 108 
rect 158 108 159 109 
rect 158 109 159 110 
rect 158 110 159 111 
rect 158 111 159 112 
rect 158 122 159 123 
rect 158 123 159 124 
rect 158 124 159 125 
rect 158 125 159 126 
rect 158 126 159 127 
rect 158 127 159 128 
rect 158 138 159 139 
rect 158 139 159 140 
rect 158 140 159 141 
rect 158 141 159 142 
rect 158 142 159 143 
rect 158 143 159 144 
rect 159 74 160 75 
rect 159 76 160 77 
rect 159 77 160 78 
rect 159 79 160 80 
rect 159 90 160 91 
rect 159 92 160 93 
rect 159 93 160 94 
rect 159 95 160 96 
rect 159 106 160 107 
rect 159 107 160 108 
rect 159 108 160 109 
rect 159 109 160 110 
rect 159 111 160 112 
rect 159 122 160 123 
rect 159 124 160 125 
rect 159 125 160 126 
rect 159 126 160 127 
rect 159 127 160 128 
rect 159 138 160 139 
rect 159 139 160 140 
rect 159 140 160 141 
rect 159 141 160 142 
rect 159 142 160 143 
rect 159 143 160 144 
<< labels >>
<< metal1 >>
rect 8 57 9 58 
rect 8 58 9 59 
rect 8 59 9 60 
rect 8 75 9 76 
rect 8 76 9 77 
rect 8 77 9 78 
rect 8 78 9 79 
rect 8 79 9 80 
rect 8 80 9 81 
rect 8 81 9 82 
rect 8 82 9 83 
rect 8 83 9 84 
rect 8 84 9 85 
rect 8 85 9 86 
rect 8 86 9 87 
rect 8 87 9 88 
rect 8 88 9 89 
rect 8 89 9 90 
rect 8 90 9 91 
rect 8 91 9 92 
rect 8 92 9 93 
rect 8 93 9 94 
rect 8 94 9 95 
rect 8 95 9 96 
rect 8 96 9 97 
rect 8 102 9 103 
rect 8 103 9 104 
rect 8 104 9 105 
rect 8 105 9 106 
rect 8 106 9 107 
rect 8 107 9 108 
rect 8 108 9 109 
rect 8 109 9 110 
rect 8 110 9 111 
rect 8 111 9 112 
rect 8 112 9 113 
rect 8 113 9 114 
rect 8 114 9 115 
rect 8 115 9 116 
rect 8 116 9 117 
rect 8 117 9 118 
rect 8 118 9 119 
rect 8 119 9 120 
rect 8 120 9 121 
rect 8 121 9 122 
rect 8 122 9 123 
rect 8 123 9 124 
rect 8 124 9 125 
rect 8 125 9 126 
rect 8 126 9 127 
rect 9 56 10 57 
rect 9 57 10 58 
rect 9 59 10 60 
rect 9 75 10 76 
rect 9 96 10 97 
rect 9 97 10 98 
rect 9 102 10 103 
rect 9 126 10 127 
rect 10 56 11 57 
rect 10 59 11 60 
rect 10 75 11 76 
rect 10 97 11 98 
rect 10 100 11 101 
rect 10 101 11 102 
rect 10 102 11 103 
rect 10 126 11 127 
rect 11 56 12 57 
rect 11 97 12 98 
rect 11 100 12 101 
rect 12 56 13 57 
rect 12 97 13 98 
rect 12 98 13 99 
rect 12 100 13 101 
rect 13 56 14 57 
rect 13 100 14 101 
rect 13 102 14 103 
rect 14 56 15 57 
rect 14 100 15 101 
rect 14 102 15 103 
rect 15 27 16 28 
rect 15 46 16 47 
rect 15 56 16 57 
rect 15 100 16 101 
rect 15 102 16 103 
rect 15 103 16 104 
rect 15 123 16 124 
rect 16 27 17 28 
rect 16 46 17 47 
rect 16 103 17 104 
rect 16 104 17 105 
rect 16 123 17 124 
rect 17 27 18 28 
rect 17 46 18 47 
rect 17 47 18 48 
rect 17 48 18 49 
rect 17 49 18 50 
rect 17 50 18 51 
rect 17 51 18 52 
rect 17 52 18 53 
rect 17 53 18 54 
rect 17 54 18 55 
rect 17 55 18 56 
rect 17 56 18 57 
rect 17 57 18 58 
rect 17 58 18 59 
rect 17 59 18 60 
rect 17 60 18 61 
rect 17 61 18 62 
rect 17 62 18 63 
rect 17 63 18 64 
rect 17 64 18 65 
rect 17 65 18 66 
rect 17 66 18 67 
rect 17 67 18 68 
rect 17 68 18 69 
rect 17 69 18 70 
rect 17 70 18 71 
rect 17 71 18 72 
rect 17 72 18 73 
rect 17 73 18 74 
rect 17 74 18 75 
rect 17 75 18 76 
rect 17 76 18 77 
rect 17 77 18 78 
rect 17 78 18 79 
rect 17 79 18 80 
rect 17 80 18 81 
rect 17 81 18 82 
rect 17 82 18 83 
rect 17 83 18 84 
rect 17 84 18 85 
rect 17 85 18 86 
rect 17 86 18 87 
rect 17 87 18 88 
rect 17 88 18 89 
rect 17 89 18 90 
rect 17 90 18 91 
rect 17 91 18 92 
rect 17 92 18 93 
rect 17 93 18 94 
rect 17 94 18 95 
rect 17 95 18 96 
rect 17 96 18 97 
rect 17 97 18 98 
rect 17 98 18 99 
rect 17 99 18 100 
rect 17 100 18 101 
rect 17 101 18 102 
rect 17 102 18 103 
rect 17 104 18 105 
rect 17 105 18 106 
rect 17 106 18 107 
rect 17 107 18 108 
rect 17 119 18 120 
rect 17 120 18 121 
rect 17 121 18 122 
rect 17 122 18 123 
rect 17 123 18 124 
rect 18 27 19 28 
rect 18 102 19 103 
rect 18 107 19 108 
rect 18 119 19 120 
rect 19 27 20 28 
rect 19 47 20 48 
rect 19 48 20 49 
rect 19 49 20 50 
rect 19 50 20 51 
rect 19 51 20 52 
rect 19 52 20 53 
rect 19 53 20 54 
rect 19 54 20 55 
rect 19 55 20 56 
rect 19 102 20 103 
rect 19 107 20 108 
rect 19 119 20 120 
rect 20 27 21 28 
rect 20 36 21 37 
rect 20 37 21 38 
rect 20 38 21 39 
rect 20 39 21 40 
rect 20 40 21 41 
rect 20 41 21 42 
rect 20 42 21 43 
rect 20 47 21 48 
rect 20 100 21 101 
rect 20 102 21 103 
rect 20 107 21 108 
rect 20 119 21 120 
rect 21 27 22 28 
rect 21 36 22 37 
rect 21 42 22 43 
rect 21 43 22 44 
rect 21 44 22 45 
rect 21 47 22 48 
rect 21 49 22 50 
rect 21 50 22 51 
rect 21 100 22 101 
rect 21 102 22 103 
rect 21 107 22 108 
rect 21 119 22 120 
rect 22 27 23 28 
rect 22 36 23 37 
rect 22 47 23 48 
rect 22 50 23 51 
rect 22 51 23 52 
rect 22 52 23 53 
rect 22 53 23 54 
rect 22 54 23 55 
rect 22 55 23 56 
rect 22 56 23 57 
rect 22 57 23 58 
rect 22 58 23 59 
rect 22 59 23 60 
rect 22 60 23 61 
rect 22 61 23 62 
rect 22 62 23 63 
rect 22 63 23 64 
rect 22 64 23 65 
rect 22 65 23 66 
rect 22 66 23 67 
rect 22 67 23 68 
rect 22 68 23 69 
rect 22 69 23 70 
rect 22 70 23 71 
rect 22 71 23 72 
rect 22 72 23 73 
rect 22 73 23 74 
rect 22 74 23 75 
rect 22 75 23 76 
rect 22 76 23 77 
rect 22 77 23 78 
rect 22 78 23 79 
rect 22 79 23 80 
rect 22 80 23 81 
rect 22 81 23 82 
rect 22 82 23 83 
rect 22 83 23 84 
rect 22 84 23 85 
rect 22 85 23 86 
rect 22 86 23 87 
rect 22 87 23 88 
rect 22 88 23 89 
rect 22 89 23 90 
rect 22 90 23 91 
rect 22 91 23 92 
rect 22 92 23 93 
rect 22 100 23 101 
rect 22 102 23 103 
rect 22 107 23 108 
rect 22 119 23 120 
rect 23 23 24 24 
rect 23 24 24 25 
rect 23 25 24 26 
rect 23 26 24 27 
rect 23 27 24 28 
rect 23 34 24 35 
rect 23 35 24 36 
rect 23 36 24 37 
rect 23 43 24 44 
rect 23 44 24 45 
rect 23 45 24 46 
rect 23 47 24 48 
rect 23 92 24 93 
rect 23 93 24 94 
rect 23 99 24 100 
rect 23 100 24 101 
rect 23 102 24 103 
rect 23 107 24 108 
rect 23 108 24 109 
rect 23 109 24 110 
rect 23 110 24 111 
rect 23 111 24 112 
rect 23 112 24 113 
rect 23 113 24 114 
rect 23 114 24 115 
rect 23 119 24 120 
rect 23 140 24 141 
rect 23 141 24 142 
rect 23 142 24 143 
rect 23 143 24 144 
rect 23 144 24 145 
rect 23 145 24 146 
rect 23 146 24 147 
rect 23 147 24 148 
rect 23 148 24 149 
rect 23 149 24 150 
rect 23 150 24 151 
rect 24 23 25 24 
rect 24 34 25 35 
rect 24 43 25 44 
rect 24 46 25 47 
rect 24 47 25 48 
rect 24 49 25 50 
rect 24 89 25 90 
rect 24 90 25 91 
rect 24 91 25 92 
rect 24 93 25 94 
rect 24 94 25 95 
rect 24 99 25 100 
rect 24 102 25 103 
rect 24 114 25 115 
rect 24 119 25 120 
rect 24 139 25 140 
rect 24 140 25 141 
rect 24 150 25 151 
rect 24 153 25 154 
rect 24 154 25 155 
rect 24 155 25 156 
rect 25 23 26 24 
rect 25 34 26 35 
rect 25 43 26 44 
rect 25 46 26 47 
rect 25 49 26 50 
rect 25 88 26 89 
rect 25 89 26 90 
rect 25 91 26 92 
rect 25 94 26 95 
rect 25 99 26 100 
rect 25 102 26 103 
rect 25 114 26 115 
rect 25 119 26 120 
rect 25 139 26 140 
rect 25 150 26 151 
rect 25 152 26 153 
rect 25 153 26 154 
rect 25 155 26 156 
rect 26 23 27 24 
rect 26 34 27 35 
rect 26 43 27 44 
rect 26 46 27 47 
rect 26 49 27 50 
rect 26 88 27 89 
rect 26 91 27 92 
rect 26 94 27 95 
rect 26 99 27 100 
rect 26 102 27 103 
rect 26 114 27 115 
rect 26 119 27 120 
rect 26 139 27 140 
rect 26 150 27 151 
rect 26 152 27 153 
rect 26 155 27 156 
rect 27 23 28 24 
rect 27 34 28 35 
rect 27 49 28 50 
rect 27 50 28 51 
rect 27 51 28 52 
rect 27 52 28 53 
rect 27 53 28 54 
rect 27 54 28 55 
rect 27 55 28 56 
rect 27 58 28 59 
rect 27 59 28 60 
rect 27 60 28 61 
rect 27 61 28 62 
rect 27 62 28 63 
rect 27 63 28 64 
rect 27 64 28 65 
rect 27 65 28 66 
rect 27 66 28 67 
rect 27 67 28 68 
rect 27 68 28 69 
rect 27 69 28 70 
rect 27 70 28 71 
rect 27 71 28 72 
rect 27 72 28 73 
rect 27 73 28 74 
rect 27 74 28 75 
rect 27 75 28 76 
rect 27 76 28 77 
rect 27 77 28 78 
rect 27 78 28 79 
rect 27 79 28 80 
rect 27 80 28 81 
rect 27 81 28 82 
rect 27 82 28 83 
rect 27 83 28 84 
rect 27 84 28 85 
rect 27 85 28 86 
rect 27 86 28 87 
rect 27 87 28 88 
rect 27 88 28 89 
rect 27 97 28 98 
rect 27 98 28 99 
rect 27 99 28 100 
rect 27 102 28 103 
rect 27 103 28 104 
rect 27 114 28 115 
rect 27 119 28 120 
rect 27 150 28 151 
rect 27 152 28 153 
rect 28 23 29 24 
rect 28 34 29 35 
rect 28 55 29 56 
rect 28 58 29 59 
rect 28 97 29 98 
rect 28 103 29 104 
rect 28 114 29 115 
rect 28 119 29 120 
rect 28 150 29 151 
rect 28 152 29 153 
rect 29 23 30 24 
rect 29 34 30 35 
rect 29 55 30 56 
rect 29 58 30 59 
rect 29 97 30 98 
rect 29 103 30 104 
rect 29 114 30 115 
rect 29 119 30 120 
rect 29 150 30 151 
rect 29 152 30 153 
rect 30 23 31 24 
rect 30 34 31 35 
rect 30 55 31 56 
rect 30 58 31 59 
rect 30 97 31 98 
rect 30 103 31 104 
rect 30 114 31 115 
rect 30 119 31 120 
rect 30 152 31 153 
rect 31 11 32 12 
rect 31 23 32 24 
rect 31 27 32 28 
rect 31 34 32 35 
rect 31 46 32 47 
rect 31 55 32 56 
rect 31 58 32 59 
rect 31 97 32 98 
rect 31 103 32 104 
rect 31 107 32 108 
rect 31 114 32 115 
rect 31 115 32 116 
rect 31 116 32 117 
rect 31 119 32 120 
rect 31 148 32 149 
rect 31 149 32 150 
rect 31 150 32 151 
rect 31 151 32 152 
rect 31 152 32 153 
rect 31 158 32 159 
rect 32 11 33 12 
rect 32 23 33 24 
rect 32 27 33 28 
rect 32 34 33 35 
rect 32 46 33 47 
rect 32 55 33 56 
rect 32 58 33 59 
rect 32 96 33 97 
rect 32 97 33 98 
rect 32 103 33 104 
rect 32 107 33 108 
rect 32 148 33 149 
rect 32 158 33 159 
rect 33 11 34 12 
rect 33 23 34 24 
rect 33 27 34 28 
rect 33 28 34 29 
rect 33 29 34 30 
rect 33 30 34 31 
rect 33 31 34 32 
rect 33 32 34 33 
rect 33 34 34 35 
rect 33 46 34 47 
rect 33 47 34 48 
rect 33 48 34 49 
rect 33 49 34 50 
rect 33 50 34 51 
rect 33 51 34 52 
rect 33 52 34 53 
rect 33 53 34 54 
rect 33 55 34 56 
rect 33 58 34 59 
rect 33 82 34 83 
rect 33 83 34 84 
rect 33 84 34 85 
rect 33 85 34 86 
rect 33 86 34 87 
rect 33 87 34 88 
rect 33 88 34 89 
rect 33 89 34 90 
rect 33 90 34 91 
rect 33 91 34 92 
rect 33 92 34 93 
rect 33 93 34 94 
rect 33 94 34 95 
rect 33 95 34 96 
rect 33 96 34 97 
rect 33 103 34 104 
rect 33 107 34 108 
rect 33 108 34 109 
rect 33 109 34 110 
rect 33 110 34 111 
rect 33 111 34 112 
rect 33 112 34 113 
rect 33 113 34 114 
rect 33 114 34 115 
rect 33 115 34 116 
rect 33 116 34 117 
rect 33 117 34 118 
rect 33 118 34 119 
rect 33 119 34 120 
rect 33 120 34 121 
rect 33 121 34 122 
rect 33 122 34 123 
rect 33 123 34 124 
rect 33 124 34 125 
rect 33 125 34 126 
rect 33 126 34 127 
rect 33 127 34 128 
rect 33 128 34 129 
rect 33 129 34 130 
rect 33 130 34 131 
rect 33 131 34 132 
rect 33 132 34 133 
rect 33 133 34 134 
rect 33 134 34 135 
rect 33 135 34 136 
rect 33 136 34 137 
rect 33 137 34 138 
rect 33 138 34 139 
rect 33 139 34 140 
rect 33 140 34 141 
rect 33 141 34 142 
rect 33 142 34 143 
rect 33 143 34 144 
rect 33 144 34 145 
rect 33 145 34 146 
rect 33 146 34 147 
rect 33 147 34 148 
rect 33 148 34 149 
rect 33 151 34 152 
rect 33 158 34 159 
rect 34 11 35 12 
rect 34 23 35 24 
rect 34 32 35 33 
rect 34 34 35 35 
rect 34 53 35 54 
rect 34 55 35 56 
rect 34 58 35 59 
rect 34 82 35 83 
rect 34 103 35 104 
rect 34 151 35 152 
rect 34 158 35 159 
rect 35 11 36 12 
rect 35 23 36 24 
rect 35 32 36 33 
rect 35 34 36 35 
rect 35 53 36 54 
rect 35 55 36 56 
rect 35 58 36 59 
rect 35 82 36 83 
rect 35 103 36 104 
rect 35 104 36 105 
rect 35 105 36 106 
rect 35 106 36 107 
rect 35 107 36 108 
rect 35 108 36 109 
rect 35 109 36 110 
rect 35 110 36 111 
rect 35 111 36 112 
rect 35 112 36 113 
rect 35 113 36 114 
rect 35 114 36 115 
rect 35 115 36 116 
rect 35 116 36 117 
rect 35 117 36 118 
rect 35 118 36 119 
rect 35 119 36 120 
rect 35 120 36 121 
rect 35 121 36 122 
rect 35 122 36 123 
rect 35 123 36 124 
rect 35 124 36 125 
rect 35 125 36 126 
rect 35 126 36 127 
rect 35 127 36 128 
rect 35 128 36 129 
rect 35 129 36 130 
rect 35 130 36 131 
rect 35 131 36 132 
rect 35 132 36 133 
rect 35 133 36 134 
rect 35 134 36 135 
rect 35 135 36 136 
rect 35 151 36 152 
rect 35 158 36 159 
rect 36 11 37 12 
rect 36 23 37 24 
rect 36 32 37 33 
rect 36 34 37 35 
rect 36 53 37 54 
rect 36 55 37 56 
rect 36 58 37 59 
rect 36 82 37 83 
rect 36 135 37 136 
rect 36 151 37 152 
rect 36 158 37 159 
rect 37 11 38 12 
rect 37 23 38 24 
rect 37 32 38 33 
rect 37 34 38 35 
rect 37 53 38 54 
rect 37 55 38 56 
rect 37 58 38 59 
rect 37 82 38 83 
rect 37 113 38 114 
rect 37 114 38 115 
rect 37 115 38 116 
rect 37 116 38 117 
rect 37 117 38 118 
rect 37 118 38 119 
rect 37 135 38 136 
rect 37 151 38 152 
rect 37 158 38 159 
rect 38 11 39 12 
rect 38 23 39 24 
rect 38 32 39 33 
rect 38 34 39 35 
rect 38 53 39 54 
rect 38 55 39 56 
rect 38 58 39 59 
rect 38 82 39 83 
rect 38 113 39 114 
rect 38 135 39 136 
rect 38 151 39 152 
rect 38 158 39 159 
rect 39 11 40 12 
rect 39 23 40 24 
rect 39 32 40 33 
rect 39 34 40 35 
rect 39 53 40 54 
rect 39 55 40 56 
rect 39 58 40 59 
rect 39 82 40 83 
rect 39 113 40 114 
rect 39 117 40 118 
rect 39 135 40 136 
rect 39 151 40 152 
rect 39 157 40 158 
rect 39 158 40 159 
rect 40 9 41 10 
rect 40 10 41 11 
rect 40 11 41 12 
rect 40 14 41 15 
rect 40 15 41 16 
rect 40 16 41 17 
rect 40 23 41 24 
rect 40 34 41 35 
rect 40 46 41 47 
rect 40 47 41 48 
rect 40 48 41 49 
rect 40 53 41 54 
rect 40 55 41 56 
rect 40 58 41 59 
rect 40 60 41 61 
rect 40 72 41 73 
rect 40 73 41 74 
rect 40 74 41 75 
rect 40 75 41 76 
rect 40 76 41 77 
rect 40 77 41 78 
rect 40 78 41 79 
rect 40 79 41 80 
rect 40 82 41 83 
rect 40 84 41 85 
rect 40 85 41 86 
rect 40 86 41 87 
rect 40 87 41 88 
rect 40 88 41 89 
rect 40 89 41 90 
rect 40 90 41 91 
rect 40 91 41 92 
rect 40 92 41 93 
rect 40 93 41 94 
rect 40 94 41 95 
rect 40 103 41 104 
rect 40 104 41 105 
rect 40 105 41 106 
rect 40 106 41 107 
rect 40 107 41 108 
rect 40 108 41 109 
rect 40 109 41 110 
rect 40 110 41 111 
rect 40 111 41 112 
rect 40 113 41 114 
rect 40 117 41 118 
rect 40 118 41 119 
rect 40 119 41 120 
rect 40 120 41 121 
rect 40 121 41 122 
rect 40 122 41 123 
rect 40 123 41 124 
rect 40 135 41 136 
rect 40 137 41 138 
rect 40 138 41 139 
rect 40 139 41 140 
rect 40 140 41 141 
rect 40 141 41 142 
rect 40 142 41 143 
rect 40 151 41 152 
rect 40 153 41 154 
rect 40 154 41 155 
rect 40 155 41 156 
rect 41 8 42 9 
rect 41 9 42 10 
rect 41 14 42 15 
rect 41 16 42 17 
rect 41 17 42 18 
rect 41 23 42 24 
rect 41 34 42 35 
rect 41 46 42 47 
rect 41 48 42 49 
rect 41 49 42 50 
rect 41 53 42 54 
rect 41 55 42 56 
rect 41 58 42 59 
rect 41 60 42 61 
rect 41 61 42 62 
rect 41 62 42 63 
rect 41 63 42 64 
rect 41 64 42 65 
rect 41 65 42 66 
rect 41 66 42 67 
rect 41 67 42 68 
rect 41 68 42 69 
rect 41 69 42 70 
rect 41 70 42 71 
rect 41 71 42 72 
rect 41 72 42 73 
rect 41 82 42 83 
rect 41 94 42 95 
rect 41 103 42 104 
rect 41 113 42 114 
rect 41 123 42 124 
rect 41 135 42 136 
rect 41 142 42 143 
rect 41 151 42 152 
rect 41 153 42 154 
rect 41 155 42 156 
rect 42 8 43 9 
rect 42 14 43 15 
rect 42 17 43 18 
rect 42 18 43 19 
rect 42 19 43 20 
rect 42 20 43 21 
rect 42 21 43 22 
rect 42 23 43 24 
rect 42 34 43 35 
rect 42 46 43 47 
rect 42 49 43 50 
rect 42 53 43 54 
rect 42 55 43 56 
rect 42 58 43 59 
rect 42 82 43 83 
rect 42 94 43 95 
rect 42 103 43 104 
rect 42 113 43 114 
rect 42 123 43 124 
rect 42 133 43 134 
rect 42 135 43 136 
rect 42 142 43 143 
rect 42 149 43 150 
rect 42 151 43 152 
rect 42 155 43 156 
rect 43 8 44 9 
rect 43 21 44 22 
rect 43 23 44 24 
rect 43 34 44 35 
rect 43 49 44 50 
rect 43 53 44 54 
rect 43 55 44 56 
rect 43 58 44 59 
rect 43 82 44 83 
rect 43 98 44 99 
rect 43 99 44 100 
rect 43 100 44 101 
rect 43 101 44 102 
rect 43 102 44 103 
rect 43 103 44 104 
rect 43 113 44 114 
rect 43 130 44 131 
rect 43 131 44 132 
rect 43 132 44 133 
rect 43 133 44 134 
rect 43 135 44 136 
rect 43 149 44 150 
rect 43 151 44 152 
rect 44 8 45 9 
rect 44 21 45 22 
rect 44 23 45 24 
rect 44 34 45 35 
rect 44 49 45 50 
rect 44 53 45 54 
rect 44 55 45 56 
rect 44 58 45 59 
rect 44 82 45 83 
rect 44 98 45 99 
rect 44 113 45 114 
rect 44 130 45 131 
rect 44 135 45 136 
rect 44 149 45 150 
rect 44 151 45 152 
rect 45 8 46 9 
rect 45 21 46 22 
rect 45 23 46 24 
rect 45 34 46 35 
rect 45 49 46 50 
rect 45 53 46 54 
rect 45 55 46 56 
rect 45 58 46 59 
rect 45 82 46 83 
rect 45 98 46 99 
rect 45 113 46 114 
rect 45 130 46 131 
rect 45 135 46 136 
rect 45 149 46 150 
rect 45 151 46 152 
rect 46 8 47 9 
rect 46 21 47 22 
rect 46 23 47 24 
rect 46 34 47 35 
rect 46 49 47 50 
rect 46 53 47 54 
rect 46 55 47 56 
rect 46 58 47 59 
rect 46 82 47 83 
rect 46 98 47 99 
rect 46 113 47 114 
rect 46 130 47 131 
rect 46 135 47 136 
rect 46 149 47 150 
rect 46 151 47 152 
rect 47 8 48 9 
rect 47 21 48 22 
rect 47 23 48 24 
rect 47 27 48 28 
rect 47 33 48 34 
rect 47 34 48 35 
rect 47 43 48 44 
rect 47 49 48 50 
rect 47 53 48 54 
rect 47 55 48 56 
rect 47 57 48 58 
rect 47 58 48 59 
rect 47 75 48 76 
rect 47 78 48 79 
rect 47 82 48 83 
rect 47 91 48 92 
rect 47 94 48 95 
rect 47 98 48 99 
rect 47 110 48 111 
rect 47 113 48 114 
rect 47 130 48 131 
rect 47 135 48 136 
rect 47 136 48 137 
rect 47 142 48 143 
rect 47 147 48 148 
rect 47 148 48 149 
rect 47 149 48 150 
rect 47 151 48 152 
rect 47 152 48 153 
rect 48 8 49 9 
rect 48 21 49 22 
rect 48 23 49 24 
rect 48 27 49 28 
rect 48 32 49 33 
rect 48 33 49 34 
rect 48 43 49 44 
rect 48 49 49 50 
rect 48 51 49 52 
rect 48 53 49 54 
rect 48 55 49 56 
rect 48 75 49 76 
rect 48 78 49 79 
rect 48 82 49 83 
rect 48 91 49 92 
rect 48 94 49 95 
rect 48 110 49 111 
rect 48 112 49 113 
rect 48 113 49 114 
rect 48 130 49 131 
rect 48 136 49 137 
rect 48 142 49 143 
rect 48 147 49 148 
rect 48 152 49 153 
rect 48 153 49 154 
rect 49 8 50 9 
rect 49 21 50 22 
rect 49 23 50 24 
rect 49 27 50 28 
rect 49 28 50 29 
rect 49 29 50 30 
rect 49 30 50 31 
rect 49 31 50 32 
rect 49 32 50 33 
rect 49 43 50 44 
rect 49 49 50 50 
rect 49 51 50 52 
rect 49 53 50 54 
rect 49 55 50 56 
rect 49 73 50 74 
rect 49 75 50 76 
rect 49 78 50 79 
rect 49 82 50 83 
rect 49 91 50 92 
rect 49 94 50 95 
rect 49 95 50 96 
rect 49 96 50 97 
rect 49 97 50 98 
rect 49 98 50 99 
rect 49 99 50 100 
rect 49 100 50 101 
rect 49 101 50 102 
rect 49 102 50 103 
rect 49 103 50 104 
rect 49 104 50 105 
rect 49 105 50 106 
rect 49 106 50 107 
rect 49 107 50 108 
rect 49 108 50 109 
rect 49 110 50 111 
rect 49 111 50 112 
rect 49 112 50 113 
rect 49 130 50 131 
rect 49 136 50 137 
rect 49 142 50 143 
rect 49 147 50 148 
rect 49 153 50 154 
rect 49 154 50 155 
rect 49 155 50 156 
rect 50 8 51 9 
rect 50 21 51 22 
rect 50 23 51 24 
rect 50 49 51 50 
rect 50 51 51 52 
rect 50 53 51 54 
rect 50 55 51 56 
rect 50 73 51 74 
rect 50 75 51 76 
rect 50 78 51 79 
rect 50 79 51 80 
rect 50 80 51 81 
rect 50 82 51 83 
rect 50 91 51 92 
rect 50 108 51 109 
rect 50 109 51 110 
rect 50 130 51 131 
rect 50 136 51 137 
rect 50 142 51 143 
rect 50 147 51 148 
rect 50 155 51 156 
rect 51 8 52 9 
rect 51 21 52 22 
rect 51 23 52 24 
rect 51 24 52 25 
rect 51 25 52 26 
rect 51 26 52 27 
rect 51 27 52 28 
rect 51 28 52 29 
rect 51 29 52 30 
rect 51 30 52 31 
rect 51 31 52 32 
rect 51 32 52 33 
rect 51 33 52 34 
rect 51 34 52 35 
rect 51 35 52 36 
rect 51 36 52 37 
rect 51 37 52 38 
rect 51 38 52 39 
rect 51 39 52 40 
rect 51 47 52 48 
rect 51 49 52 50 
rect 51 51 52 52 
rect 51 53 52 54 
rect 51 55 52 56 
rect 51 73 52 74 
rect 51 75 52 76 
rect 51 80 52 81 
rect 51 82 52 83 
rect 51 91 52 92 
rect 51 109 52 110 
rect 51 110 52 111 
rect 51 111 52 112 
rect 51 112 52 113 
rect 51 113 52 114 
rect 51 114 52 115 
rect 51 115 52 116 
rect 51 116 52 117 
rect 51 117 52 118 
rect 51 118 52 119 
rect 51 119 52 120 
rect 51 120 52 121 
rect 51 121 52 122 
rect 51 122 52 123 
rect 51 123 52 124 
rect 51 130 52 131 
rect 51 136 52 137 
rect 51 142 52 143 
rect 51 147 52 148 
rect 51 155 52 156 
rect 52 8 53 9 
rect 52 21 53 22 
rect 52 22 53 23 
rect 52 39 53 40 
rect 52 47 53 48 
rect 52 49 53 50 
rect 52 51 53 52 
rect 52 53 53 54 
rect 52 55 53 56 
rect 52 57 53 58 
rect 52 58 53 59 
rect 52 59 53 60 
rect 52 60 53 61 
rect 52 61 53 62 
rect 52 62 53 63 
rect 52 63 53 64 
rect 52 64 53 65 
rect 52 65 53 66 
rect 52 66 53 67 
rect 52 67 53 68 
rect 52 68 53 69 
rect 52 69 53 70 
rect 52 70 53 71 
rect 52 71 53 72 
rect 52 72 53 73 
rect 52 73 53 74 
rect 52 75 53 76 
rect 52 80 53 81 
rect 52 82 53 83 
rect 52 91 53 92 
rect 52 94 53 95 
rect 52 95 53 96 
rect 52 123 53 124 
rect 52 130 53 131 
rect 52 136 53 137 
rect 52 142 53 143 
rect 52 147 53 148 
rect 52 155 53 156 
rect 53 8 54 9 
rect 53 22 54 23 
rect 53 23 54 24 
rect 53 24 54 25 
rect 53 25 54 26 
rect 53 26 54 27 
rect 53 27 54 28 
rect 53 28 54 29 
rect 53 29 54 30 
rect 53 30 54 31 
rect 53 31 54 32 
rect 53 32 54 33 
rect 53 37 54 38 
rect 53 39 54 40 
rect 53 47 54 48 
rect 53 49 54 50 
rect 53 51 54 52 
rect 53 53 54 54 
rect 53 55 54 56 
rect 53 75 54 76 
rect 53 80 54 81 
rect 53 82 54 83 
rect 53 91 54 92 
rect 53 95 54 96 
rect 53 96 54 97 
rect 53 97 54 98 
rect 53 98 54 99 
rect 53 99 54 100 
rect 53 100 54 101 
rect 53 101 54 102 
rect 53 102 54 103 
rect 53 103 54 104 
rect 53 104 54 105 
rect 53 105 54 106 
rect 53 106 54 107 
rect 53 107 54 108 
rect 53 108 54 109 
rect 53 109 54 110 
rect 53 110 54 111 
rect 53 111 54 112 
rect 53 112 54 113 
rect 53 113 54 114 
rect 53 114 54 115 
rect 53 115 54 116 
rect 53 116 54 117 
rect 53 117 54 118 
rect 53 118 54 119 
rect 53 119 54 120 
rect 53 120 54 121 
rect 53 121 54 122 
rect 53 123 54 124 
rect 53 126 54 127 
rect 53 127 54 128 
rect 53 128 54 129 
rect 53 129 54 130 
rect 53 130 54 131 
rect 53 136 54 137 
rect 53 142 54 143 
rect 53 147 54 148 
rect 53 155 54 156 
rect 54 8 55 9 
rect 54 32 55 33 
rect 54 34 55 35 
rect 54 37 55 38 
rect 54 39 55 40 
rect 54 47 55 48 
rect 54 49 55 50 
rect 54 51 55 52 
rect 54 53 55 54 
rect 54 55 55 56 
rect 54 58 55 59 
rect 54 59 55 60 
rect 54 60 55 61 
rect 54 61 55 62 
rect 54 62 55 63 
rect 54 63 55 64 
rect 54 64 55 65 
rect 54 65 55 66 
rect 54 66 55 67 
rect 54 67 55 68 
rect 54 68 55 69 
rect 54 69 55 70 
rect 54 70 55 71 
rect 54 71 55 72 
rect 54 72 55 73 
rect 54 73 55 74 
rect 54 74 55 75 
rect 54 75 55 76 
rect 54 82 55 83 
rect 54 91 55 92 
rect 54 93 55 94 
rect 54 123 55 124 
rect 54 132 55 133 
rect 54 133 55 134 
rect 54 136 55 137 
rect 54 138 55 139 
rect 54 139 55 140 
rect 54 140 55 141 
rect 54 142 55 143 
rect 54 143 55 144 
rect 54 147 55 148 
rect 54 155 55 156 
rect 55 8 56 9 
rect 55 30 56 31 
rect 55 32 56 33 
rect 55 34 56 35 
rect 55 37 56 38 
rect 55 39 56 40 
rect 55 47 56 48 
rect 55 49 56 50 
rect 55 51 56 52 
rect 55 53 56 54 
rect 55 55 56 56 
rect 55 58 56 59 
rect 55 82 56 83 
rect 55 91 56 92 
rect 55 93 56 94 
rect 55 120 56 121 
rect 55 123 56 124 
rect 55 125 56 126 
rect 55 126 56 127 
rect 55 127 56 128 
rect 55 128 56 129 
rect 55 129 56 130 
rect 55 130 56 131 
rect 55 131 56 132 
rect 55 132 56 133 
rect 55 136 56 137 
rect 55 140 56 141 
rect 55 141 56 142 
rect 55 143 56 144 
rect 55 144 56 145 
rect 55 147 56 148 
rect 55 155 56 156 
rect 56 8 57 9 
rect 56 11 57 12 
rect 56 12 57 13 
rect 56 13 57 14 
rect 56 14 57 15 
rect 56 15 57 16 
rect 56 16 57 17 
rect 56 17 57 18 
rect 56 18 57 19 
rect 56 19 57 20 
rect 56 20 57 21 
rect 56 21 57 22 
rect 56 22 57 23 
rect 56 23 57 24 
rect 56 24 57 25 
rect 56 25 57 26 
rect 56 26 57 27 
rect 56 27 57 28 
rect 56 28 57 29 
rect 56 29 57 30 
rect 56 30 57 31 
rect 56 32 57 33 
rect 56 34 57 35 
rect 56 37 57 38 
rect 56 39 57 40 
rect 56 46 57 47 
rect 56 47 57 48 
rect 56 49 57 50 
rect 56 51 57 52 
rect 56 53 57 54 
rect 56 55 57 56 
rect 56 59 57 60 
rect 56 60 57 61 
rect 56 61 57 62 
rect 56 62 57 63 
rect 56 63 57 64 
rect 56 64 57 65 
rect 56 65 57 66 
rect 56 66 57 67 
rect 56 67 57 68 
rect 56 68 57 69 
rect 56 69 57 70 
rect 56 70 57 71 
rect 56 71 57 72 
rect 56 72 57 73 
rect 56 73 57 74 
rect 56 74 57 75 
rect 56 75 57 76 
rect 56 76 57 77 
rect 56 77 57 78 
rect 56 78 57 79 
rect 56 79 57 80 
rect 56 80 57 81 
rect 56 82 57 83 
rect 56 91 57 92 
rect 56 93 57 94 
rect 56 94 57 95 
rect 56 95 57 96 
rect 56 96 57 97 
rect 56 97 57 98 
rect 56 98 57 99 
rect 56 99 57 100 
rect 56 100 57 101 
rect 56 101 57 102 
rect 56 102 57 103 
rect 56 103 57 104 
rect 56 104 57 105 
rect 56 105 57 106 
rect 56 106 57 107 
rect 56 107 57 108 
rect 56 108 57 109 
rect 56 109 57 110 
rect 56 110 57 111 
rect 56 111 57 112 
rect 56 112 57 113 
rect 56 113 57 114 
rect 56 114 57 115 
rect 56 115 57 116 
rect 56 116 57 117 
rect 56 117 57 118 
rect 56 118 57 119 
rect 56 119 57 120 
rect 56 120 57 121 
rect 56 123 57 124 
rect 56 136 57 137 
rect 56 138 57 139 
rect 56 139 57 140 
rect 56 141 57 142 
rect 56 142 57 143 
rect 56 144 57 145 
rect 56 147 57 148 
rect 56 155 57 156 
rect 57 8 58 9 
rect 57 11 58 12 
rect 57 32 58 33 
rect 57 34 58 35 
rect 57 37 58 38 
rect 57 39 58 40 
rect 57 46 58 47 
rect 57 49 58 50 
rect 57 51 58 52 
rect 57 53 58 54 
rect 57 55 58 56 
rect 57 59 58 60 
rect 57 80 58 81 
rect 57 81 58 82 
rect 57 123 58 124 
rect 57 134 58 135 
rect 57 136 58 137 
rect 57 139 58 140 
rect 57 142 58 143 
rect 57 144 58 145 
rect 57 145 58 146 
rect 57 147 58 148 
rect 57 155 58 156 
rect 58 8 59 9 
rect 58 11 59 12 
rect 58 34 59 35 
rect 58 36 59 37 
rect 58 37 59 38 
rect 58 39 59 40 
rect 58 46 59 47 
rect 58 49 59 50 
rect 58 51 59 52 
rect 58 53 59 54 
rect 58 55 59 56 
rect 58 59 59 60 
rect 58 81 59 82 
rect 58 82 59 83 
rect 58 83 59 84 
rect 58 84 59 85 
rect 58 85 59 86 
rect 58 86 59 87 
rect 58 87 59 88 
rect 58 88 59 89 
rect 58 89 59 90 
rect 58 90 59 91 
rect 58 91 59 92 
rect 58 92 59 93 
rect 58 93 59 94 
rect 58 94 59 95 
rect 58 95 59 96 
rect 58 96 59 97 
rect 58 97 59 98 
rect 58 98 59 99 
rect 58 99 59 100 
rect 58 100 59 101 
rect 58 101 59 102 
rect 58 102 59 103 
rect 58 123 59 124 
rect 58 133 59 134 
rect 58 134 59 135 
rect 58 136 59 137 
rect 58 139 59 140 
rect 58 142 59 143 
rect 58 145 59 146 
rect 58 147 59 148 
rect 58 155 59 156 
rect 59 8 60 9 
rect 59 34 60 35 
rect 59 36 60 37 
rect 59 39 60 40 
rect 59 49 60 50 
rect 59 51 60 52 
rect 59 53 60 54 
rect 59 55 60 56 
rect 59 102 60 103 
rect 59 123 60 124 
rect 59 133 60 134 
rect 59 136 60 137 
rect 59 145 60 146 
rect 59 147 60 148 
rect 60 8 61 9 
rect 60 34 61 35 
rect 60 36 61 37 
rect 60 39 61 40 
rect 60 49 61 50 
rect 60 51 61 52 
rect 60 53 61 54 
rect 60 55 61 56 
rect 60 102 61 103 
rect 60 123 61 124 
rect 60 133 61 134 
rect 60 136 61 137 
rect 60 145 61 146 
rect 60 147 61 148 
rect 61 8 62 9 
rect 61 34 62 35 
rect 61 36 62 37 
rect 61 39 62 40 
rect 61 49 62 50 
rect 61 51 62 52 
rect 61 53 62 54 
rect 61 55 62 56 
rect 61 102 62 103 
rect 61 123 62 124 
rect 61 133 62 134 
rect 61 136 62 137 
rect 61 145 62 146 
rect 61 147 62 148 
rect 62 8 63 9 
rect 62 34 63 35 
rect 62 36 63 37 
rect 62 39 63 40 
rect 62 49 63 50 
rect 62 51 63 52 
rect 62 53 63 54 
rect 62 55 63 56 
rect 62 102 63 103 
rect 62 123 63 124 
rect 62 133 63 134 
rect 62 136 63 137 
rect 62 145 63 146 
rect 62 147 63 148 
rect 63 8 64 9 
rect 63 27 64 28 
rect 63 34 64 35 
rect 63 39 64 40 
rect 63 43 64 44 
rect 63 49 64 50 
rect 63 51 64 52 
rect 63 53 64 54 
rect 63 55 64 56 
rect 63 59 64 60 
rect 63 62 64 63 
rect 63 102 64 103 
rect 63 123 64 124 
rect 63 133 64 134 
rect 63 136 64 137 
rect 63 142 64 143 
rect 63 145 64 146 
rect 63 147 64 148 
rect 64 8 65 9 
rect 64 27 65 28 
rect 64 34 65 35 
rect 64 39 65 40 
rect 64 43 65 44 
rect 64 49 65 50 
rect 64 51 65 52 
rect 64 53 65 54 
rect 64 55 65 56 
rect 64 59 65 60 
rect 64 62 65 63 
rect 64 102 65 103 
rect 64 123 65 124 
rect 64 133 65 134 
rect 64 136 65 137 
rect 64 137 65 138 
rect 64 142 65 143 
rect 64 144 65 145 
rect 64 145 65 146 
rect 64 147 65 148 
rect 65 8 66 9 
rect 65 34 66 35 
rect 65 39 66 40 
rect 65 41 66 42 
rect 65 42 66 43 
rect 65 43 66 44 
rect 65 49 66 50 
rect 65 51 66 52 
rect 65 53 66 54 
rect 65 55 66 56 
rect 65 59 66 60 
rect 65 62 66 63 
rect 65 102 66 103 
rect 65 123 66 124 
rect 65 133 66 134 
rect 65 137 66 138 
rect 65 138 66 139 
rect 65 139 66 140 
rect 65 140 66 141 
rect 65 141 66 142 
rect 65 142 66 143 
rect 65 144 66 145 
rect 65 147 66 148 
rect 66 8 67 9 
rect 66 34 67 35 
rect 66 39 67 40 
rect 66 51 67 52 
rect 66 53 67 54 
rect 66 55 67 56 
rect 66 59 67 60 
rect 66 102 67 103 
rect 66 123 67 124 
rect 66 133 67 134 
rect 66 143 67 144 
rect 66 144 67 145 
rect 66 147 67 148 
rect 67 8 68 9 
rect 67 9 68 10 
rect 67 10 68 11 
rect 67 11 68 12 
rect 67 12 68 13 
rect 67 13 68 14 
rect 67 14 68 15 
rect 67 15 68 16 
rect 67 16 68 17 
rect 67 17 68 18 
rect 67 18 68 19 
rect 67 19 68 20 
rect 67 20 68 21 
rect 67 21 68 22 
rect 67 22 68 23 
rect 67 23 68 24 
rect 67 24 68 25 
rect 67 25 68 26 
rect 67 26 68 27 
rect 67 27 68 28 
rect 67 28 68 29 
rect 67 29 68 30 
rect 67 30 68 31 
rect 67 31 68 32 
rect 67 32 68 33 
rect 67 34 68 35 
rect 67 35 68 36 
rect 67 39 68 40 
rect 67 40 68 41 
rect 67 41 68 42 
rect 67 42 68 43 
rect 67 43 68 44 
rect 67 44 68 45 
rect 67 45 68 46 
rect 67 46 68 47 
rect 67 47 68 48 
rect 67 49 68 50 
rect 67 50 68 51 
rect 67 51 68 52 
rect 67 53 68 54 
rect 67 55 68 56 
rect 67 56 68 57 
rect 67 59 68 60 
rect 67 60 68 61 
rect 67 61 68 62 
rect 67 62 68 63 
rect 67 63 68 64 
rect 67 64 68 65 
rect 67 65 68 66 
rect 67 66 68 67 
rect 67 67 68 68 
rect 67 68 68 69 
rect 67 69 68 70 
rect 67 70 68 71 
rect 67 71 68 72 
rect 67 72 68 73 
rect 67 73 68 74 
rect 67 74 68 75 
rect 67 75 68 76 
rect 67 76 68 77 
rect 67 77 68 78 
rect 67 78 68 79 
rect 67 79 68 80 
rect 67 80 68 81 
rect 67 81 68 82 
rect 67 82 68 83 
rect 67 83 68 84 
rect 67 84 68 85 
rect 67 85 68 86 
rect 67 86 68 87 
rect 67 87 68 88 
rect 67 88 68 89 
rect 67 89 68 90 
rect 67 90 68 91 
rect 67 91 68 92 
rect 67 92 68 93 
rect 67 93 68 94 
rect 67 94 68 95 
rect 67 95 68 96 
rect 67 96 68 97 
rect 67 97 68 98 
rect 67 98 68 99 
rect 67 99 68 100 
rect 67 100 68 101 
rect 67 102 68 103 
rect 67 123 68 124 
rect 67 127 68 128 
rect 67 128 68 129 
rect 67 129 68 130 
rect 67 130 68 131 
rect 67 131 68 132 
rect 67 132 68 133 
rect 67 133 68 134 
rect 67 142 68 143 
rect 67 143 68 144 
rect 67 147 68 148 
rect 68 32 69 33 
rect 68 33 69 34 
rect 68 35 69 36 
rect 68 47 69 48 
rect 68 49 69 50 
rect 68 53 69 54 
rect 68 54 69 55 
rect 68 56 69 57 
rect 68 100 69 101 
rect 68 102 69 103 
rect 68 123 69 124 
rect 68 127 69 128 
rect 68 142 69 143 
rect 68 147 69 148 
rect 69 27 70 28 
rect 69 33 70 34 
rect 69 35 70 36 
rect 69 36 70 37 
rect 69 47 70 48 
rect 69 49 70 50 
rect 69 54 70 55 
rect 69 56 70 57 
rect 69 63 70 64 
rect 69 64 70 65 
rect 69 65 70 66 
rect 69 66 70 67 
rect 69 67 70 68 
rect 69 100 70 101 
rect 69 102 70 103 
rect 69 123 70 124 
rect 69 127 70 128 
rect 69 142 70 143 
rect 69 147 70 148 
rect 70 27 71 28 
rect 70 33 71 34 
rect 70 34 71 35 
rect 70 36 71 37 
rect 70 47 71 48 
rect 70 49 71 50 
rect 70 51 71 52 
rect 70 52 71 53 
rect 70 54 71 55 
rect 70 56 71 57 
rect 70 67 71 68 
rect 70 69 71 70 
rect 70 70 71 71 
rect 70 71 71 72 
rect 70 72 71 73 
rect 70 73 71 74 
rect 70 74 71 75 
rect 70 75 71 76 
rect 70 76 71 77 
rect 70 77 71 78 
rect 70 78 71 79 
rect 70 88 71 89 
rect 70 89 71 90 
rect 70 90 71 91 
rect 70 91 71 92 
rect 70 92 71 93 
rect 70 93 71 94 
rect 70 94 71 95 
rect 70 95 71 96 
rect 70 96 71 97 
rect 70 97 71 98 
rect 70 98 71 99 
rect 70 100 71 101 
rect 70 102 71 103 
rect 70 123 71 124 
rect 70 127 71 128 
rect 70 142 71 143 
rect 70 147 71 148 
rect 71 23 72 24 
rect 71 24 72 25 
rect 71 25 72 26 
rect 71 27 72 28 
rect 71 34 72 35 
rect 71 36 72 37 
rect 71 47 72 48 
rect 71 49 72 50 
rect 71 52 72 53 
rect 71 54 72 55 
rect 71 56 72 57 
rect 71 67 72 68 
rect 71 78 72 79 
rect 71 87 72 88 
rect 71 88 72 89 
rect 71 100 72 101 
rect 71 102 72 103 
rect 71 104 72 105 
rect 71 105 72 106 
rect 71 106 72 107 
rect 71 107 72 108 
rect 71 108 72 109 
rect 71 123 72 124 
rect 71 127 72 128 
rect 71 142 72 143 
rect 71 147 72 148 
rect 72 14 73 15 
rect 72 15 73 16 
rect 72 16 73 17 
rect 72 17 73 18 
rect 72 18 73 19 
rect 72 19 73 20 
rect 72 20 73 21 
rect 72 21 73 22 
rect 72 22 73 23 
rect 72 23 73 24 
rect 72 27 73 28 
rect 72 34 73 35 
rect 72 36 73 37 
rect 72 49 73 50 
rect 72 52 73 53 
rect 72 54 73 55 
rect 72 56 73 57 
rect 72 62 73 63 
rect 72 63 73 64 
rect 72 64 73 65 
rect 72 67 73 68 
rect 72 75 73 76 
rect 72 76 73 77 
rect 72 78 73 79 
rect 72 81 73 82 
rect 72 82 73 83 
rect 72 83 73 84 
rect 72 84 73 85 
rect 72 85 73 86 
rect 72 86 73 87 
rect 72 87 73 88 
rect 72 89 73 90 
rect 72 90 73 91 
rect 72 91 73 92 
rect 72 100 73 101 
rect 72 102 73 103 
rect 72 108 73 109 
rect 72 109 73 110 
rect 72 110 73 111 
rect 72 111 73 112 
rect 72 112 73 113 
rect 72 123 73 124 
rect 72 125 73 126 
rect 72 126 73 127 
rect 72 127 73 128 
rect 72 142 73 143 
rect 72 147 73 148 
rect 73 14 74 15 
rect 73 27 74 28 
rect 73 34 74 35 
rect 73 36 74 37 
rect 73 49 74 50 
rect 73 52 74 53 
rect 73 54 74 55 
rect 73 56 74 57 
rect 73 62 74 63 
rect 73 64 74 65 
rect 73 65 74 66 
rect 73 67 74 68 
rect 73 68 74 69 
rect 73 69 74 70 
rect 73 70 74 71 
rect 73 71 74 72 
rect 73 72 74 73 
rect 73 75 74 76 
rect 73 78 74 79 
rect 73 88 74 89 
rect 73 89 74 90 
rect 73 91 74 92 
rect 73 100 74 101 
rect 73 102 74 103 
rect 73 112 74 113 
rect 73 113 74 114 
rect 73 123 74 124 
rect 73 142 74 143 
rect 73 147 74 148 
rect 74 14 75 15 
rect 74 27 75 28 
rect 74 34 75 35 
rect 74 36 75 37 
rect 74 49 75 50 
rect 74 52 75 53 
rect 74 54 75 55 
rect 74 56 75 57 
rect 74 62 75 63 
rect 74 65 75 66 
rect 74 66 75 67 
rect 74 72 75 73 
rect 74 75 75 76 
rect 74 78 75 79 
rect 74 88 75 89 
rect 74 91 75 92 
rect 74 100 75 101 
rect 74 102 75 103 
rect 74 113 75 114 
rect 74 114 75 115 
rect 74 115 75 116 
rect 74 116 75 117 
rect 74 117 75 118 
rect 74 118 75 119 
rect 74 119 75 120 
rect 74 120 75 121 
rect 74 123 75 124 
rect 74 142 75 143 
rect 74 147 75 148 
rect 75 27 76 28 
rect 75 34 76 35 
rect 75 36 76 37 
rect 75 37 76 38 
rect 75 49 76 50 
rect 75 52 76 53 
rect 75 54 76 55 
rect 75 56 76 57 
rect 75 66 76 67 
rect 75 67 76 68 
rect 75 68 76 69 
rect 75 72 76 73 
rect 75 88 76 89 
rect 75 100 76 101 
rect 75 102 76 103 
rect 75 120 76 121 
rect 75 123 76 124 
rect 75 147 76 148 
rect 76 27 77 28 
rect 76 34 77 35 
rect 76 35 77 36 
rect 76 37 77 38 
rect 76 49 77 50 
rect 76 52 77 53 
rect 76 54 77 55 
rect 76 56 77 57 
rect 76 68 77 69 
rect 76 72 77 73 
rect 76 88 77 89 
rect 76 100 77 101 
rect 76 102 77 103 
rect 76 120 77 121 
rect 76 123 77 124 
rect 76 147 77 148 
rect 77 27 78 28 
rect 77 35 78 36 
rect 77 37 78 38 
rect 77 49 78 50 
rect 77 52 78 53 
rect 77 54 78 55 
rect 77 56 78 57 
rect 77 68 78 69 
rect 77 72 78 73 
rect 77 88 78 89 
rect 77 100 78 101 
rect 77 102 78 103 
rect 77 120 78 121 
rect 77 123 78 124 
rect 77 147 78 148 
rect 78 27 79 28 
rect 78 35 79 36 
rect 78 37 79 38 
rect 78 49 79 50 
rect 78 52 79 53 
rect 78 54 79 55 
rect 78 56 79 57 
rect 78 68 79 69 
rect 78 72 79 73 
rect 78 88 79 89 
rect 78 100 79 101 
rect 78 102 79 103 
rect 78 120 79 121 
rect 78 123 79 124 
rect 78 124 79 125 
rect 78 125 79 126 
rect 78 126 79 127 
rect 78 127 79 128 
rect 78 147 79 148 
rect 79 27 80 28 
rect 79 35 80 36 
rect 79 37 80 38 
rect 79 49 80 50 
rect 79 52 80 53 
rect 79 54 80 55 
rect 79 56 80 57 
rect 79 68 80 69 
rect 79 72 80 73 
rect 79 87 80 88 
rect 79 88 80 89 
rect 79 100 80 101 
rect 79 102 80 103 
rect 79 147 80 148 
rect 80 27 81 28 
rect 80 35 81 36 
rect 80 37 81 38 
rect 80 49 81 50 
rect 80 52 81 53 
rect 80 54 81 55 
rect 80 56 81 57 
rect 80 57 81 58 
rect 80 72 81 73 
rect 80 73 81 74 
rect 80 100 81 101 
rect 80 102 81 103 
rect 80 113 81 114 
rect 80 114 81 115 
rect 80 115 81 116 
rect 80 116 81 117 
rect 80 117 81 118 
rect 80 118 81 119 
rect 80 119 81 120 
rect 80 120 81 121 
rect 80 121 81 122 
rect 80 122 81 123 
rect 80 123 81 124 
rect 80 124 81 125 
rect 80 125 81 126 
rect 80 126 81 127 
rect 80 127 81 128 
rect 80 128 81 129 
rect 80 129 81 130 
rect 80 130 81 131 
rect 80 131 81 132 
rect 80 132 81 133 
rect 80 133 81 134 
rect 80 134 81 135 
rect 80 135 81 136 
rect 80 136 81 137 
rect 80 137 81 138 
rect 80 147 81 148 
rect 81 27 82 28 
rect 81 35 82 36 
rect 81 37 82 38 
rect 81 38 82 39 
rect 81 49 82 50 
rect 81 52 82 53 
rect 81 54 82 55 
rect 81 55 82 56 
rect 81 57 82 58 
rect 81 58 82 59 
rect 81 59 82 60 
rect 81 60 82 61 
rect 81 61 82 62 
rect 81 62 82 63 
rect 81 63 82 64 
rect 81 64 82 65 
rect 81 65 82 66 
rect 81 66 82 67 
rect 81 67 82 68 
rect 81 68 82 69 
rect 81 69 82 70 
rect 81 70 82 71 
rect 81 71 82 72 
rect 81 73 82 74 
rect 81 74 82 75 
rect 81 75 82 76 
rect 81 76 82 77 
rect 81 77 82 78 
rect 81 78 82 79 
rect 81 79 82 80 
rect 81 80 82 81 
rect 81 81 82 82 
rect 81 82 82 83 
rect 81 83 82 84 
rect 81 84 82 85 
rect 81 85 82 86 
rect 81 86 82 87 
rect 81 87 82 88 
rect 81 88 82 89 
rect 81 89 82 90 
rect 81 90 82 91 
rect 81 91 82 92 
rect 81 92 82 93 
rect 81 93 82 94 
rect 81 94 82 95 
rect 81 95 82 96 
rect 81 96 82 97 
rect 81 97 82 98 
rect 81 98 82 99 
rect 81 100 82 101 
rect 81 102 82 103 
rect 81 105 82 106 
rect 81 106 82 107 
rect 81 107 82 108 
rect 81 108 82 109 
rect 81 109 82 110 
rect 81 110 82 111 
rect 81 111 82 112 
rect 81 112 82 113 
rect 81 113 82 114 
rect 81 137 82 138 
rect 81 138 82 139 
rect 81 139 82 140 
rect 81 140 82 141 
rect 81 141 82 142 
rect 81 142 82 143 
rect 81 147 82 148 
rect 82 27 83 28 
rect 82 35 83 36 
rect 82 36 83 37 
rect 82 38 83 39 
rect 82 49 83 50 
rect 82 52 83 53 
rect 82 53 83 54 
rect 82 55 83 56 
rect 82 56 83 57 
rect 82 71 83 72 
rect 82 72 83 73 
rect 82 98 83 99 
rect 82 99 83 100 
rect 82 102 83 103 
rect 82 114 83 115 
rect 82 115 83 116 
rect 82 116 83 117 
rect 82 117 83 118 
rect 82 118 83 119 
rect 82 119 83 120 
rect 82 120 83 121 
rect 82 121 83 122 
rect 82 122 83 123 
rect 82 123 83 124 
rect 82 124 83 125 
rect 82 125 83 126 
rect 82 126 83 127 
rect 82 127 83 128 
rect 82 128 83 129 
rect 82 129 83 130 
rect 82 130 83 131 
rect 82 131 83 132 
rect 82 132 83 133 
rect 82 133 83 134 
rect 82 134 83 135 
rect 82 135 83 136 
rect 82 136 83 137 
rect 82 142 83 143 
rect 82 147 83 148 
rect 83 27 84 28 
rect 83 28 84 29 
rect 83 36 84 37 
rect 83 38 84 39 
rect 83 49 84 50 
rect 83 53 84 54 
rect 83 56 84 57 
rect 83 57 84 58 
rect 83 58 84 59 
rect 83 59 84 60 
rect 83 69 84 70 
rect 83 70 84 71 
rect 83 72 84 73 
rect 83 73 84 74 
rect 83 74 84 75 
rect 83 75 84 76 
rect 83 76 84 77 
rect 83 77 84 78 
rect 83 78 84 79 
rect 83 79 84 80 
rect 83 80 84 81 
rect 83 81 84 82 
rect 83 82 84 83 
rect 83 83 84 84 
rect 83 84 84 85 
rect 83 85 84 86 
rect 83 86 84 87 
rect 83 87 84 88 
rect 83 88 84 89 
rect 83 89 84 90 
rect 83 90 84 91 
rect 83 91 84 92 
rect 83 92 84 93 
rect 83 93 84 94 
rect 83 94 84 95 
rect 83 95 84 96 
rect 83 96 84 97 
rect 83 99 84 100 
rect 83 100 84 101 
rect 83 102 84 103 
rect 83 105 84 106 
rect 83 106 84 107 
rect 83 107 84 108 
rect 83 108 84 109 
rect 83 109 84 110 
rect 83 110 84 111 
rect 83 111 84 112 
rect 83 112 84 113 
rect 83 113 84 114 
rect 83 114 84 115 
rect 83 136 84 137 
rect 83 137 84 138 
rect 83 138 84 139 
rect 83 142 84 143 
rect 83 147 84 148 
rect 84 28 85 29 
rect 84 36 85 37 
rect 84 38 85 39 
rect 84 49 85 50 
rect 84 53 85 54 
rect 84 59 85 60 
rect 84 70 85 71 
rect 84 96 85 97 
rect 84 102 85 103 
rect 84 138 85 139 
rect 84 142 85 143 
rect 84 147 85 148 
rect 85 28 86 29 
rect 85 36 86 37 
rect 85 38 86 39 
rect 85 49 86 50 
rect 85 53 86 54 
rect 85 59 86 60 
rect 85 70 86 71 
rect 85 89 86 90 
rect 85 96 86 97 
rect 85 102 86 103 
rect 85 127 86 128 
rect 85 138 86 139 
rect 85 142 86 143 
rect 85 147 86 148 
rect 86 28 87 29 
rect 86 36 87 37 
rect 86 38 87 39 
rect 86 49 87 50 
rect 86 53 87 54 
rect 86 59 87 60 
rect 86 70 87 71 
rect 86 82 87 83 
rect 86 89 87 90 
rect 86 96 87 97 
rect 86 102 87 103 
rect 86 127 87 128 
rect 86 138 87 139 
rect 86 142 87 143 
rect 86 147 87 148 
rect 87 28 88 29 
rect 87 36 88 37 
rect 87 38 88 39 
rect 87 39 88 40 
rect 87 49 88 50 
rect 87 53 88 54 
rect 87 54 88 55 
rect 87 55 88 56 
rect 87 56 88 57 
rect 87 59 88 60 
rect 87 70 88 71 
rect 87 71 88 72 
rect 87 78 88 79 
rect 87 79 88 80 
rect 87 80 88 81 
rect 87 81 88 82 
rect 87 82 88 83 
rect 87 87 88 88 
rect 87 88 88 89 
rect 87 89 88 90 
rect 87 96 88 97 
rect 87 97 88 98 
rect 87 98 88 99 
rect 87 99 88 100 
rect 87 100 88 101 
rect 87 102 88 103 
rect 87 105 88 106 
rect 87 106 88 107 
rect 87 107 88 108 
rect 87 127 88 128 
rect 87 128 88 129 
rect 87 129 88 130 
rect 87 138 88 139 
rect 87 139 88 140 
rect 87 142 88 143 
rect 87 147 88 148 
rect 88 28 89 29 
rect 88 29 89 30 
rect 88 30 89 31 
rect 88 31 89 32 
rect 88 32 89 33 
rect 88 36 89 37 
rect 88 37 89 38 
rect 88 39 89 40 
rect 88 46 89 47 
rect 88 47 89 48 
rect 88 49 89 50 
rect 88 56 89 57 
rect 88 59 89 60 
rect 88 71 89 72 
rect 88 78 89 79 
rect 88 83 89 84 
rect 88 84 89 85 
rect 88 85 89 86 
rect 88 86 89 87 
rect 88 87 89 88 
rect 88 102 89 103 
rect 88 107 89 108 
rect 88 129 89 130 
rect 88 139 89 140 
rect 88 142 89 143 
rect 88 147 89 148 
rect 88 153 89 154 
rect 88 154 89 155 
rect 88 155 89 156 
rect 88 156 89 157 
rect 88 157 89 158 
rect 88 158 89 159 
rect 89 32 90 33 
rect 89 33 90 34 
rect 89 37 90 38 
rect 89 39 90 40 
rect 89 46 90 47 
rect 89 49 90 50 
rect 89 56 90 57 
rect 89 59 90 60 
rect 89 71 90 72 
rect 89 78 90 79 
rect 89 82 90 83 
rect 89 83 90 84 
rect 89 102 90 103 
rect 89 107 90 108 
rect 89 129 90 130 
rect 89 139 90 140 
rect 89 142 90 143 
rect 89 147 90 148 
rect 89 152 90 153 
rect 89 153 90 154 
rect 89 158 90 159 
rect 90 33 91 34 
rect 90 37 91 38 
rect 90 39 91 40 
rect 90 46 91 47 
rect 90 49 91 50 
rect 90 56 91 57 
rect 90 59 91 60 
rect 90 71 91 72 
rect 90 78 91 79 
rect 90 82 91 83 
rect 90 85 91 86 
rect 90 86 91 87 
rect 90 87 91 88 
rect 90 88 91 89 
rect 90 102 91 103 
rect 90 107 91 108 
rect 90 129 91 130 
rect 90 139 91 140 
rect 90 142 91 143 
rect 90 147 91 148 
rect 90 152 91 153 
rect 90 158 91 159 
rect 91 33 92 34 
rect 91 37 92 38 
rect 91 39 92 40 
rect 91 49 92 50 
rect 91 56 92 57 
rect 91 71 92 72 
rect 91 78 92 79 
rect 91 82 92 83 
rect 91 88 92 89 
rect 91 102 92 103 
rect 91 107 92 108 
rect 91 129 92 130 
rect 91 147 92 148 
rect 91 152 92 153 
rect 92 33 93 34 
rect 92 37 93 38 
rect 92 39 93 40 
rect 92 40 93 41 
rect 92 49 93 50 
rect 92 56 93 57 
rect 92 71 93 72 
rect 92 78 93 79 
rect 92 82 93 83 
rect 92 86 93 87 
rect 92 88 93 89 
rect 92 102 93 103 
rect 92 107 93 108 
rect 92 129 93 130 
rect 92 147 93 148 
rect 92 152 93 153 
rect 93 33 94 34 
rect 93 37 94 38 
rect 93 38 94 39 
rect 93 40 94 41 
rect 93 49 94 50 
rect 93 56 94 57 
rect 93 71 94 72 
rect 93 78 94 79 
rect 93 82 94 83 
rect 93 86 94 87 
rect 93 88 94 89 
rect 93 102 94 103 
rect 93 107 94 108 
rect 93 129 94 130 
rect 93 147 94 148 
rect 93 152 94 153 
rect 94 33 95 34 
rect 94 38 95 39 
rect 94 40 95 41 
rect 94 49 95 50 
rect 94 56 95 57 
rect 94 71 95 72 
rect 94 78 95 79 
rect 94 82 95 83 
rect 94 86 95 87 
rect 94 88 95 89 
rect 94 102 95 103 
rect 94 107 95 108 
rect 94 129 95 130 
rect 94 147 95 148 
rect 94 152 95 153 
rect 95 30 96 31 
rect 95 33 96 34 
rect 95 38 96 39 
rect 95 40 96 41 
rect 95 49 96 50 
rect 95 56 96 57 
rect 95 71 96 72 
rect 95 78 96 79 
rect 95 82 96 83 
rect 95 86 96 87 
rect 95 88 96 89 
rect 95 102 96 103 
rect 95 107 96 108 
rect 95 129 96 130 
rect 95 147 96 148 
rect 95 152 96 153 
rect 95 155 96 156 
rect 96 30 97 31 
rect 96 33 97 34 
rect 96 38 97 39 
rect 96 40 97 41 
rect 96 49 97 50 
rect 96 56 97 57 
rect 96 57 97 58 
rect 96 71 97 72 
rect 96 78 97 79 
rect 96 82 97 83 
rect 96 86 97 87 
rect 96 88 97 89 
rect 96 89 97 90 
rect 96 102 97 103 
rect 96 107 97 108 
rect 96 128 97 129 
rect 96 129 97 130 
rect 96 147 97 148 
rect 96 152 97 153 
rect 96 155 97 156 
rect 97 30 98 31 
rect 97 31 98 32 
rect 97 33 98 34 
rect 97 38 98 39 
rect 97 40 98 41 
rect 97 49 98 50 
rect 97 57 98 58 
rect 97 58 98 59 
rect 97 59 98 60 
rect 97 60 98 61 
rect 97 61 98 62 
rect 97 62 98 63 
rect 97 63 98 64 
rect 97 64 98 65 
rect 97 65 98 66 
rect 97 66 98 67 
rect 97 67 98 68 
rect 97 68 98 69 
rect 97 69 98 70 
rect 97 71 98 72 
rect 97 78 98 79 
rect 97 82 98 83 
rect 97 86 98 87 
rect 97 87 98 88 
rect 97 89 98 90 
rect 97 90 98 91 
rect 97 91 98 92 
rect 97 92 98 93 
rect 97 93 98 94 
rect 97 94 98 95 
rect 97 95 98 96 
rect 97 96 98 97 
rect 97 97 98 98 
rect 97 98 98 99 
rect 97 102 98 103 
rect 97 107 98 108 
rect 97 128 98 129 
rect 97 130 98 131 
rect 97 131 98 132 
rect 97 132 98 133 
rect 97 133 98 134 
rect 97 134 98 135 
rect 97 135 98 136 
rect 97 136 98 137 
rect 97 137 98 138 
rect 97 138 98 139 
rect 97 139 98 140 
rect 97 140 98 141 
rect 97 141 98 142 
rect 97 142 98 143 
rect 97 143 98 144 
rect 97 144 98 145 
rect 97 145 98 146 
rect 97 146 98 147 
rect 97 147 98 148 
rect 97 152 98 153 
rect 97 154 98 155 
rect 97 155 98 156 
rect 98 31 99 32 
rect 98 33 99 34 
rect 98 38 99 39 
rect 98 40 99 41 
rect 98 49 99 50 
rect 98 71 99 72 
rect 98 78 99 79 
rect 98 80 99 81 
rect 98 82 99 83 
rect 98 87 99 88 
rect 98 98 99 99 
rect 98 102 99 103 
rect 98 107 99 108 
rect 98 128 99 129 
rect 98 130 99 131 
rect 98 152 99 153 
rect 98 154 99 155 
rect 99 31 100 32 
rect 99 33 100 34 
rect 99 38 100 39 
rect 99 40 100 41 
rect 99 49 100 50 
rect 99 71 100 72 
rect 99 78 100 79 
rect 99 80 100 81 
rect 99 82 100 83 
rect 99 87 100 88 
rect 99 98 100 99 
rect 99 102 100 103 
rect 99 107 100 108 
rect 99 128 100 129 
rect 99 130 100 131 
rect 99 152 100 153 
rect 99 154 100 155 
rect 100 31 101 32 
rect 100 33 101 34 
rect 100 38 101 39 
rect 100 40 101 41 
rect 100 49 101 50 
rect 100 69 101 70 
rect 100 71 101 72 
rect 100 78 101 79 
rect 100 80 101 81 
rect 100 87 101 88 
rect 100 98 101 99 
rect 100 102 101 103 
rect 100 107 101 108 
rect 100 128 101 129 
rect 100 130 101 131 
rect 100 152 101 153 
rect 100 154 101 155 
rect 101 31 102 32 
rect 101 33 102 34 
rect 101 38 102 39 
rect 101 40 102 41 
rect 101 49 102 50 
rect 101 69 102 70 
rect 101 71 102 72 
rect 101 78 102 79 
rect 101 80 102 81 
rect 101 87 102 88 
rect 101 98 102 99 
rect 101 102 102 103 
rect 101 107 102 108 
rect 101 128 102 129 
rect 101 130 102 131 
rect 101 152 102 153 
rect 101 154 102 155 
rect 102 31 103 32 
rect 102 33 103 34 
rect 102 38 103 39 
rect 102 40 103 41 
rect 102 49 103 50 
rect 102 68 103 69 
rect 102 69 103 70 
rect 102 71 103 72 
rect 102 78 103 79 
rect 102 80 103 81 
rect 102 87 103 88 
rect 102 98 103 99 
rect 102 102 103 103 
rect 102 107 103 108 
rect 102 128 103 129 
rect 102 130 103 131 
rect 102 152 103 153 
rect 102 154 103 155 
rect 103 33 104 34 
rect 103 34 104 35 
rect 103 35 104 36 
rect 103 38 104 39 
rect 103 40 104 41 
rect 103 49 104 50 
rect 103 51 104 52 
rect 103 52 104 53 
rect 103 53 104 54 
rect 103 54 104 55 
rect 103 55 104 56 
rect 103 56 104 57 
rect 103 57 104 58 
rect 103 58 104 59 
rect 103 59 104 60 
rect 103 60 104 61 
rect 103 61 104 62 
rect 103 62 104 63 
rect 103 63 104 64 
rect 103 64 104 65 
rect 103 65 104 66 
rect 103 68 104 69 
rect 103 71 104 72 
rect 103 78 104 79 
rect 103 80 104 81 
rect 103 81 104 82 
rect 103 87 104 88 
rect 103 98 104 99 
rect 103 102 104 103 
rect 103 107 104 108 
rect 103 108 104 109 
rect 103 109 104 110 
rect 103 110 104 111 
rect 103 111 104 112 
rect 103 112 104 113 
rect 103 113 104 114 
rect 103 114 104 115 
rect 103 115 104 116 
rect 103 116 104 117 
rect 103 117 104 118 
rect 103 118 104 119 
rect 103 119 104 120 
rect 103 120 104 121 
rect 103 121 104 122 
rect 103 122 104 123 
rect 103 123 104 124 
rect 103 128 104 129 
rect 103 130 104 131 
rect 103 150 104 151 
rect 103 152 104 153 
rect 104 35 105 36 
rect 104 38 105 39 
rect 104 40 105 41 
rect 104 49 105 50 
rect 104 68 105 69 
rect 104 71 105 72 
rect 104 78 105 79 
rect 104 81 105 82 
rect 104 87 105 88 
rect 104 98 105 99 
rect 104 102 105 103 
rect 104 123 105 124 
rect 104 126 105 127 
rect 104 128 105 129 
rect 104 150 105 151 
rect 104 152 105 153 
rect 105 35 106 36 
rect 105 38 106 39 
rect 105 40 106 41 
rect 105 49 106 50 
rect 105 68 106 69 
rect 105 71 106 72 
rect 105 78 106 79 
rect 105 81 106 82 
rect 105 87 106 88 
rect 105 98 106 99 
rect 105 102 106 103 
rect 105 123 106 124 
rect 105 126 106 127 
rect 105 128 106 129 
rect 105 129 106 130 
rect 105 150 106 151 
rect 105 152 106 153 
rect 106 35 107 36 
rect 106 38 107 39 
rect 106 40 107 41 
rect 106 49 107 50 
rect 106 68 107 69 
rect 106 71 107 72 
rect 106 78 107 79 
rect 106 81 107 82 
rect 106 98 107 99 
rect 106 102 107 103 
rect 106 123 107 124 
rect 106 126 107 127 
rect 106 129 107 130 
rect 106 150 107 151 
rect 106 152 107 153 
rect 107 35 108 36 
rect 107 38 108 39 
rect 107 40 108 41 
rect 107 49 108 50 
rect 107 67 108 68 
rect 107 68 108 69 
rect 107 71 108 72 
rect 107 81 108 82 
rect 107 82 108 83 
rect 107 83 108 84 
rect 107 84 108 85 
rect 107 85 108 86 
rect 107 86 108 87 
rect 107 87 108 88 
rect 107 88 108 89 
rect 107 98 108 99 
rect 107 102 108 103 
rect 107 129 108 130 
rect 107 150 108 151 
rect 107 152 108 153 
rect 108 35 109 36 
rect 108 40 109 41 
rect 108 42 109 43 
rect 108 49 109 50 
rect 108 67 109 68 
rect 108 71 109 72 
rect 108 88 109 89 
rect 108 98 109 99 
rect 108 102 109 103 
rect 108 129 109 130 
rect 108 150 109 151 
rect 108 152 109 153 
rect 109 35 110 36 
rect 109 40 110 41 
rect 109 42 110 43 
rect 109 49 110 50 
rect 109 67 110 68 
rect 109 71 110 72 
rect 109 88 110 89 
rect 109 98 110 99 
rect 109 102 110 103 
rect 109 129 110 130 
rect 109 150 110 151 
rect 109 152 110 153 
rect 110 35 111 36 
rect 110 40 111 41 
rect 110 42 111 43 
rect 110 49 111 50 
rect 110 67 111 68 
rect 110 71 111 72 
rect 110 88 111 89 
rect 110 98 111 99 
rect 110 102 111 103 
rect 110 129 111 130 
rect 110 150 111 151 
rect 110 152 111 153 
rect 111 35 112 36 
rect 111 40 112 41 
rect 111 42 112 43 
rect 111 49 112 50 
rect 111 67 112 68 
rect 111 71 112 72 
rect 111 88 112 89 
rect 111 98 112 99 
rect 111 102 112 103 
rect 111 126 112 127 
rect 111 129 112 130 
rect 111 150 112 151 
rect 111 152 112 153 
rect 112 35 113 36 
rect 112 40 113 41 
rect 112 42 113 43 
rect 112 43 113 44 
rect 112 44 113 45 
rect 112 45 113 46 
rect 112 46 113 47 
rect 112 47 113 48 
rect 112 49 113 50 
rect 112 67 113 68 
rect 112 71 113 72 
rect 112 88 113 89 
rect 112 89 113 90 
rect 112 102 113 103 
rect 112 113 113 114 
rect 112 114 113 115 
rect 112 115 113 116 
rect 112 116 113 117 
rect 112 117 113 118 
rect 112 118 113 119 
rect 112 119 113 120 
rect 112 120 113 121 
rect 112 126 113 127 
rect 112 129 113 130 
rect 112 150 113 151 
rect 112 152 113 153 
rect 113 35 114 36 
rect 113 40 114 41 
rect 113 47 114 48 
rect 113 49 114 50 
rect 113 51 114 52 
rect 113 52 114 53 
rect 113 53 114 54 
rect 113 54 114 55 
rect 113 55 114 56 
rect 113 56 114 57 
rect 113 57 114 58 
rect 113 58 114 59 
rect 113 59 114 60 
rect 113 60 114 61 
rect 113 61 114 62 
rect 113 62 114 63 
rect 113 63 114 64 
rect 113 64 114 65 
rect 113 65 114 66 
rect 113 66 114 67 
rect 113 67 114 68 
rect 113 71 114 72 
rect 113 89 114 90 
rect 113 90 114 91 
rect 113 91 114 92 
rect 113 92 114 93 
rect 113 93 114 94 
rect 113 94 114 95 
rect 113 95 114 96 
rect 113 96 114 97 
rect 113 97 114 98 
rect 113 98 114 99 
rect 113 99 114 100 
rect 113 100 114 101 
rect 113 102 114 103 
rect 113 105 114 106 
rect 113 106 114 107 
rect 113 107 114 108 
rect 113 108 114 109 
rect 113 109 114 110 
rect 113 110 114 111 
rect 113 111 114 112 
rect 113 112 114 113 
rect 113 113 114 114 
rect 113 120 114 121 
rect 113 123 114 124 
rect 113 124 114 125 
rect 113 125 114 126 
rect 113 126 114 127 
rect 113 129 114 130 
rect 113 150 114 151 
rect 113 152 114 153 
rect 114 35 115 36 
rect 114 38 115 39 
rect 114 40 115 41 
rect 114 47 115 48 
rect 114 49 115 50 
rect 114 71 115 72 
rect 114 102 115 103 
rect 114 120 115 121 
rect 114 129 115 130 
rect 114 150 115 151 
rect 114 152 115 153 
rect 115 35 116 36 
rect 115 38 116 39 
rect 115 40 116 41 
rect 115 47 116 48 
rect 115 49 116 50 
rect 115 71 116 72 
rect 115 88 116 89 
rect 115 102 116 103 
rect 115 120 116 121 
rect 115 123 116 124 
rect 115 129 116 130 
rect 115 150 116 151 
rect 115 152 116 153 
rect 116 35 117 36 
rect 116 38 117 39 
rect 116 40 117 41 
rect 116 47 117 48 
rect 116 49 117 50 
rect 116 71 117 72 
rect 116 88 117 89 
rect 116 91 117 92 
rect 116 102 117 103 
rect 116 120 117 121 
rect 116 123 117 124 
rect 116 129 117 130 
rect 116 150 117 151 
rect 116 152 117 153 
rect 117 35 118 36 
rect 117 38 118 39 
rect 117 40 118 41 
rect 117 47 118 48 
rect 117 49 118 50 
rect 117 71 118 72 
rect 117 88 118 89 
rect 117 91 118 92 
rect 117 102 118 103 
rect 117 120 118 121 
rect 117 123 118 124 
rect 117 129 118 130 
rect 117 150 118 151 
rect 117 152 118 153 
rect 118 35 119 36 
rect 118 38 119 39 
rect 118 40 119 41 
rect 118 47 119 48 
rect 118 49 119 50 
rect 118 51 119 52 
rect 118 52 119 53 
rect 118 53 119 54 
rect 118 71 119 72 
rect 118 88 119 89 
rect 118 91 119 92 
rect 118 102 119 103 
rect 118 120 119 121 
rect 118 123 119 124 
rect 118 129 119 130 
rect 118 150 119 151 
rect 118 152 119 153 
rect 119 33 120 34 
rect 119 35 120 36 
rect 119 38 120 39 
rect 119 40 120 41 
rect 119 47 120 48 
rect 119 49 120 50 
rect 119 53 120 54 
rect 119 54 120 55 
rect 119 71 120 72 
rect 119 88 120 89 
rect 119 91 120 92 
rect 119 102 120 103 
rect 119 120 120 121 
rect 119 123 120 124 
rect 119 129 120 130 
rect 119 150 120 151 
rect 119 152 120 153 
rect 120 30 121 31 
rect 120 31 121 32 
rect 120 32 121 33 
rect 120 33 121 34 
rect 120 35 121 36 
rect 120 37 121 38 
rect 120 38 121 39 
rect 120 40 121 41 
rect 120 47 121 48 
rect 120 49 121 50 
rect 120 52 121 53 
rect 120 54 121 55 
rect 120 55 121 56 
rect 120 56 121 57 
rect 120 57 121 58 
rect 120 58 121 59 
rect 120 59 121 60 
rect 120 60 121 61 
rect 120 61 121 62 
rect 120 62 121 63 
rect 120 63 121 64 
rect 120 64 121 65 
rect 120 71 121 72 
rect 120 78 121 79 
rect 120 79 121 80 
rect 120 80 121 81 
rect 120 81 121 82 
rect 120 82 121 83 
rect 120 83 121 84 
rect 120 84 121 85 
rect 120 85 121 86 
rect 120 86 121 87 
rect 120 88 121 89 
rect 120 91 121 92 
rect 120 92 121 93 
rect 120 93 121 94 
rect 120 94 121 95 
rect 120 95 121 96 
rect 120 96 121 97 
rect 120 102 121 103 
rect 120 105 121 106 
rect 120 106 121 107 
rect 120 107 121 108 
rect 120 120 121 121 
rect 120 123 121 124 
rect 120 129 121 130 
rect 120 150 121 151 
rect 120 152 121 153 
rect 121 30 122 31 
rect 121 35 122 36 
rect 121 37 122 38 
rect 121 40 122 41 
rect 121 49 122 50 
rect 121 52 122 53 
rect 121 64 122 65 
rect 121 65 122 66 
rect 121 71 122 72 
rect 121 78 122 79 
rect 121 88 122 89 
rect 121 96 122 97 
rect 121 97 122 98 
rect 121 102 122 103 
rect 121 107 122 108 
rect 121 108 122 109 
rect 121 109 122 110 
rect 121 110 122 111 
rect 121 111 122 112 
rect 121 112 122 113 
rect 121 113 122 114 
rect 121 114 122 115 
rect 121 115 122 116 
rect 121 116 122 117 
rect 121 117 122 118 
rect 121 118 122 119 
rect 121 120 122 121 
rect 121 123 122 124 
rect 121 129 122 130 
rect 121 131 122 132 
rect 121 132 122 133 
rect 121 133 122 134 
rect 121 134 122 135 
rect 121 135 122 136 
rect 121 136 122 137 
rect 121 137 122 138 
rect 121 138 122 139 
rect 121 139 122 140 
rect 121 140 122 141 
rect 121 141 122 142 
rect 121 142 122 143 
rect 121 143 122 144 
rect 121 144 122 145 
rect 121 145 122 146 
rect 121 146 122 147 
rect 121 147 122 148 
rect 121 148 122 149 
rect 121 149 122 150 
rect 121 150 122 151 
rect 121 152 122 153 
rect 122 30 123 31 
rect 122 35 123 36 
rect 122 37 123 38 
rect 122 40 123 41 
rect 122 49 123 50 
rect 122 52 123 53 
rect 122 65 123 66 
rect 122 66 123 67 
rect 122 67 123 68 
rect 122 71 123 72 
rect 122 78 123 79 
rect 122 88 123 89 
rect 122 97 123 98 
rect 122 102 123 103 
rect 122 120 123 121 
rect 122 123 123 124 
rect 122 129 123 130 
rect 122 152 123 153 
rect 123 37 124 38 
rect 123 40 124 41 
rect 123 49 124 50 
rect 123 52 124 53 
rect 123 67 124 68 
rect 123 68 124 69 
rect 123 69 124 70 
rect 123 71 124 72 
rect 123 88 124 89 
rect 123 97 124 98 
rect 123 98 124 99 
rect 123 102 124 103 
rect 123 120 124 121 
rect 123 129 124 130 
rect 123 152 124 153 
rect 124 37 125 38 
rect 124 40 125 41 
rect 124 49 125 50 
rect 124 52 125 53 
rect 124 69 125 70 
rect 124 71 125 72 
rect 124 88 125 89 
rect 124 98 125 99 
rect 124 102 125 103 
rect 124 120 125 121 
rect 124 129 125 130 
rect 124 152 125 153 
rect 125 37 126 38 
rect 125 40 126 41 
rect 125 49 126 50 
rect 125 52 126 53 
rect 125 69 126 70 
rect 125 71 126 72 
rect 125 88 126 89 
rect 125 98 126 99 
rect 125 102 126 103 
rect 125 120 126 121 
rect 125 129 126 130 
rect 125 152 126 153 
rect 126 37 127 38 
rect 126 40 127 41 
rect 126 49 127 50 
rect 126 52 127 53 
rect 126 69 127 70 
rect 126 71 127 72 
rect 126 88 127 89 
rect 126 98 127 99 
rect 126 102 127 103 
rect 126 120 127 121 
rect 126 129 127 130 
rect 126 152 127 153 
rect 127 33 128 34 
rect 127 34 128 35 
rect 127 35 128 36 
rect 127 36 128 37 
rect 127 37 128 38 
rect 127 40 128 41 
rect 127 49 128 50 
rect 127 52 128 53 
rect 127 53 128 54 
rect 127 54 128 55 
rect 127 55 128 56 
rect 127 56 128 57 
rect 127 71 128 72 
rect 127 75 128 76 
rect 127 78 128 79 
rect 127 88 128 89 
rect 127 94 128 95 
rect 127 98 128 99 
rect 127 102 128 103 
rect 127 120 128 121 
rect 127 126 128 127 
rect 127 129 128 130 
rect 127 152 128 153 
rect 128 32 129 33 
rect 128 33 129 34 
rect 128 40 129 41 
rect 128 49 129 50 
rect 128 56 129 57 
rect 128 57 129 58 
rect 128 71 129 72 
rect 128 73 129 74 
rect 128 75 129 76 
rect 128 78 129 79 
rect 128 88 129 89 
rect 128 89 129 90 
rect 128 94 129 95 
rect 128 98 129 99 
rect 128 102 129 103 
rect 128 120 129 121 
rect 128 121 129 122 
rect 128 126 129 127 
rect 128 128 129 129 
rect 128 129 129 130 
rect 128 152 129 153 
rect 129 17 130 18 
rect 129 18 130 19 
rect 129 19 130 20 
rect 129 20 130 21 
rect 129 21 130 22 
rect 129 22 130 23 
rect 129 23 130 24 
rect 129 24 130 25 
rect 129 25 130 26 
rect 129 26 130 27 
rect 129 27 130 28 
rect 129 28 130 29 
rect 129 29 130 30 
rect 129 30 130 31 
rect 129 31 130 32 
rect 129 32 130 33 
rect 129 40 130 41 
rect 129 42 130 43 
rect 129 49 130 50 
rect 129 57 130 58 
rect 129 58 130 59 
rect 129 59 130 60 
rect 129 60 130 61 
rect 129 61 130 62 
rect 129 62 130 63 
rect 129 63 130 64 
rect 129 64 130 65 
rect 129 65 130 66 
rect 129 66 130 67 
rect 129 67 130 68 
rect 129 68 130 69 
rect 129 69 130 70 
rect 129 71 130 72 
rect 129 73 130 74 
rect 129 74 130 75 
rect 129 75 130 76 
rect 129 77 130 78 
rect 129 78 130 79 
rect 129 89 130 90 
rect 129 90 130 91 
rect 129 91 130 92 
rect 129 92 130 93 
rect 129 93 130 94 
rect 129 94 130 95 
rect 129 98 130 99 
rect 129 102 130 103 
rect 129 121 130 122 
rect 129 122 130 123 
rect 129 123 130 124 
rect 129 126 130 127 
rect 129 127 130 128 
rect 129 128 130 129 
rect 129 152 130 153 
rect 130 17 131 18 
rect 130 40 131 41 
rect 130 42 131 43 
rect 130 49 131 50 
rect 130 69 131 70 
rect 130 71 131 72 
rect 130 98 131 99 
rect 130 102 131 103 
rect 130 123 131 124 
rect 130 152 131 153 
rect 131 17 132 18 
rect 131 40 132 41 
rect 131 42 132 43 
rect 131 49 132 50 
rect 131 69 132 70 
rect 131 71 132 72 
rect 131 98 132 99 
rect 131 102 132 103 
rect 131 123 132 124 
rect 131 152 132 153 
rect 132 17 133 18 
rect 132 40 133 41 
rect 132 42 133 43 
rect 132 49 133 50 
rect 132 69 133 70 
rect 132 71 133 72 
rect 132 98 133 99 
rect 132 102 133 103 
rect 132 123 133 124 
rect 132 152 133 153 
rect 133 17 134 18 
rect 133 40 134 41 
rect 133 42 134 43 
rect 133 49 134 50 
rect 133 69 134 70 
rect 133 71 134 72 
rect 133 98 134 99 
rect 133 102 134 103 
rect 133 123 134 124 
rect 133 152 134 153 
rect 134 17 135 18 
rect 134 40 135 41 
rect 134 42 135 43 
rect 134 49 135 50 
rect 134 69 135 70 
rect 134 71 135 72 
rect 134 98 135 99 
rect 134 102 135 103 
rect 134 123 135 124 
rect 134 152 135 153 
rect 135 17 136 18 
rect 135 40 136 41 
rect 135 42 136 43 
rect 135 49 136 50 
rect 135 69 136 70 
rect 135 71 136 72 
rect 135 98 136 99 
rect 135 102 136 103 
rect 135 123 136 124 
rect 135 152 136 153 
rect 136 17 137 18 
rect 136 40 137 41 
rect 136 42 137 43 
rect 136 43 137 44 
rect 136 44 137 45 
rect 136 45 137 46 
rect 136 46 137 47 
rect 136 49 137 50 
rect 136 69 137 70 
rect 136 71 137 72 
rect 136 98 137 99 
rect 136 102 137 103 
rect 136 123 137 124 
rect 136 152 137 153 
rect 137 17 138 18 
rect 137 40 138 41 
rect 137 46 138 47 
rect 137 49 138 50 
rect 137 71 138 72 
rect 137 98 138 99 
rect 137 102 138 103 
rect 137 104 138 105 
rect 137 123 138 124 
rect 137 152 138 153 
rect 138 17 139 18 
rect 138 40 139 41 
rect 138 46 139 47 
rect 138 49 139 50 
rect 138 71 139 72 
rect 138 98 139 99 
rect 138 102 139 103 
rect 138 104 139 105 
rect 138 123 139 124 
rect 138 152 139 153 
rect 139 17 140 18 
rect 139 40 140 41 
rect 139 49 140 50 
rect 139 71 140 72 
rect 139 98 140 99 
rect 139 102 140 103 
rect 139 104 140 105 
rect 139 152 140 153 
rect 140 17 141 18 
rect 140 40 141 41 
rect 140 49 141 50 
rect 140 71 141 72 
rect 140 98 141 99 
rect 140 102 141 103 
rect 140 104 141 105 
rect 140 152 141 153 
rect 141 17 142 18 
rect 141 40 142 41 
rect 141 49 142 50 
rect 141 71 142 72 
rect 141 98 142 99 
rect 141 102 142 103 
rect 141 104 142 105 
rect 141 152 142 153 
rect 142 17 143 18 
rect 142 40 143 41 
rect 142 49 143 50 
rect 142 71 143 72 
rect 142 98 143 99 
rect 142 102 143 103 
rect 142 104 143 105 
rect 142 152 143 153 
rect 143 14 144 15 
rect 143 17 144 18 
rect 143 40 144 41 
rect 143 43 144 44 
rect 143 49 144 50 
rect 143 71 144 72 
rect 143 98 144 99 
rect 143 99 144 100 
rect 143 100 144 101 
rect 143 102 144 103 
rect 143 104 144 105 
rect 143 107 144 108 
rect 143 110 144 111 
rect 143 152 144 153 
rect 144 14 145 15 
rect 144 16 145 17 
rect 144 17 145 18 
rect 144 40 145 41 
rect 144 43 145 44 
rect 144 48 145 49 
rect 144 49 145 50 
rect 144 71 145 72 
rect 144 100 145 101 
rect 144 102 145 103 
rect 144 104 145 105 
rect 144 105 145 106 
rect 144 107 145 108 
rect 144 110 145 111 
rect 144 152 145 153 
rect 145 14 146 15 
rect 145 15 146 16 
rect 145 16 146 17 
rect 145 40 146 41 
rect 145 43 146 44 
rect 145 44 146 45 
rect 145 45 146 46 
rect 145 46 146 47 
rect 145 47 146 48 
rect 145 48 146 49 
rect 145 71 146 72 
rect 145 100 146 101 
rect 145 102 146 103 
rect 145 105 146 106 
rect 145 106 146 107 
rect 145 107 146 108 
rect 145 109 146 110 
rect 145 110 146 111 
rect 145 152 146 153 
rect 146 40 147 41 
rect 146 71 147 72 
rect 146 100 147 101 
rect 146 102 147 103 
rect 146 109 147 110 
rect 146 152 147 153 
rect 147 40 148 41 
rect 147 41 148 42 
rect 147 42 148 43 
rect 147 43 148 44 
rect 147 44 148 45 
rect 147 45 148 46 
rect 147 46 148 47 
rect 147 47 148 48 
rect 147 48 148 49 
rect 147 49 148 50 
rect 147 50 148 51 
rect 147 51 148 52 
rect 147 52 148 53 
rect 147 53 148 54 
rect 147 54 148 55 
rect 147 55 148 56 
rect 147 56 148 57 
rect 147 57 148 58 
rect 147 58 148 59 
rect 147 59 148 60 
rect 147 60 148 61 
rect 147 61 148 62 
rect 147 62 148 63 
rect 147 63 148 64 
rect 147 64 148 65 
rect 147 65 148 66 
rect 147 66 148 67 
rect 147 67 148 68 
rect 147 68 148 69 
rect 147 69 148 70 
rect 147 71 148 72 
rect 147 72 148 73 
rect 147 102 148 103 
rect 147 103 148 104 
rect 147 105 148 106 
rect 147 106 148 107 
rect 147 107 148 108 
rect 147 108 148 109 
rect 147 109 148 110 
rect 147 152 148 153 
rect 148 69 149 70 
rect 148 70 149 71 
rect 148 72 149 73 
rect 148 103 149 104 
rect 148 152 149 153 
rect 149 70 150 71 
rect 149 72 150 73 
rect 149 103 150 104 
rect 149 152 150 153 
rect 150 70 151 71 
rect 150 72 151 73 
rect 150 103 151 104 
rect 150 152 151 153 
rect 151 70 152 71 
rect 151 72 152 73 
rect 151 103 152 104 
rect 151 152 152 153 
rect 152 70 153 71 
rect 152 72 153 73 
rect 152 101 153 102 
rect 152 103 153 104 
rect 152 106 153 107 
rect 152 107 153 108 
rect 152 108 153 109 
rect 152 109 153 110 
rect 152 110 153 111 
rect 152 111 153 112 
rect 152 112 153 113 
rect 152 113 153 114 
rect 152 121 153 122 
rect 152 122 153 123 
rect 152 123 153 124 
rect 152 124 153 125 
rect 152 125 153 126 
rect 152 126 153 127 
rect 152 127 153 128 
rect 152 128 153 129 
rect 152 129 153 130 
rect 152 130 153 131 
rect 152 131 153 132 
rect 152 132 153 133 
rect 152 133 153 134 
rect 152 134 153 135 
rect 152 135 153 136 
rect 152 136 153 137 
rect 152 137 153 138 
rect 152 138 153 139 
rect 152 139 153 140 
rect 152 140 153 141 
rect 152 141 153 142 
rect 152 142 153 143 
rect 152 143 153 144 
rect 152 144 153 145 
rect 152 145 153 146 
rect 152 146 153 147 
rect 152 147 153 148 
rect 152 148 153 149 
rect 152 149 153 150 
rect 152 150 153 151 
rect 152 151 153 152 
rect 152 152 153 153 
rect 153 70 154 71 
rect 153 72 154 73 
rect 153 101 154 102 
rect 153 103 154 104 
rect 153 113 154 114 
rect 153 114 154 115 
rect 153 115 154 116 
rect 153 116 154 117 
rect 153 117 154 118 
rect 153 118 154 119 
rect 153 119 154 120 
rect 153 120 154 121 
rect 153 121 154 122 
rect 154 70 155 71 
rect 154 72 155 73 
rect 154 101 155 102 
rect 154 103 155 104 
rect 155 70 156 71 
rect 155 72 156 73 
rect 155 101 156 102 
rect 155 103 156 104 
rect 156 70 157 71 
rect 156 72 157 73 
rect 156 101 157 102 
rect 156 103 157 104 
rect 157 70 158 71 
rect 157 72 158 73 
rect 157 101 158 102 
rect 157 103 158 104 
rect 158 70 159 71 
rect 158 72 159 73 
rect 158 101 159 102 
rect 158 103 159 104 
rect 159 70 160 71 
rect 159 72 160 73 
rect 159 75 160 76 
rect 159 78 160 79 
rect 159 97 160 98 
rect 159 98 160 99 
rect 159 99 160 100 
rect 159 100 160 101 
rect 159 101 160 102 
rect 159 103 160 104 
rect 159 104 160 105 
rect 159 110 160 111 
rect 159 123 160 124 
rect 160 70 161 71 
rect 160 72 161 73 
rect 160 73 161 74 
rect 160 75 161 76 
rect 160 78 161 79 
rect 160 96 161 97 
rect 160 97 161 98 
rect 160 104 161 105 
rect 160 105 161 106 
rect 160 110 161 111 
rect 160 123 161 124 
rect 161 70 162 71 
rect 161 71 162 72 
rect 161 73 162 74 
rect 161 74 162 75 
rect 161 75 162 76 
rect 161 78 162 79 
rect 161 79 162 80 
rect 161 80 162 81 
rect 161 81 162 82 
rect 161 82 162 83 
rect 161 83 162 84 
rect 161 84 162 85 
rect 161 85 162 86 
rect 161 86 162 87 
rect 161 87 162 88 
rect 161 88 162 89 
rect 161 89 162 90 
rect 161 90 162 91 
rect 161 91 162 92 
rect 161 92 162 93 
rect 161 93 162 94 
rect 161 94 162 95 
rect 161 95 162 96 
rect 161 96 162 97 
rect 161 105 162 106 
rect 161 106 162 107 
rect 161 107 162 108 
rect 161 108 162 109 
rect 161 109 162 110 
rect 161 110 162 111 
rect 161 112 162 113 
rect 161 113 162 114 
rect 161 114 162 115 
rect 161 115 162 116 
rect 161 116 162 117 
rect 161 117 162 118 
rect 161 118 162 119 
rect 161 119 162 120 
rect 161 120 162 121 
rect 161 121 162 122 
rect 161 122 162 123 
rect 161 123 162 124 
rect 162 71 163 72 
rect 162 72 163 73 
rect 162 111 163 112 
rect 162 112 163 113 
rect 163 72 164 73 
rect 163 73 164 74 
rect 163 74 164 75 
rect 163 75 164 76 
rect 163 76 164 77 
rect 163 77 164 78 
rect 163 78 164 79 
rect 163 79 164 80 
rect 163 80 164 81 
rect 163 81 164 82 
rect 163 82 164 83 
rect 163 83 164 84 
rect 163 84 164 85 
rect 163 85 164 86 
rect 163 86 164 87 
rect 163 87 164 88 
rect 163 88 164 89 
rect 163 89 164 90 
rect 163 90 164 91 
rect 163 91 164 92 
rect 163 92 164 93 
rect 163 93 164 94 
rect 163 94 164 95 
rect 163 95 164 96 
rect 163 96 164 97 
rect 163 97 164 98 
rect 163 98 164 99 
rect 163 99 164 100 
rect 163 100 164 101 
rect 163 101 164 102 
rect 163 102 164 103 
rect 163 103 164 104 
rect 163 104 164 105 
rect 163 105 164 106 
rect 163 106 164 107 
rect 163 107 164 108 
rect 163 108 164 109 
rect 163 109 164 110 
rect 163 110 164 111 
rect 163 111 164 112 
<< metal2 >>
rect 13 98 14 99 
rect 13 99 14 100 
rect 13 100 14 101 
rect 13 101 14 102 
rect 16 56 17 57 
rect 16 100 17 101 
rect 17 56 18 57 
rect 17 100 18 101 
rect 18 56 19 57 
rect 18 100 19 101 
rect 19 56 20 57 
rect 19 100 20 101 
rect 21 45 22 46 
rect 21 46 22 47 
rect 21 47 22 48 
rect 21 48 22 49 
rect 23 46 24 47 
rect 23 47 24 48 
rect 23 48 24 49 
rect 23 49 24 50 
rect 30 150 31 151 
rect 31 117 32 118 
rect 31 150 32 151 
rect 32 117 33 118 
rect 32 119 33 120 
rect 32 150 33 151 
rect 33 117 34 118 
rect 33 119 34 120 
rect 33 150 34 151 
rect 34 117 35 118 
rect 34 119 35 120 
rect 35 117 36 118 
rect 35 119 36 120 
rect 36 117 37 118 
rect 36 119 37 120 
rect 37 117 38 118 
rect 37 119 38 120 
rect 38 117 39 118 
rect 39 135 40 136 
rect 39 136 40 137 
rect 39 137 40 138 
rect 39 138 40 139 
rect 39 139 40 140 
rect 39 140 40 141 
rect 39 141 40 142 
rect 39 142 40 143 
rect 39 143 40 144 
rect 39 144 40 145 
rect 39 145 40 146 
rect 39 146 40 147 
rect 39 147 40 148 
rect 39 148 40 149 
rect 39 149 40 150 
rect 39 150 40 151 
rect 39 151 40 152 
rect 39 152 40 153 
rect 39 153 40 154 
rect 39 154 40 155 
rect 39 155 40 156 
rect 39 156 40 157 
rect 40 32 41 33 
rect 40 33 41 34 
rect 40 34 41 35 
rect 40 35 41 36 
rect 40 36 41 37 
rect 40 37 41 38 
rect 40 38 41 39 
rect 40 39 41 40 
rect 40 40 41 41 
rect 40 41 41 42 
rect 40 42 41 43 
rect 40 43 41 44 
rect 40 44 41 45 
rect 40 45 41 46 
rect 40 46 41 47 
rect 40 47 41 48 
rect 40 48 41 49 
rect 40 49 41 50 
rect 40 50 41 51 
rect 40 51 41 52 
rect 40 52 41 53 
rect 40 53 41 54 
rect 40 54 41 55 
rect 40 55 41 56 
rect 40 56 41 57 
rect 40 57 41 58 
rect 40 58 41 59 
rect 40 59 41 60 
rect 40 80 41 81 
rect 40 81 41 82 
rect 40 82 41 83 
rect 40 83 41 84 
rect 40 112 41 113 
rect 40 113 41 114 
rect 40 114 41 115 
rect 40 115 41 116 
rect 40 116 41 117 
rect 40 121 41 122 
rect 40 122 41 123 
rect 40 123 41 124 
rect 40 124 41 125 
rect 40 125 41 126 
rect 40 126 41 127 
rect 40 127 41 128 
rect 40 128 41 129 
rect 40 129 41 130 
rect 40 130 41 131 
rect 40 131 41 132 
rect 40 132 41 133 
rect 40 133 41 134 
rect 40 134 41 135 
rect 40 135 41 136 
rect 41 116 42 117 
rect 41 117 42 118 
rect 41 118 42 119 
rect 41 119 42 120 
rect 41 120 42 121 
rect 41 121 42 122 
rect 41 136 42 137 
rect 41 137 42 138 
rect 41 149 42 150 
rect 41 150 42 151 
rect 41 151 42 152 
rect 41 152 42 153 
rect 42 134 43 135 
rect 42 135 43 136 
rect 42 136 43 137 
rect 47 51 48 52 
rect 47 52 48 53 
rect 47 53 48 54 
rect 47 54 48 55 
rect 47 55 48 56 
rect 47 56 48 57 
rect 47 97 48 98 
rect 48 97 49 98 
rect 49 34 50 35 
rect 49 35 50 36 
rect 49 36 50 37 
rect 49 37 50 38 
rect 49 38 50 39 
rect 49 39 50 40 
rect 49 40 50 41 
rect 49 41 50 42 
rect 49 42 50 43 
rect 49 74 50 75 
rect 49 75 50 76 
rect 49 76 50 77 
rect 49 77 50 78 
rect 49 78 50 79 
rect 49 79 50 80 
rect 49 80 50 81 
rect 49 81 50 82 
rect 49 82 50 83 
rect 49 83 50 84 
rect 49 84 50 85 
rect 49 85 50 86 
rect 49 86 50 87 
rect 49 87 50 88 
rect 49 88 50 89 
rect 49 89 50 90 
rect 49 90 50 91 
rect 49 91 50 92 
rect 49 92 50 93 
rect 49 93 50 94 
rect 49 94 50 95 
rect 49 95 50 96 
rect 49 96 50 97 
rect 49 97 50 98 
rect 50 34 51 35 
rect 51 34 52 35 
rect 51 48 52 49 
rect 51 49 52 50 
rect 51 50 52 51 
rect 51 51 52 52 
rect 51 52 52 53 
rect 51 53 52 54 
rect 51 54 52 55 
rect 51 55 52 56 
rect 51 56 52 57 
rect 51 57 52 58 
rect 52 34 53 35 
rect 52 79 53 80 
rect 52 80 53 81 
rect 52 81 53 82 
rect 52 82 53 83 
rect 52 83 53 84 
rect 52 84 53 85 
rect 52 85 53 86 
rect 52 86 53 87 
rect 52 87 53 88 
rect 52 88 53 89 
rect 52 89 53 90 
rect 52 90 53 91 
rect 52 91 53 92 
rect 52 92 53 93 
rect 52 93 53 94 
rect 53 34 54 35 
rect 53 38 54 39 
rect 53 39 54 40 
rect 53 40 54 41 
rect 53 41 54 42 
rect 53 42 54 43 
rect 53 43 54 44 
rect 53 44 54 45 
rect 53 45 54 46 
rect 53 46 54 47 
rect 53 47 54 48 
rect 53 48 54 49 
rect 53 49 54 50 
rect 53 50 54 51 
rect 53 51 54 52 
rect 53 52 54 53 
rect 53 53 54 54 
rect 53 54 54 55 
rect 53 55 54 56 
rect 53 56 54 57 
rect 53 57 54 58 
rect 53 58 54 59 
rect 53 59 54 60 
rect 53 60 54 61 
rect 53 61 54 62 
rect 53 62 54 63 
rect 53 63 54 64 
rect 53 64 54 65 
rect 53 65 54 66 
rect 53 66 54 67 
rect 53 67 54 68 
rect 53 68 54 69 
rect 53 69 54 70 
rect 53 70 54 71 
rect 53 71 54 72 
rect 53 72 54 73 
rect 53 73 54 74 
rect 53 74 54 75 
rect 53 75 54 76 
rect 53 76 54 77 
rect 53 77 54 78 
rect 53 78 54 79 
rect 53 79 54 80 
rect 53 122 54 123 
rect 53 123 54 124 
rect 53 124 54 125 
rect 53 125 54 126 
rect 54 80 55 81 
rect 54 81 55 82 
rect 54 82 55 83 
rect 54 83 55 84 
rect 54 84 55 85 
rect 54 85 55 86 
rect 54 86 55 87 
rect 54 87 55 88 
rect 54 88 55 89 
rect 54 89 55 90 
rect 54 90 55 91 
rect 54 91 55 92 
rect 54 92 55 93 
rect 54 134 55 135 
rect 54 135 55 136 
rect 54 136 55 137 
rect 54 137 55 138 
rect 55 31 56 32 
rect 55 32 56 33 
rect 55 33 56 34 
rect 55 34 56 35 
rect 55 35 56 36 
rect 55 36 56 37 
rect 55 37 56 38 
rect 55 38 56 39 
rect 55 39 56 40 
rect 55 40 56 41 
rect 55 41 56 42 
rect 55 42 56 43 
rect 55 43 56 44 
rect 55 44 56 45 
rect 55 45 56 46 
rect 55 46 56 47 
rect 55 47 56 48 
rect 55 48 56 49 
rect 55 49 56 50 
rect 55 50 56 51 
rect 55 51 56 52 
rect 55 52 56 53 
rect 55 53 56 54 
rect 55 54 56 55 
rect 55 55 56 56 
rect 55 56 56 57 
rect 55 57 56 58 
rect 55 121 56 122 
rect 55 122 56 123 
rect 55 123 56 124 
rect 55 124 56 125 
rect 56 88 57 89 
rect 56 89 57 90 
rect 56 90 57 91 
rect 56 134 57 135 
rect 56 135 57 136 
rect 56 136 57 137 
rect 56 137 57 138 
rect 57 33 58 34 
rect 57 34 58 35 
rect 57 35 58 36 
rect 57 36 58 37 
rect 57 37 58 38 
rect 57 38 58 39 
rect 57 39 58 40 
rect 57 40 58 41 
rect 57 82 58 83 
rect 57 88 58 89 
rect 58 40 59 41 
rect 58 82 59 83 
rect 58 88 59 89 
rect 59 40 60 41 
rect 59 82 60 83 
rect 59 88 60 89 
rect 60 40 61 41 
rect 60 82 61 83 
rect 60 88 61 89 
rect 61 40 62 41 
rect 61 82 62 83 
rect 61 88 62 89 
rect 62 40 63 41 
rect 62 82 63 83 
rect 62 88 63 89 
rect 63 35 64 36 
rect 63 36 64 37 
rect 63 40 64 41 
rect 63 82 64 83 
rect 63 88 64 89 
rect 64 35 65 36 
rect 64 40 65 41 
rect 64 41 65 42 
rect 64 82 65 83 
rect 64 88 65 89 
rect 65 27 66 28 
rect 65 35 66 36 
rect 65 82 66 83 
rect 65 88 66 89 
rect 66 27 67 28 
rect 66 35 67 36 
rect 66 49 67 50 
rect 66 62 67 63 
rect 66 82 67 83 
rect 66 88 67 89 
rect 67 27 68 28 
rect 67 35 68 36 
rect 67 49 68 50 
rect 67 50 68 51 
rect 67 62 68 63 
rect 67 82 68 83 
rect 67 88 68 89 
rect 68 27 69 28 
rect 68 35 69 36 
rect 68 50 69 51 
rect 68 51 69 52 
rect 68 62 69 63 
rect 68 82 69 83 
rect 68 88 69 89 
rect 69 35 70 36 
rect 69 51 70 52 
rect 69 62 70 63 
rect 69 82 70 83 
rect 69 88 70 89 
rect 70 35 71 36 
rect 70 82 71 83 
rect 70 88 71 89 
rect 70 99 71 100 
rect 70 100 71 101 
rect 70 101 71 102 
rect 70 102 71 103 
rect 70 103 71 104 
rect 70 104 71 105 
rect 71 26 72 27 
rect 71 27 72 28 
rect 71 28 72 29 
rect 71 29 72 30 
rect 71 30 72 31 
rect 71 31 72 32 
rect 71 32 72 33 
rect 71 33 72 34 
rect 71 34 72 35 
rect 71 35 72 36 
rect 71 48 72 49 
rect 71 49 72 50 
rect 71 50 72 51 
rect 71 51 72 52 
rect 71 52 72 53 
rect 71 53 72 54 
rect 71 54 72 55 
rect 71 55 72 56 
rect 71 56 72 57 
rect 71 57 72 58 
rect 71 58 72 59 
rect 71 59 72 60 
rect 71 60 72 61 
rect 71 61 72 62 
rect 71 62 72 63 
rect 71 63 72 64 
rect 71 64 72 65 
rect 71 65 72 66 
rect 71 66 72 67 
rect 71 67 72 68 
rect 71 68 72 69 
rect 71 69 72 70 
rect 71 82 72 83 
rect 71 88 72 89 
rect 72 77 73 78 
rect 72 78 73 79 
rect 72 79 73 80 
rect 72 80 73 81 
rect 72 82 73 83 
rect 72 88 73 89 
rect 72 97 73 98 
rect 72 98 73 99 
rect 72 99 73 100 
rect 72 100 73 101 
rect 72 101 73 102 
rect 72 102 73 103 
rect 72 103 73 104 
rect 72 104 73 105 
rect 72 105 73 106 
rect 72 106 73 107 
rect 72 107 73 108 
rect 72 108 73 109 
rect 72 109 73 110 
rect 72 110 73 111 
rect 72 111 73 112 
rect 72 112 73 113 
rect 72 113 73 114 
rect 72 114 73 115 
rect 72 115 73 116 
rect 72 116 73 117 
rect 72 117 73 118 
rect 72 118 73 119 
rect 72 119 73 120 
rect 72 120 73 121 
rect 72 121 73 122 
rect 72 122 73 123 
rect 72 123 73 124 
rect 72 124 73 125 
rect 73 82 74 83 
rect 73 88 74 89 
rect 73 97 74 98 
rect 74 82 75 83 
rect 74 88 75 89 
rect 74 97 75 98 
rect 75 82 76 83 
rect 75 88 76 89 
rect 75 97 76 98 
rect 76 82 77 83 
rect 76 88 77 89 
rect 76 97 77 98 
rect 77 82 78 83 
rect 77 88 78 89 
rect 77 97 78 98 
rect 78 82 79 83 
rect 78 88 79 89 
rect 78 97 79 98 
rect 79 82 80 83 
rect 79 86 80 87 
rect 79 88 80 89 
rect 79 97 80 98 
rect 79 120 80 121 
rect 79 127 80 128 
rect 80 68 81 69 
rect 80 82 81 83 
rect 80 86 81 87 
rect 80 88 81 89 
rect 80 96 81 97 
rect 80 97 81 98 
rect 80 120 81 121 
rect 80 127 81 128 
rect 81 68 82 69 
rect 81 82 82 83 
rect 81 86 82 87 
rect 81 88 82 89 
rect 81 90 82 91 
rect 81 91 82 92 
rect 81 92 82 93 
rect 81 93 82 94 
rect 81 94 82 95 
rect 81 95 82 96 
rect 81 96 82 97 
rect 81 101 82 102 
rect 81 102 82 103 
rect 81 103 82 104 
rect 81 104 82 105 
rect 81 120 82 121 
rect 81 127 82 128 
rect 82 68 83 69 
rect 82 82 83 83 
rect 82 86 83 87 
rect 82 88 83 89 
rect 82 90 83 91 
rect 82 120 83 121 
rect 82 127 83 128 
rect 83 68 84 69 
rect 83 82 84 83 
rect 83 86 84 87 
rect 83 88 84 89 
rect 83 90 84 91 
rect 83 101 84 102 
rect 83 102 84 103 
rect 83 103 84 104 
rect 83 104 84 105 
rect 83 120 84 121 
rect 83 127 84 128 
rect 84 82 85 83 
rect 84 86 85 87 
rect 84 88 85 89 
rect 84 90 85 91 
rect 84 120 85 121 
rect 84 127 85 128 
rect 85 82 86 83 
rect 85 86 86 87 
rect 85 88 86 89 
rect 85 90 86 91 
rect 85 120 86 121 
rect 86 86 87 87 
rect 86 88 87 89 
rect 86 120 87 121 
rect 87 86 88 87 
rect 87 88 88 89 
rect 87 101 88 102 
rect 87 102 88 103 
rect 87 103 88 104 
rect 87 104 88 105 
rect 87 120 88 121 
rect 88 48 89 49 
rect 88 49 89 50 
rect 88 50 89 51 
rect 88 51 89 52 
rect 88 52 89 53 
rect 88 53 89 54 
rect 88 54 89 55 
rect 88 55 89 56 
rect 88 56 89 57 
rect 88 57 89 58 
rect 88 58 89 59 
rect 88 59 89 60 
rect 88 60 89 61 
rect 88 61 89 62 
rect 88 62 89 63 
rect 88 63 89 64 
rect 88 64 89 65 
rect 88 65 89 66 
rect 88 66 89 67 
rect 88 67 89 68 
rect 88 68 89 69 
rect 88 86 89 87 
rect 88 88 89 89 
rect 88 120 89 121 
rect 89 68 90 69 
rect 89 86 90 87 
rect 89 88 90 89 
rect 89 120 90 121 
rect 90 68 91 69 
rect 90 69 91 70 
rect 90 70 91 71 
rect 90 71 91 72 
rect 90 72 91 73 
rect 90 73 91 74 
rect 90 74 91 75 
rect 90 75 91 76 
rect 90 76 91 77 
rect 90 77 91 78 
rect 90 78 91 79 
rect 90 79 91 80 
rect 90 80 91 81 
rect 90 81 91 82 
rect 90 82 91 83 
rect 90 83 91 84 
rect 90 84 91 85 
rect 90 86 91 87 
rect 90 88 91 89 
rect 90 120 91 121 
rect 91 86 92 87 
rect 91 88 92 89 
rect 91 120 92 121 
rect 92 88 93 89 
rect 92 120 93 121 
rect 93 88 94 89 
rect 93 120 94 121 
rect 94 88 95 89 
rect 94 120 95 121 
rect 95 88 96 89 
rect 95 120 96 121 
rect 96 88 97 89 
rect 96 120 97 121 
rect 97 70 98 71 
rect 97 71 98 72 
rect 97 72 98 73 
rect 97 73 98 74 
rect 97 74 98 75 
rect 97 75 98 76 
rect 97 76 98 77 
rect 97 77 98 78 
rect 97 78 98 79 
rect 97 79 98 80 
rect 97 80 98 81 
rect 97 88 98 89 
rect 97 120 98 121 
rect 98 88 99 89 
rect 98 120 99 121 
rect 99 69 100 70 
rect 99 70 100 71 
rect 99 71 100 72 
rect 99 72 100 73 
rect 99 73 100 74 
rect 99 74 100 75 
rect 99 75 100 76 
rect 99 76 100 77 
rect 99 77 100 78 
rect 99 78 100 79 
rect 99 79 100 80 
rect 99 80 100 81 
rect 99 81 100 82 
rect 99 88 100 89 
rect 99 120 100 121 
rect 100 88 101 89 
rect 100 120 101 121 
rect 101 88 102 89 
rect 101 120 102 121 
rect 102 88 103 89 
rect 102 120 103 121 
rect 103 31 104 32 
rect 103 32 104 33 
rect 103 33 104 34 
rect 103 34 104 35 
rect 103 35 104 36 
rect 103 36 104 37 
rect 103 37 104 38 
rect 103 38 104 39 
rect 103 39 104 40 
rect 103 40 104 41 
rect 103 41 104 42 
rect 103 42 104 43 
rect 103 43 104 44 
rect 103 44 104 45 
rect 103 45 104 46 
rect 103 46 104 47 
rect 103 47 104 48 
rect 103 48 104 49 
rect 103 49 104 50 
rect 103 50 104 51 
rect 103 66 104 67 
rect 103 67 104 68 
rect 103 88 104 89 
rect 103 120 104 121 
rect 103 126 104 127 
rect 103 127 104 128 
rect 103 128 104 129 
rect 103 129 104 130 
rect 103 151 104 152 
rect 103 152 104 153 
rect 103 153 104 154 
rect 103 154 104 155 
rect 104 67 105 68 
rect 104 88 105 89 
rect 104 120 105 121 
rect 105 67 106 68 
rect 105 86 106 87 
rect 105 88 106 89 
rect 105 120 106 121 
rect 106 67 107 68 
rect 106 86 107 87 
rect 106 88 107 89 
rect 106 120 107 121 
rect 107 39 108 40 
rect 107 40 108 41 
rect 107 41 108 42 
rect 107 42 108 43 
rect 107 67 108 68 
rect 107 86 108 87 
rect 107 88 108 89 
rect 107 120 108 121 
rect 108 67 109 68 
rect 108 86 109 87 
rect 108 88 109 89 
rect 108 120 109 121 
rect 109 67 110 68 
rect 109 86 110 87 
rect 109 88 110 89 
rect 109 120 110 121 
rect 110 67 111 68 
rect 110 86 111 87 
rect 110 88 111 89 
rect 110 120 111 121 
rect 111 67 112 68 
rect 111 86 112 87 
rect 111 88 112 89 
rect 111 120 112 121 
rect 112 67 113 68 
rect 112 86 113 87 
rect 112 88 113 89 
rect 112 98 113 99 
rect 112 120 113 121 
rect 112 121 113 122 
rect 113 38 114 39 
rect 113 39 114 40 
rect 113 40 114 41 
rect 113 41 114 42 
rect 113 42 114 43 
rect 113 43 114 44 
rect 113 44 114 45 
rect 113 45 114 46 
rect 113 46 114 47 
rect 113 47 114 48 
rect 113 48 114 49 
rect 113 49 114 50 
rect 113 50 114 51 
rect 113 67 114 68 
rect 113 86 114 87 
rect 113 88 114 89 
rect 113 98 114 99 
rect 113 101 114 102 
rect 113 102 114 103 
rect 113 103 114 104 
rect 113 104 114 105 
rect 113 121 114 122 
rect 113 122 114 123 
rect 114 67 115 68 
rect 114 86 115 87 
rect 114 88 115 89 
rect 114 98 115 99 
rect 114 99 115 100 
rect 115 67 116 68 
rect 115 86 116 87 
rect 115 87 116 88 
rect 115 99 116 100 
rect 115 100 116 101 
rect 115 101 116 102 
rect 115 102 116 103 
rect 115 103 116 104 
rect 115 104 116 105 
rect 115 105 116 106 
rect 115 106 116 107 
rect 115 107 116 108 
rect 115 108 116 109 
rect 115 109 116 110 
rect 115 110 116 111 
rect 115 111 116 112 
rect 115 112 116 113 
rect 115 113 116 114 
rect 115 114 116 115 
rect 115 115 116 116 
rect 115 116 116 117 
rect 115 117 116 118 
rect 115 118 116 119 
rect 115 119 116 120 
rect 115 120 116 121 
rect 115 121 116 122 
rect 115 122 116 123 
rect 116 67 117 68 
rect 116 87 117 88 
rect 116 88 117 89 
rect 116 89 117 90 
rect 116 90 117 91 
rect 117 67 118 68 
rect 118 33 119 34 
rect 118 34 119 35 
rect 118 35 119 36 
rect 118 36 119 37 
rect 118 37 119 38 
rect 118 38 119 39 
rect 118 39 119 40 
rect 118 40 119 41 
rect 118 41 119 42 
rect 118 42 119 43 
rect 118 43 119 44 
rect 118 44 119 45 
rect 118 45 119 46 
rect 118 46 119 47 
rect 118 47 119 48 
rect 118 48 119 49 
rect 118 49 119 50 
rect 118 50 119 51 
rect 118 67 119 68 
rect 119 67 120 68 
rect 120 48 121 49 
rect 120 49 121 50 
rect 120 50 121 51 
rect 120 51 121 52 
rect 120 67 121 68 
rect 120 87 121 88 
rect 120 88 121 89 
rect 120 89 121 90 
rect 120 90 121 91 
rect 120 91 121 92 
rect 120 92 121 93 
rect 120 93 121 94 
rect 120 94 121 95 
rect 120 95 121 96 
rect 120 96 121 97 
rect 120 97 121 98 
rect 120 98 121 99 
rect 120 99 121 100 
rect 120 100 121 101 
rect 120 101 121 102 
rect 120 102 121 103 
rect 120 103 121 104 
rect 120 104 121 105 
rect 120 121 121 122 
rect 120 122 121 123 
rect 120 123 121 124 
rect 120 124 121 125 
rect 120 125 121 126 
rect 120 126 121 127 
rect 120 127 121 128 
rect 120 128 121 129 
rect 120 129 121 130 
rect 120 130 121 131 
rect 120 131 121 132 
rect 121 67 122 68 
rect 121 119 122 120 
rect 121 120 122 121 
rect 121 121 122 122 
rect 122 67 123 68 
rect 123 35 124 36 
rect 123 36 124 37 
rect 123 67 124 68 
rect 124 36 125 37 
rect 124 67 125 68 
rect 125 36 126 37 
rect 125 67 126 68 
rect 126 36 127 37 
rect 126 67 127 68 
rect 127 36 128 37 
rect 127 67 128 68 
rect 127 69 128 70 
rect 127 70 128 71 
rect 127 71 128 72 
rect 127 72 128 73 
rect 128 36 129 37 
rect 128 67 129 68 
rect 128 68 129 69 
rect 128 72 129 73 
rect 129 36 130 37 
rect 129 37 130 38 
rect 129 38 130 39 
rect 129 39 130 40 
rect 129 40 130 41 
rect 129 41 130 42 
rect 129 68 130 69 
rect 129 69 130 70 
rect 129 70 130 71 
rect 129 71 130 72 
rect 129 74 130 75 
rect 129 75 130 76 
rect 129 76 130 77 
rect 130 71 131 72 
rect 130 72 131 73 
rect 130 73 131 74 
rect 130 74 131 75 
rect 136 70 137 71 
rect 136 71 137 72 
rect 136 72 137 73 
rect 136 73 137 74 
rect 136 74 137 75 
rect 136 75 137 76 
rect 136 76 137 77 
rect 136 77 137 78 
rect 136 78 137 79 
rect 136 79 137 80 
rect 136 80 137 81 
rect 136 81 137 82 
rect 136 82 137 83 
rect 136 83 137 84 
rect 136 84 137 85 
rect 136 85 137 86 
rect 136 86 137 87 
rect 136 87 137 88 
rect 136 88 137 89 
rect 136 89 137 90 
rect 136 90 137 91 
rect 136 91 137 92 
rect 136 92 137 93 
rect 136 93 137 94 
rect 136 94 137 95 
rect 136 95 137 96 
rect 136 96 137 97 
rect 136 97 137 98 
rect 136 98 137 99 
rect 136 99 137 100 
rect 136 100 137 101 
rect 136 101 137 102 
rect 136 102 137 103 
rect 136 103 137 104 
rect 136 104 137 105 
rect 147 100 148 101 
rect 147 101 148 102 
rect 147 102 148 103 
rect 147 103 148 104 
rect 147 104 148 105 
rect 152 102 153 103 
rect 152 103 153 104 
rect 152 104 153 105 
rect 152 105 153 106 
<< m2contact >>
rect 13 98 14 99 
rect 19 56 20 57 
rect 19 100 20 101 
rect 21 45 22 46 
rect 23 49 24 50 
rect 31 117 32 118 
rect 33 150 34 151 
rect 37 119 38 120 
rect 39 156 40 157 
rect 40 32 41 33 
rect 40 80 41 81 
rect 41 137 42 138 
rect 41 149 42 150 
rect 47 51 48 52 
rect 47 97 48 98 
rect 51 57 52 58 
rect 52 93 53 94 
rect 53 34 54 35 
rect 53 125 54 126 
rect 54 80 55 81 
rect 54 134 55 135 
rect 55 57 56 58 
rect 55 121 56 122 
rect 56 134 57 135 
rect 63 36 64 37 
rect 64 41 65 42 
rect 65 27 66 28 
rect 69 51 70 52 
rect 69 62 70 63 
rect 70 104 71 105 
rect 71 69 72 70 
rect 72 80 73 81 
rect 79 86 80 87 
rect 81 104 82 105 
rect 83 68 84 69 
rect 83 104 84 105 
rect 84 127 85 128 
rect 85 82 86 83 
rect 85 90 86 91 
rect 87 104 88 105 
rect 90 84 91 85 
rect 97 80 98 81 
rect 99 69 100 70 
rect 103 31 104 32 
rect 103 66 104 67 
rect 103 126 104 127 
rect 103 154 104 155 
rect 105 86 106 87 
rect 107 42 108 43 
rect 113 38 114 39 
rect 113 104 114 105 
rect 113 122 114 123 
rect 114 88 115 89 
rect 115 122 116 123 
rect 118 33 119 34 
rect 120 51 121 52 
rect 120 104 121 105 
rect 120 131 121 132 
rect 123 35 124 36 
rect 127 69 128 70 
rect 136 104 137 105 
rect 147 100 148 101 
rect 152 105 153 106 
rect 13 102 14 103 
rect 15 56 16 57 
rect 15 100 16 101 
rect 21 49 22 50 
rect 23 45 24 46 
rect 29 150 30 151 
rect 31 119 32 120 
rect 39 117 40 118 
rect 40 60 41 61 
rect 40 84 41 85 
rect 40 111 41 112 
rect 41 153 42 154 
rect 42 133 43 134 
rect 47 57 48 58 
rect 49 43 50 44 
rect 49 73 50 74 
rect 51 47 52 48 
rect 53 37 54 38 
rect 53 121 54 122 
rect 54 93 55 94 
rect 54 138 55 139 
rect 55 30 56 31 
rect 55 125 56 126 
rect 56 82 57 83 
rect 56 91 57 92 
rect 56 138 57 139 
rect 57 32 58 33 
rect 65 49 66 50 
rect 65 62 66 63 
rect 69 27 70 28 
rect 70 98 71 99 
rect 71 25 72 26 
rect 71 47 72 48 
rect 72 76 73 77 
rect 72 125 73 126 
rect 78 120 79 121 
rect 78 127 79 128 
rect 79 68 80 69 
rect 81 100 82 101 
rect 83 100 84 101 
rect 87 100 88 101 
rect 88 47 89 48 
rect 92 86 93 87 
rect 97 69 98 70 
rect 99 82 100 83 
rect 103 51 104 52 
rect 103 130 104 131 
rect 103 150 104 151 
rect 107 38 108 39 
rect 111 98 112 99 
rect 113 51 114 52 
rect 113 100 114 101 
rect 116 91 117 92 
rect 118 51 119 52 
rect 120 47 121 48 
rect 120 86 121 87 
rect 121 118 122 119 
rect 128 73 129 74 
rect 129 42 130 43 
rect 129 77 130 78 
rect 136 69 137 70 
rect 147 105 148 106 
rect 152 101 153 102 
<< end >>
3.99seconds.
