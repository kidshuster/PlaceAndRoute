magic
tech scmos
timestamp 58.9684
<< polysilicon >>
rect 10 10 11 11 
rect 10 11 11 12 
rect 10 12 11 13 
rect 10 13 11 14 
rect 10 14 11 15 
rect 10 15 11 16 
rect 10 26 11 27 
rect 10 27 11 28 
rect 10 28 11 29 
rect 10 29 11 30 
rect 10 30 11 31 
rect 10 31 11 32 
rect 10 42 11 43 
rect 10 43 11 44 
rect 10 44 11 45 
rect 10 45 11 46 
rect 10 46 11 47 
rect 10 47 11 48 
rect 10 58 11 59 
rect 10 59 11 60 
rect 10 60 11 61 
rect 10 61 11 62 
rect 10 63 11 64 
rect 10 74 11 75 
rect 10 76 11 77 
rect 10 77 11 78 
rect 10 79 11 80 
rect 10 90 11 91 
rect 10 91 11 92 
rect 10 92 11 93 
rect 10 93 11 94 
rect 10 94 11 95 
rect 10 95 11 96 
rect 10 106 11 107 
rect 10 107 11 108 
rect 10 108 11 109 
rect 10 109 11 110 
rect 10 110 11 111 
rect 10 111 11 112 
rect 10 138 11 139 
rect 10 140 11 141 
rect 10 141 11 142 
rect 10 143 11 144 
rect 10 154 11 155 
rect 10 155 11 156 
rect 10 156 11 157 
rect 10 157 11 158 
rect 10 158 11 159 
rect 10 159 11 160 
rect 10 170 11 171 
rect 10 172 11 173 
rect 10 173 11 174 
rect 10 174 11 175 
rect 10 175 11 176 
rect 10 186 11 187 
rect 10 188 11 189 
rect 10 189 11 190 
rect 10 191 11 192 
rect 10 202 11 203 
rect 10 204 11 205 
rect 10 205 11 206 
rect 10 207 11 208 
rect 10 218 11 219 
rect 10 220 11 221 
rect 10 221 11 222 
rect 10 222 11 223 
rect 10 223 11 224 
rect 10 234 11 235 
rect 10 236 11 237 
rect 10 237 11 238 
rect 10 238 11 239 
rect 10 239 11 240 
rect 10 250 11 251 
rect 10 252 11 253 
rect 10 253 11 254 
rect 10 254 11 255 
rect 10 255 11 256 
rect 10 266 11 267 
rect 10 267 11 268 
rect 10 268 11 269 
rect 10 269 11 270 
rect 10 270 11 271 
rect 10 271 11 272 
rect 10 282 11 283 
rect 10 283 11 284 
rect 10 284 11 285 
rect 10 285 11 286 
rect 10 286 11 287 
rect 10 287 11 288 
rect 10 298 11 299 
rect 10 300 11 301 
rect 10 301 11 302 
rect 10 302 11 303 
rect 10 303 11 304 
rect 11 10 12 11 
rect 11 11 12 12 
rect 11 12 12 13 
rect 11 13 12 14 
rect 11 14 12 15 
rect 11 15 12 16 
rect 11 26 12 27 
rect 11 27 12 28 
rect 11 28 12 29 
rect 11 29 12 30 
rect 11 30 12 31 
rect 11 31 12 32 
rect 11 42 12 43 
rect 11 43 12 44 
rect 11 44 12 45 
rect 11 45 12 46 
rect 11 46 12 47 
rect 11 47 12 48 
rect 11 58 12 59 
rect 11 59 12 60 
rect 11 60 12 61 
rect 11 61 12 62 
rect 11 62 12 63 
rect 11 63 12 64 
rect 11 74 12 75 
rect 11 75 12 76 
rect 11 76 12 77 
rect 11 77 12 78 
rect 11 78 12 79 
rect 11 79 12 80 
rect 11 90 12 91 
rect 11 91 12 92 
rect 11 92 12 93 
rect 11 93 12 94 
rect 11 94 12 95 
rect 11 95 12 96 
rect 11 106 12 107 
rect 11 107 12 108 
rect 11 108 12 109 
rect 11 109 12 110 
rect 11 110 12 111 
rect 11 111 12 112 
rect 11 138 12 139 
rect 11 139 12 140 
rect 11 140 12 141 
rect 11 141 12 142 
rect 11 142 12 143 
rect 11 143 12 144 
rect 11 154 12 155 
rect 11 155 12 156 
rect 11 156 12 157 
rect 11 157 12 158 
rect 11 158 12 159 
rect 11 159 12 160 
rect 11 170 12 171 
rect 11 171 12 172 
rect 11 172 12 173 
rect 11 173 12 174 
rect 11 174 12 175 
rect 11 175 12 176 
rect 11 186 12 187 
rect 11 187 12 188 
rect 11 188 12 189 
rect 11 189 12 190 
rect 11 190 12 191 
rect 11 191 12 192 
rect 11 202 12 203 
rect 11 203 12 204 
rect 11 204 12 205 
rect 11 205 12 206 
rect 11 206 12 207 
rect 11 207 12 208 
rect 11 218 12 219 
rect 11 219 12 220 
rect 11 220 12 221 
rect 11 221 12 222 
rect 11 222 12 223 
rect 11 223 12 224 
rect 11 234 12 235 
rect 11 235 12 236 
rect 11 236 12 237 
rect 11 237 12 238 
rect 11 238 12 239 
rect 11 239 12 240 
rect 11 250 12 251 
rect 11 251 12 252 
rect 11 252 12 253 
rect 11 253 12 254 
rect 11 254 12 255 
rect 11 255 12 256 
rect 11 266 12 267 
rect 11 267 12 268 
rect 11 268 12 269 
rect 11 269 12 270 
rect 11 270 12 271 
rect 11 271 12 272 
rect 11 282 12 283 
rect 11 283 12 284 
rect 11 284 12 285 
rect 11 285 12 286 
rect 11 286 12 287 
rect 11 287 12 288 
rect 11 298 12 299 
rect 11 299 12 300 
rect 11 300 12 301 
rect 11 301 12 302 
rect 11 302 12 303 
rect 11 303 12 304 
rect 12 10 13 11 
rect 12 11 13 12 
rect 12 12 13 13 
rect 12 13 13 14 
rect 12 14 13 15 
rect 12 15 13 16 
rect 12 26 13 27 
rect 12 27 13 28 
rect 12 28 13 29 
rect 12 29 13 30 
rect 12 30 13 31 
rect 12 31 13 32 
rect 12 42 13 43 
rect 12 43 13 44 
rect 12 44 13 45 
rect 12 45 13 46 
rect 12 46 13 47 
rect 12 47 13 48 
rect 12 58 13 59 
rect 12 59 13 60 
rect 12 60 13 61 
rect 12 61 13 62 
rect 12 62 13 63 
rect 12 63 13 64 
rect 12 74 13 75 
rect 12 75 13 76 
rect 12 76 13 77 
rect 12 77 13 78 
rect 12 78 13 79 
rect 12 79 13 80 
rect 12 90 13 91 
rect 12 91 13 92 
rect 12 92 13 93 
rect 12 93 13 94 
rect 12 94 13 95 
rect 12 95 13 96 
rect 12 106 13 107 
rect 12 107 13 108 
rect 12 108 13 109 
rect 12 109 13 110 
rect 12 110 13 111 
rect 12 111 13 112 
rect 12 138 13 139 
rect 12 139 13 140 
rect 12 140 13 141 
rect 12 141 13 142 
rect 12 142 13 143 
rect 12 143 13 144 
rect 12 154 13 155 
rect 12 155 13 156 
rect 12 156 13 157 
rect 12 157 13 158 
rect 12 158 13 159 
rect 12 159 13 160 
rect 12 170 13 171 
rect 12 171 13 172 
rect 12 172 13 173 
rect 12 173 13 174 
rect 12 174 13 175 
rect 12 175 13 176 
rect 12 186 13 187 
rect 12 187 13 188 
rect 12 188 13 189 
rect 12 189 13 190 
rect 12 190 13 191 
rect 12 191 13 192 
rect 12 202 13 203 
rect 12 203 13 204 
rect 12 204 13 205 
rect 12 205 13 206 
rect 12 206 13 207 
rect 12 207 13 208 
rect 12 218 13 219 
rect 12 219 13 220 
rect 12 220 13 221 
rect 12 221 13 222 
rect 12 222 13 223 
rect 12 223 13 224 
rect 12 234 13 235 
rect 12 235 13 236 
rect 12 236 13 237 
rect 12 237 13 238 
rect 12 238 13 239 
rect 12 239 13 240 
rect 12 250 13 251 
rect 12 251 13 252 
rect 12 252 13 253 
rect 12 253 13 254 
rect 12 254 13 255 
rect 12 255 13 256 
rect 12 266 13 267 
rect 12 267 13 268 
rect 12 268 13 269 
rect 12 269 13 270 
rect 12 270 13 271 
rect 12 271 13 272 
rect 12 282 13 283 
rect 12 283 13 284 
rect 12 284 13 285 
rect 12 285 13 286 
rect 12 286 13 287 
rect 12 287 13 288 
rect 12 298 13 299 
rect 12 299 13 300 
rect 12 300 13 301 
rect 12 301 13 302 
rect 12 302 13 303 
rect 12 303 13 304 
rect 13 10 14 11 
rect 13 11 14 12 
rect 13 12 14 13 
rect 13 13 14 14 
rect 13 14 14 15 
rect 13 15 14 16 
rect 13 26 14 27 
rect 13 27 14 28 
rect 13 28 14 29 
rect 13 29 14 30 
rect 13 30 14 31 
rect 13 31 14 32 
rect 13 42 14 43 
rect 13 43 14 44 
rect 13 44 14 45 
rect 13 45 14 46 
rect 13 46 14 47 
rect 13 47 14 48 
rect 13 58 14 59 
rect 13 59 14 60 
rect 13 60 14 61 
rect 13 61 14 62 
rect 13 62 14 63 
rect 13 63 14 64 
rect 13 74 14 75 
rect 13 75 14 76 
rect 13 76 14 77 
rect 13 77 14 78 
rect 13 78 14 79 
rect 13 79 14 80 
rect 13 90 14 91 
rect 13 91 14 92 
rect 13 92 14 93 
rect 13 93 14 94 
rect 13 94 14 95 
rect 13 95 14 96 
rect 13 106 14 107 
rect 13 107 14 108 
rect 13 108 14 109 
rect 13 109 14 110 
rect 13 110 14 111 
rect 13 111 14 112 
rect 13 138 14 139 
rect 13 139 14 140 
rect 13 140 14 141 
rect 13 141 14 142 
rect 13 142 14 143 
rect 13 143 14 144 
rect 13 154 14 155 
rect 13 155 14 156 
rect 13 156 14 157 
rect 13 157 14 158 
rect 13 158 14 159 
rect 13 159 14 160 
rect 13 170 14 171 
rect 13 171 14 172 
rect 13 172 14 173 
rect 13 173 14 174 
rect 13 174 14 175 
rect 13 175 14 176 
rect 13 186 14 187 
rect 13 187 14 188 
rect 13 188 14 189 
rect 13 189 14 190 
rect 13 190 14 191 
rect 13 191 14 192 
rect 13 202 14 203 
rect 13 203 14 204 
rect 13 204 14 205 
rect 13 205 14 206 
rect 13 206 14 207 
rect 13 207 14 208 
rect 13 218 14 219 
rect 13 219 14 220 
rect 13 220 14 221 
rect 13 221 14 222 
rect 13 222 14 223 
rect 13 223 14 224 
rect 13 234 14 235 
rect 13 235 14 236 
rect 13 236 14 237 
rect 13 237 14 238 
rect 13 238 14 239 
rect 13 239 14 240 
rect 13 250 14 251 
rect 13 251 14 252 
rect 13 252 14 253 
rect 13 253 14 254 
rect 13 254 14 255 
rect 13 255 14 256 
rect 13 266 14 267 
rect 13 267 14 268 
rect 13 268 14 269 
rect 13 269 14 270 
rect 13 270 14 271 
rect 13 271 14 272 
rect 13 282 14 283 
rect 13 283 14 284 
rect 13 284 14 285 
rect 13 285 14 286 
rect 13 286 14 287 
rect 13 287 14 288 
rect 13 298 14 299 
rect 13 299 14 300 
rect 13 300 14 301 
rect 13 301 14 302 
rect 13 302 14 303 
rect 13 303 14 304 
rect 14 10 15 11 
rect 14 11 15 12 
rect 14 12 15 13 
rect 14 13 15 14 
rect 14 14 15 15 
rect 14 15 15 16 
rect 14 26 15 27 
rect 14 27 15 28 
rect 14 28 15 29 
rect 14 29 15 30 
rect 14 30 15 31 
rect 14 31 15 32 
rect 14 42 15 43 
rect 14 43 15 44 
rect 14 44 15 45 
rect 14 45 15 46 
rect 14 46 15 47 
rect 14 47 15 48 
rect 14 58 15 59 
rect 14 59 15 60 
rect 14 60 15 61 
rect 14 61 15 62 
rect 14 62 15 63 
rect 14 63 15 64 
rect 14 74 15 75 
rect 14 75 15 76 
rect 14 76 15 77 
rect 14 77 15 78 
rect 14 78 15 79 
rect 14 79 15 80 
rect 14 90 15 91 
rect 14 91 15 92 
rect 14 92 15 93 
rect 14 93 15 94 
rect 14 94 15 95 
rect 14 95 15 96 
rect 14 106 15 107 
rect 14 107 15 108 
rect 14 108 15 109 
rect 14 109 15 110 
rect 14 110 15 111 
rect 14 111 15 112 
rect 14 138 15 139 
rect 14 139 15 140 
rect 14 140 15 141 
rect 14 141 15 142 
rect 14 142 15 143 
rect 14 143 15 144 
rect 14 154 15 155 
rect 14 155 15 156 
rect 14 156 15 157 
rect 14 157 15 158 
rect 14 158 15 159 
rect 14 159 15 160 
rect 14 170 15 171 
rect 14 171 15 172 
rect 14 172 15 173 
rect 14 173 15 174 
rect 14 174 15 175 
rect 14 175 15 176 
rect 14 186 15 187 
rect 14 187 15 188 
rect 14 188 15 189 
rect 14 189 15 190 
rect 14 190 15 191 
rect 14 191 15 192 
rect 14 202 15 203 
rect 14 203 15 204 
rect 14 204 15 205 
rect 14 205 15 206 
rect 14 206 15 207 
rect 14 207 15 208 
rect 14 218 15 219 
rect 14 219 15 220 
rect 14 220 15 221 
rect 14 221 15 222 
rect 14 222 15 223 
rect 14 223 15 224 
rect 14 234 15 235 
rect 14 235 15 236 
rect 14 236 15 237 
rect 14 237 15 238 
rect 14 238 15 239 
rect 14 239 15 240 
rect 14 250 15 251 
rect 14 251 15 252 
rect 14 252 15 253 
rect 14 253 15 254 
rect 14 254 15 255 
rect 14 255 15 256 
rect 14 266 15 267 
rect 14 267 15 268 
rect 14 268 15 269 
rect 14 269 15 270 
rect 14 270 15 271 
rect 14 271 15 272 
rect 14 282 15 283 
rect 14 283 15 284 
rect 14 284 15 285 
rect 14 285 15 286 
rect 14 286 15 287 
rect 14 287 15 288 
rect 14 298 15 299 
rect 14 299 15 300 
rect 14 300 15 301 
rect 14 301 15 302 
rect 14 302 15 303 
rect 14 303 15 304 
rect 15 10 16 11 
rect 15 11 16 12 
rect 15 12 16 13 
rect 15 13 16 14 
rect 15 14 16 15 
rect 15 15 16 16 
rect 15 26 16 27 
rect 15 27 16 28 
rect 15 28 16 29 
rect 15 29 16 30 
rect 15 30 16 31 
rect 15 31 16 32 
rect 15 42 16 43 
rect 15 43 16 44 
rect 15 44 16 45 
rect 15 45 16 46 
rect 15 46 16 47 
rect 15 47 16 48 
rect 15 58 16 59 
rect 15 59 16 60 
rect 15 60 16 61 
rect 15 61 16 62 
rect 15 62 16 63 
rect 15 63 16 64 
rect 15 74 16 75 
rect 15 75 16 76 
rect 15 76 16 77 
rect 15 77 16 78 
rect 15 79 16 80 
rect 15 90 16 91 
rect 15 91 16 92 
rect 15 92 16 93 
rect 15 93 16 94 
rect 15 94 16 95 
rect 15 95 16 96 
rect 15 106 16 107 
rect 15 108 16 109 
rect 15 109 16 110 
rect 15 110 16 111 
rect 15 111 16 112 
rect 15 138 16 139 
rect 15 140 16 141 
rect 15 141 16 142 
rect 15 143 16 144 
rect 15 154 16 155 
rect 15 156 16 157 
rect 15 157 16 158 
rect 15 158 16 159 
rect 15 159 16 160 
rect 15 170 16 171 
rect 15 171 16 172 
rect 15 172 16 173 
rect 15 173 16 174 
rect 15 175 16 176 
rect 15 186 16 187 
rect 15 187 16 188 
rect 15 188 16 189 
rect 15 189 16 190 
rect 15 191 16 192 
rect 15 202 16 203 
rect 15 204 16 205 
rect 15 205 16 206 
rect 15 206 16 207 
rect 15 207 16 208 
rect 15 218 16 219 
rect 15 219 16 220 
rect 15 220 16 221 
rect 15 221 16 222 
rect 15 222 16 223 
rect 15 223 16 224 
rect 15 234 16 235 
rect 15 235 16 236 
rect 15 236 16 237 
rect 15 237 16 238 
rect 15 238 16 239 
rect 15 239 16 240 
rect 15 250 16 251 
rect 15 251 16 252 
rect 15 252 16 253 
rect 15 253 16 254 
rect 15 254 16 255 
rect 15 255 16 256 
rect 15 266 16 267 
rect 15 267 16 268 
rect 15 268 16 269 
rect 15 269 16 270 
rect 15 270 16 271 
rect 15 271 16 272 
rect 15 282 16 283 
rect 15 283 16 284 
rect 15 284 16 285 
rect 15 285 16 286 
rect 15 287 16 288 
rect 15 298 16 299 
rect 15 299 16 300 
rect 15 300 16 301 
rect 15 301 16 302 
rect 15 302 16 303 
rect 15 303 16 304 
rect 26 10 27 11 
rect 26 11 27 12 
rect 26 12 27 13 
rect 26 13 27 14 
rect 26 14 27 15 
rect 26 15 27 16 
rect 26 26 27 27 
rect 26 27 27 28 
rect 26 28 27 29 
rect 26 29 27 30 
rect 26 30 27 31 
rect 26 31 27 32 
rect 26 42 27 43 
rect 26 43 27 44 
rect 26 44 27 45 
rect 26 45 27 46 
rect 26 46 27 47 
rect 26 47 27 48 
rect 26 58 27 59 
rect 26 59 27 60 
rect 26 60 27 61 
rect 26 61 27 62 
rect 26 62 27 63 
rect 26 63 27 64 
rect 26 74 27 75 
rect 26 76 27 77 
rect 26 77 27 78 
rect 26 79 27 80 
rect 26 90 27 91 
rect 26 91 27 92 
rect 26 92 27 93 
rect 26 93 27 94 
rect 26 94 27 95 
rect 26 95 27 96 
rect 26 106 27 107 
rect 26 108 27 109 
rect 26 109 27 110 
rect 26 111 27 112 
rect 26 138 27 139 
rect 26 140 27 141 
rect 26 141 27 142 
rect 26 142 27 143 
rect 26 143 27 144 
rect 26 154 27 155 
rect 26 156 27 157 
rect 26 157 27 158 
rect 26 158 27 159 
rect 26 159 27 160 
rect 26 170 27 171 
rect 26 171 27 172 
rect 26 172 27 173 
rect 26 173 27 174 
rect 26 175 27 176 
rect 26 186 27 187 
rect 26 187 27 188 
rect 26 188 27 189 
rect 26 189 27 190 
rect 26 190 27 191 
rect 26 191 27 192 
rect 26 202 27 203 
rect 26 204 27 205 
rect 26 205 27 206 
rect 26 207 27 208 
rect 26 218 27 219 
rect 26 220 27 221 
rect 26 221 27 222 
rect 26 222 27 223 
rect 26 223 27 224 
rect 26 234 27 235 
rect 26 235 27 236 
rect 26 236 27 237 
rect 26 237 27 238 
rect 26 238 27 239 
rect 26 239 27 240 
rect 26 250 27 251 
rect 26 252 27 253 
rect 26 253 27 254 
rect 26 254 27 255 
rect 26 255 27 256 
rect 26 266 27 267 
rect 26 267 27 268 
rect 26 268 27 269 
rect 26 269 27 270 
rect 26 270 27 271 
rect 26 271 27 272 
rect 26 282 27 283 
rect 26 283 27 284 
rect 26 284 27 285 
rect 26 285 27 286 
rect 26 287 27 288 
rect 26 298 27 299 
rect 26 300 27 301 
rect 26 301 27 302 
rect 26 302 27 303 
rect 26 303 27 304 
rect 27 10 28 11 
rect 27 11 28 12 
rect 27 12 28 13 
rect 27 13 28 14 
rect 27 14 28 15 
rect 27 15 28 16 
rect 27 26 28 27 
rect 27 27 28 28 
rect 27 28 28 29 
rect 27 29 28 30 
rect 27 30 28 31 
rect 27 31 28 32 
rect 27 42 28 43 
rect 27 43 28 44 
rect 27 44 28 45 
rect 27 45 28 46 
rect 27 46 28 47 
rect 27 47 28 48 
rect 27 58 28 59 
rect 27 59 28 60 
rect 27 60 28 61 
rect 27 61 28 62 
rect 27 62 28 63 
rect 27 63 28 64 
rect 27 74 28 75 
rect 27 75 28 76 
rect 27 76 28 77 
rect 27 77 28 78 
rect 27 78 28 79 
rect 27 79 28 80 
rect 27 90 28 91 
rect 27 91 28 92 
rect 27 92 28 93 
rect 27 93 28 94 
rect 27 94 28 95 
rect 27 95 28 96 
rect 27 106 28 107 
rect 27 107 28 108 
rect 27 108 28 109 
rect 27 109 28 110 
rect 27 110 28 111 
rect 27 111 28 112 
rect 27 138 28 139 
rect 27 139 28 140 
rect 27 140 28 141 
rect 27 141 28 142 
rect 27 142 28 143 
rect 27 143 28 144 
rect 27 154 28 155 
rect 27 155 28 156 
rect 27 156 28 157 
rect 27 157 28 158 
rect 27 158 28 159 
rect 27 159 28 160 
rect 27 170 28 171 
rect 27 171 28 172 
rect 27 172 28 173 
rect 27 173 28 174 
rect 27 174 28 175 
rect 27 175 28 176 
rect 27 186 28 187 
rect 27 187 28 188 
rect 27 188 28 189 
rect 27 189 28 190 
rect 27 190 28 191 
rect 27 191 28 192 
rect 27 202 28 203 
rect 27 203 28 204 
rect 27 204 28 205 
rect 27 205 28 206 
rect 27 206 28 207 
rect 27 207 28 208 
rect 27 218 28 219 
rect 27 219 28 220 
rect 27 220 28 221 
rect 27 221 28 222 
rect 27 222 28 223 
rect 27 223 28 224 
rect 27 234 28 235 
rect 27 235 28 236 
rect 27 236 28 237 
rect 27 237 28 238 
rect 27 238 28 239 
rect 27 239 28 240 
rect 27 250 28 251 
rect 27 251 28 252 
rect 27 252 28 253 
rect 27 253 28 254 
rect 27 254 28 255 
rect 27 255 28 256 
rect 27 266 28 267 
rect 27 267 28 268 
rect 27 268 28 269 
rect 27 269 28 270 
rect 27 270 28 271 
rect 27 271 28 272 
rect 27 282 28 283 
rect 27 283 28 284 
rect 27 284 28 285 
rect 27 285 28 286 
rect 27 286 28 287 
rect 27 287 28 288 
rect 27 298 28 299 
rect 27 299 28 300 
rect 27 300 28 301 
rect 27 301 28 302 
rect 27 302 28 303 
rect 27 303 28 304 
rect 28 10 29 11 
rect 28 11 29 12 
rect 28 12 29 13 
rect 28 13 29 14 
rect 28 14 29 15 
rect 28 15 29 16 
rect 28 26 29 27 
rect 28 27 29 28 
rect 28 28 29 29 
rect 28 29 29 30 
rect 28 30 29 31 
rect 28 31 29 32 
rect 28 42 29 43 
rect 28 43 29 44 
rect 28 44 29 45 
rect 28 45 29 46 
rect 28 46 29 47 
rect 28 47 29 48 
rect 28 58 29 59 
rect 28 59 29 60 
rect 28 60 29 61 
rect 28 61 29 62 
rect 28 62 29 63 
rect 28 63 29 64 
rect 28 74 29 75 
rect 28 75 29 76 
rect 28 76 29 77 
rect 28 77 29 78 
rect 28 78 29 79 
rect 28 79 29 80 
rect 28 90 29 91 
rect 28 91 29 92 
rect 28 92 29 93 
rect 28 93 29 94 
rect 28 94 29 95 
rect 28 95 29 96 
rect 28 106 29 107 
rect 28 107 29 108 
rect 28 108 29 109 
rect 28 109 29 110 
rect 28 110 29 111 
rect 28 111 29 112 
rect 28 138 29 139 
rect 28 139 29 140 
rect 28 140 29 141 
rect 28 141 29 142 
rect 28 142 29 143 
rect 28 143 29 144 
rect 28 154 29 155 
rect 28 155 29 156 
rect 28 156 29 157 
rect 28 157 29 158 
rect 28 158 29 159 
rect 28 159 29 160 
rect 28 170 29 171 
rect 28 171 29 172 
rect 28 172 29 173 
rect 28 173 29 174 
rect 28 174 29 175 
rect 28 175 29 176 
rect 28 186 29 187 
rect 28 187 29 188 
rect 28 188 29 189 
rect 28 189 29 190 
rect 28 190 29 191 
rect 28 191 29 192 
rect 28 202 29 203 
rect 28 203 29 204 
rect 28 204 29 205 
rect 28 205 29 206 
rect 28 206 29 207 
rect 28 207 29 208 
rect 28 218 29 219 
rect 28 219 29 220 
rect 28 220 29 221 
rect 28 221 29 222 
rect 28 222 29 223 
rect 28 223 29 224 
rect 28 234 29 235 
rect 28 235 29 236 
rect 28 236 29 237 
rect 28 237 29 238 
rect 28 238 29 239 
rect 28 239 29 240 
rect 28 250 29 251 
rect 28 251 29 252 
rect 28 252 29 253 
rect 28 253 29 254 
rect 28 254 29 255 
rect 28 255 29 256 
rect 28 266 29 267 
rect 28 267 29 268 
rect 28 268 29 269 
rect 28 269 29 270 
rect 28 270 29 271 
rect 28 271 29 272 
rect 28 282 29 283 
rect 28 283 29 284 
rect 28 284 29 285 
rect 28 285 29 286 
rect 28 286 29 287 
rect 28 287 29 288 
rect 28 298 29 299 
rect 28 299 29 300 
rect 28 300 29 301 
rect 28 301 29 302 
rect 28 302 29 303 
rect 28 303 29 304 
rect 29 10 30 11 
rect 29 11 30 12 
rect 29 12 30 13 
rect 29 13 30 14 
rect 29 14 30 15 
rect 29 15 30 16 
rect 29 26 30 27 
rect 29 27 30 28 
rect 29 28 30 29 
rect 29 29 30 30 
rect 29 30 30 31 
rect 29 31 30 32 
rect 29 42 30 43 
rect 29 43 30 44 
rect 29 44 30 45 
rect 29 45 30 46 
rect 29 46 30 47 
rect 29 47 30 48 
rect 29 58 30 59 
rect 29 59 30 60 
rect 29 60 30 61 
rect 29 61 30 62 
rect 29 62 30 63 
rect 29 63 30 64 
rect 29 74 30 75 
rect 29 75 30 76 
rect 29 76 30 77 
rect 29 77 30 78 
rect 29 78 30 79 
rect 29 79 30 80 
rect 29 90 30 91 
rect 29 91 30 92 
rect 29 92 30 93 
rect 29 93 30 94 
rect 29 94 30 95 
rect 29 95 30 96 
rect 29 106 30 107 
rect 29 107 30 108 
rect 29 108 30 109 
rect 29 109 30 110 
rect 29 110 30 111 
rect 29 111 30 112 
rect 29 138 30 139 
rect 29 139 30 140 
rect 29 140 30 141 
rect 29 141 30 142 
rect 29 142 30 143 
rect 29 143 30 144 
rect 29 154 30 155 
rect 29 155 30 156 
rect 29 156 30 157 
rect 29 157 30 158 
rect 29 158 30 159 
rect 29 159 30 160 
rect 29 170 30 171 
rect 29 171 30 172 
rect 29 172 30 173 
rect 29 173 30 174 
rect 29 174 30 175 
rect 29 175 30 176 
rect 29 186 30 187 
rect 29 187 30 188 
rect 29 188 30 189 
rect 29 189 30 190 
rect 29 190 30 191 
rect 29 191 30 192 
rect 29 202 30 203 
rect 29 203 30 204 
rect 29 204 30 205 
rect 29 205 30 206 
rect 29 206 30 207 
rect 29 207 30 208 
rect 29 218 30 219 
rect 29 219 30 220 
rect 29 220 30 221 
rect 29 221 30 222 
rect 29 222 30 223 
rect 29 223 30 224 
rect 29 234 30 235 
rect 29 235 30 236 
rect 29 236 30 237 
rect 29 237 30 238 
rect 29 238 30 239 
rect 29 239 30 240 
rect 29 250 30 251 
rect 29 251 30 252 
rect 29 252 30 253 
rect 29 253 30 254 
rect 29 254 30 255 
rect 29 255 30 256 
rect 29 266 30 267 
rect 29 267 30 268 
rect 29 268 30 269 
rect 29 269 30 270 
rect 29 270 30 271 
rect 29 271 30 272 
rect 29 282 30 283 
rect 29 283 30 284 
rect 29 284 30 285 
rect 29 285 30 286 
rect 29 286 30 287 
rect 29 287 30 288 
rect 29 298 30 299 
rect 29 299 30 300 
rect 29 300 30 301 
rect 29 301 30 302 
rect 29 302 30 303 
rect 29 303 30 304 
rect 30 10 31 11 
rect 30 11 31 12 
rect 30 12 31 13 
rect 30 13 31 14 
rect 30 14 31 15 
rect 30 15 31 16 
rect 30 26 31 27 
rect 30 27 31 28 
rect 30 28 31 29 
rect 30 29 31 30 
rect 30 30 31 31 
rect 30 31 31 32 
rect 30 42 31 43 
rect 30 43 31 44 
rect 30 44 31 45 
rect 30 45 31 46 
rect 30 46 31 47 
rect 30 47 31 48 
rect 30 58 31 59 
rect 30 59 31 60 
rect 30 60 31 61 
rect 30 61 31 62 
rect 30 62 31 63 
rect 30 63 31 64 
rect 30 74 31 75 
rect 30 75 31 76 
rect 30 76 31 77 
rect 30 77 31 78 
rect 30 78 31 79 
rect 30 79 31 80 
rect 30 90 31 91 
rect 30 91 31 92 
rect 30 92 31 93 
rect 30 93 31 94 
rect 30 94 31 95 
rect 30 95 31 96 
rect 30 106 31 107 
rect 30 107 31 108 
rect 30 108 31 109 
rect 30 109 31 110 
rect 30 110 31 111 
rect 30 111 31 112 
rect 30 138 31 139 
rect 30 139 31 140 
rect 30 140 31 141 
rect 30 141 31 142 
rect 30 142 31 143 
rect 30 143 31 144 
rect 30 154 31 155 
rect 30 155 31 156 
rect 30 156 31 157 
rect 30 157 31 158 
rect 30 158 31 159 
rect 30 159 31 160 
rect 30 170 31 171 
rect 30 171 31 172 
rect 30 172 31 173 
rect 30 173 31 174 
rect 30 174 31 175 
rect 30 175 31 176 
rect 30 186 31 187 
rect 30 187 31 188 
rect 30 188 31 189 
rect 30 189 31 190 
rect 30 190 31 191 
rect 30 191 31 192 
rect 30 202 31 203 
rect 30 203 31 204 
rect 30 204 31 205 
rect 30 205 31 206 
rect 30 206 31 207 
rect 30 207 31 208 
rect 30 218 31 219 
rect 30 219 31 220 
rect 30 220 31 221 
rect 30 221 31 222 
rect 30 222 31 223 
rect 30 223 31 224 
rect 30 234 31 235 
rect 30 235 31 236 
rect 30 236 31 237 
rect 30 237 31 238 
rect 30 238 31 239 
rect 30 239 31 240 
rect 30 250 31 251 
rect 30 251 31 252 
rect 30 252 31 253 
rect 30 253 31 254 
rect 30 254 31 255 
rect 30 255 31 256 
rect 30 266 31 267 
rect 30 267 31 268 
rect 30 268 31 269 
rect 30 269 31 270 
rect 30 270 31 271 
rect 30 271 31 272 
rect 30 282 31 283 
rect 30 283 31 284 
rect 30 284 31 285 
rect 30 285 31 286 
rect 30 286 31 287 
rect 30 287 31 288 
rect 30 298 31 299 
rect 30 299 31 300 
rect 30 300 31 301 
rect 30 301 31 302 
rect 30 302 31 303 
rect 30 303 31 304 
rect 31 10 32 11 
rect 31 11 32 12 
rect 31 12 32 13 
rect 31 13 32 14 
rect 31 15 32 16 
rect 31 26 32 27 
rect 31 27 32 28 
rect 31 28 32 29 
rect 31 29 32 30 
rect 31 30 32 31 
rect 31 31 32 32 
rect 31 42 32 43 
rect 31 43 32 44 
rect 31 44 32 45 
rect 31 45 32 46 
rect 31 46 32 47 
rect 31 47 32 48 
rect 31 58 32 59 
rect 31 60 32 61 
rect 31 61 32 62 
rect 31 63 32 64 
rect 31 74 32 75 
rect 31 75 32 76 
rect 31 76 32 77 
rect 31 77 32 78 
rect 31 78 32 79 
rect 31 79 32 80 
rect 31 90 32 91 
rect 31 91 32 92 
rect 31 92 32 93 
rect 31 93 32 94 
rect 31 94 32 95 
rect 31 95 32 96 
rect 31 106 32 107 
rect 31 108 32 109 
rect 31 109 32 110 
rect 31 110 32 111 
rect 31 111 32 112 
rect 31 138 32 139 
rect 31 140 32 141 
rect 31 141 32 142 
rect 31 142 32 143 
rect 31 143 32 144 
rect 31 154 32 155 
rect 31 156 32 157 
rect 31 157 32 158 
rect 31 158 32 159 
rect 31 159 32 160 
rect 31 170 32 171 
rect 31 171 32 172 
rect 31 172 32 173 
rect 31 173 32 174 
rect 31 174 32 175 
rect 31 175 32 176 
rect 31 186 32 187 
rect 31 187 32 188 
rect 31 188 32 189 
rect 31 189 32 190 
rect 31 190 32 191 
rect 31 191 32 192 
rect 31 202 32 203 
rect 31 203 32 204 
rect 31 204 32 205 
rect 31 205 32 206 
rect 31 206 32 207 
rect 31 207 32 208 
rect 31 218 32 219 
rect 31 220 32 221 
rect 31 221 32 222 
rect 31 223 32 224 
rect 31 234 32 235 
rect 31 236 32 237 
rect 31 237 32 238 
rect 31 238 32 239 
rect 31 239 32 240 
rect 31 250 32 251 
rect 31 252 32 253 
rect 31 253 32 254 
rect 31 255 32 256 
rect 31 266 32 267 
rect 31 267 32 268 
rect 31 268 32 269 
rect 31 269 32 270 
rect 31 271 32 272 
rect 31 282 32 283 
rect 31 284 32 285 
rect 31 285 32 286 
rect 31 286 32 287 
rect 31 287 32 288 
rect 31 298 32 299 
rect 31 300 32 301 
rect 31 301 32 302 
rect 31 302 32 303 
rect 31 303 32 304 
rect 42 10 43 11 
rect 42 11 43 12 
rect 42 12 43 13 
rect 42 13 43 14 
rect 42 14 43 15 
rect 42 15 43 16 
rect 42 26 43 27 
rect 42 27 43 28 
rect 42 28 43 29 
rect 42 29 43 30 
rect 42 31 43 32 
rect 42 42 43 43 
rect 42 44 43 45 
rect 42 45 43 46 
rect 42 47 43 48 
rect 42 58 43 59 
rect 42 60 43 61 
rect 42 61 43 62 
rect 42 62 43 63 
rect 42 63 43 64 
rect 42 74 43 75 
rect 42 75 43 76 
rect 42 76 43 77 
rect 42 77 43 78 
rect 42 79 43 80 
rect 42 90 43 91 
rect 42 92 43 93 
rect 42 93 43 94 
rect 42 94 43 95 
rect 42 95 43 96 
rect 42 106 43 107 
rect 42 107 43 108 
rect 42 108 43 109 
rect 42 109 43 110 
rect 42 111 43 112 
rect 42 122 43 123 
rect 42 124 43 125 
rect 42 125 43 126 
rect 42 127 43 128 
rect 42 138 43 139 
rect 42 139 43 140 
rect 42 140 43 141 
rect 42 141 43 142 
rect 42 143 43 144 
rect 42 154 43 155 
rect 42 155 43 156 
rect 42 156 43 157 
rect 42 157 43 158 
rect 42 158 43 159 
rect 42 159 43 160 
rect 42 170 43 171 
rect 42 172 43 173 
rect 42 173 43 174 
rect 42 175 43 176 
rect 42 186 43 187 
rect 42 188 43 189 
rect 42 189 43 190 
rect 42 190 43 191 
rect 42 191 43 192 
rect 42 202 43 203 
rect 42 203 43 204 
rect 42 204 43 205 
rect 42 205 43 206 
rect 42 207 43 208 
rect 42 218 43 219 
rect 42 220 43 221 
rect 42 221 43 222 
rect 42 223 43 224 
rect 42 234 43 235 
rect 42 235 43 236 
rect 42 236 43 237 
rect 42 237 43 238 
rect 42 238 43 239 
rect 42 239 43 240 
rect 42 250 43 251 
rect 42 252 43 253 
rect 42 253 43 254 
rect 42 255 43 256 
rect 42 266 43 267 
rect 42 268 43 269 
rect 42 269 43 270 
rect 42 270 43 271 
rect 42 271 43 272 
rect 42 282 43 283 
rect 42 283 43 284 
rect 42 284 43 285 
rect 42 285 43 286 
rect 42 286 43 287 
rect 42 287 43 288 
rect 42 298 43 299 
rect 42 299 43 300 
rect 42 300 43 301 
rect 42 301 43 302 
rect 42 303 43 304 
rect 43 10 44 11 
rect 43 11 44 12 
rect 43 12 44 13 
rect 43 13 44 14 
rect 43 14 44 15 
rect 43 15 44 16 
rect 43 26 44 27 
rect 43 27 44 28 
rect 43 28 44 29 
rect 43 29 44 30 
rect 43 30 44 31 
rect 43 31 44 32 
rect 43 42 44 43 
rect 43 43 44 44 
rect 43 44 44 45 
rect 43 45 44 46 
rect 43 46 44 47 
rect 43 47 44 48 
rect 43 58 44 59 
rect 43 59 44 60 
rect 43 60 44 61 
rect 43 61 44 62 
rect 43 62 44 63 
rect 43 63 44 64 
rect 43 74 44 75 
rect 43 75 44 76 
rect 43 76 44 77 
rect 43 77 44 78 
rect 43 78 44 79 
rect 43 79 44 80 
rect 43 90 44 91 
rect 43 91 44 92 
rect 43 92 44 93 
rect 43 93 44 94 
rect 43 94 44 95 
rect 43 95 44 96 
rect 43 106 44 107 
rect 43 107 44 108 
rect 43 108 44 109 
rect 43 109 44 110 
rect 43 110 44 111 
rect 43 111 44 112 
rect 43 122 44 123 
rect 43 123 44 124 
rect 43 124 44 125 
rect 43 125 44 126 
rect 43 126 44 127 
rect 43 127 44 128 
rect 43 138 44 139 
rect 43 139 44 140 
rect 43 140 44 141 
rect 43 141 44 142 
rect 43 142 44 143 
rect 43 143 44 144 
rect 43 154 44 155 
rect 43 155 44 156 
rect 43 156 44 157 
rect 43 157 44 158 
rect 43 158 44 159 
rect 43 159 44 160 
rect 43 170 44 171 
rect 43 171 44 172 
rect 43 172 44 173 
rect 43 173 44 174 
rect 43 174 44 175 
rect 43 175 44 176 
rect 43 186 44 187 
rect 43 187 44 188 
rect 43 188 44 189 
rect 43 189 44 190 
rect 43 190 44 191 
rect 43 191 44 192 
rect 43 202 44 203 
rect 43 203 44 204 
rect 43 204 44 205 
rect 43 205 44 206 
rect 43 206 44 207 
rect 43 207 44 208 
rect 43 218 44 219 
rect 43 219 44 220 
rect 43 220 44 221 
rect 43 221 44 222 
rect 43 222 44 223 
rect 43 223 44 224 
rect 43 234 44 235 
rect 43 235 44 236 
rect 43 236 44 237 
rect 43 237 44 238 
rect 43 238 44 239 
rect 43 239 44 240 
rect 43 250 44 251 
rect 43 251 44 252 
rect 43 252 44 253 
rect 43 253 44 254 
rect 43 254 44 255 
rect 43 255 44 256 
rect 43 266 44 267 
rect 43 267 44 268 
rect 43 268 44 269 
rect 43 269 44 270 
rect 43 270 44 271 
rect 43 271 44 272 
rect 43 282 44 283 
rect 43 283 44 284 
rect 43 284 44 285 
rect 43 285 44 286 
rect 43 286 44 287 
rect 43 287 44 288 
rect 43 298 44 299 
rect 43 299 44 300 
rect 43 300 44 301 
rect 43 301 44 302 
rect 43 302 44 303 
rect 43 303 44 304 
rect 44 10 45 11 
rect 44 11 45 12 
rect 44 12 45 13 
rect 44 13 45 14 
rect 44 14 45 15 
rect 44 15 45 16 
rect 44 26 45 27 
rect 44 27 45 28 
rect 44 28 45 29 
rect 44 29 45 30 
rect 44 30 45 31 
rect 44 31 45 32 
rect 44 42 45 43 
rect 44 43 45 44 
rect 44 44 45 45 
rect 44 45 45 46 
rect 44 46 45 47 
rect 44 47 45 48 
rect 44 58 45 59 
rect 44 59 45 60 
rect 44 60 45 61 
rect 44 61 45 62 
rect 44 62 45 63 
rect 44 63 45 64 
rect 44 74 45 75 
rect 44 75 45 76 
rect 44 76 45 77 
rect 44 77 45 78 
rect 44 78 45 79 
rect 44 79 45 80 
rect 44 90 45 91 
rect 44 91 45 92 
rect 44 92 45 93 
rect 44 93 45 94 
rect 44 94 45 95 
rect 44 95 45 96 
rect 44 106 45 107 
rect 44 107 45 108 
rect 44 108 45 109 
rect 44 109 45 110 
rect 44 110 45 111 
rect 44 111 45 112 
rect 44 122 45 123 
rect 44 123 45 124 
rect 44 124 45 125 
rect 44 125 45 126 
rect 44 126 45 127 
rect 44 127 45 128 
rect 44 138 45 139 
rect 44 139 45 140 
rect 44 140 45 141 
rect 44 141 45 142 
rect 44 142 45 143 
rect 44 143 45 144 
rect 44 154 45 155 
rect 44 155 45 156 
rect 44 156 45 157 
rect 44 157 45 158 
rect 44 158 45 159 
rect 44 159 45 160 
rect 44 170 45 171 
rect 44 171 45 172 
rect 44 172 45 173 
rect 44 173 45 174 
rect 44 174 45 175 
rect 44 175 45 176 
rect 44 186 45 187 
rect 44 187 45 188 
rect 44 188 45 189 
rect 44 189 45 190 
rect 44 190 45 191 
rect 44 191 45 192 
rect 44 202 45 203 
rect 44 203 45 204 
rect 44 204 45 205 
rect 44 205 45 206 
rect 44 206 45 207 
rect 44 207 45 208 
rect 44 218 45 219 
rect 44 219 45 220 
rect 44 220 45 221 
rect 44 221 45 222 
rect 44 222 45 223 
rect 44 223 45 224 
rect 44 234 45 235 
rect 44 235 45 236 
rect 44 236 45 237 
rect 44 237 45 238 
rect 44 238 45 239 
rect 44 239 45 240 
rect 44 250 45 251 
rect 44 251 45 252 
rect 44 252 45 253 
rect 44 253 45 254 
rect 44 254 45 255 
rect 44 255 45 256 
rect 44 266 45 267 
rect 44 267 45 268 
rect 44 268 45 269 
rect 44 269 45 270 
rect 44 270 45 271 
rect 44 271 45 272 
rect 44 282 45 283 
rect 44 283 45 284 
rect 44 284 45 285 
rect 44 285 45 286 
rect 44 286 45 287 
rect 44 287 45 288 
rect 44 298 45 299 
rect 44 299 45 300 
rect 44 300 45 301 
rect 44 301 45 302 
rect 44 302 45 303 
rect 44 303 45 304 
rect 45 10 46 11 
rect 45 11 46 12 
rect 45 12 46 13 
rect 45 13 46 14 
rect 45 14 46 15 
rect 45 15 46 16 
rect 45 26 46 27 
rect 45 27 46 28 
rect 45 28 46 29 
rect 45 29 46 30 
rect 45 30 46 31 
rect 45 31 46 32 
rect 45 42 46 43 
rect 45 43 46 44 
rect 45 44 46 45 
rect 45 45 46 46 
rect 45 46 46 47 
rect 45 47 46 48 
rect 45 58 46 59 
rect 45 59 46 60 
rect 45 60 46 61 
rect 45 61 46 62 
rect 45 62 46 63 
rect 45 63 46 64 
rect 45 74 46 75 
rect 45 75 46 76 
rect 45 76 46 77 
rect 45 77 46 78 
rect 45 78 46 79 
rect 45 79 46 80 
rect 45 90 46 91 
rect 45 91 46 92 
rect 45 92 46 93 
rect 45 93 46 94 
rect 45 94 46 95 
rect 45 95 46 96 
rect 45 106 46 107 
rect 45 107 46 108 
rect 45 108 46 109 
rect 45 109 46 110 
rect 45 110 46 111 
rect 45 111 46 112 
rect 45 122 46 123 
rect 45 123 46 124 
rect 45 124 46 125 
rect 45 125 46 126 
rect 45 126 46 127 
rect 45 127 46 128 
rect 45 138 46 139 
rect 45 139 46 140 
rect 45 140 46 141 
rect 45 141 46 142 
rect 45 142 46 143 
rect 45 143 46 144 
rect 45 154 46 155 
rect 45 155 46 156 
rect 45 156 46 157 
rect 45 157 46 158 
rect 45 158 46 159 
rect 45 159 46 160 
rect 45 170 46 171 
rect 45 171 46 172 
rect 45 172 46 173 
rect 45 173 46 174 
rect 45 174 46 175 
rect 45 175 46 176 
rect 45 186 46 187 
rect 45 187 46 188 
rect 45 188 46 189 
rect 45 189 46 190 
rect 45 190 46 191 
rect 45 191 46 192 
rect 45 202 46 203 
rect 45 203 46 204 
rect 45 204 46 205 
rect 45 205 46 206 
rect 45 206 46 207 
rect 45 207 46 208 
rect 45 218 46 219 
rect 45 219 46 220 
rect 45 220 46 221 
rect 45 221 46 222 
rect 45 222 46 223 
rect 45 223 46 224 
rect 45 234 46 235 
rect 45 235 46 236 
rect 45 236 46 237 
rect 45 237 46 238 
rect 45 238 46 239 
rect 45 239 46 240 
rect 45 250 46 251 
rect 45 251 46 252 
rect 45 252 46 253 
rect 45 253 46 254 
rect 45 254 46 255 
rect 45 255 46 256 
rect 45 266 46 267 
rect 45 267 46 268 
rect 45 268 46 269 
rect 45 269 46 270 
rect 45 270 46 271 
rect 45 271 46 272 
rect 45 282 46 283 
rect 45 283 46 284 
rect 45 284 46 285 
rect 45 285 46 286 
rect 45 286 46 287 
rect 45 287 46 288 
rect 45 298 46 299 
rect 45 299 46 300 
rect 45 300 46 301 
rect 45 301 46 302 
rect 45 302 46 303 
rect 45 303 46 304 
rect 46 10 47 11 
rect 46 11 47 12 
rect 46 12 47 13 
rect 46 13 47 14 
rect 46 14 47 15 
rect 46 15 47 16 
rect 46 26 47 27 
rect 46 27 47 28 
rect 46 28 47 29 
rect 46 29 47 30 
rect 46 30 47 31 
rect 46 31 47 32 
rect 46 42 47 43 
rect 46 43 47 44 
rect 46 44 47 45 
rect 46 45 47 46 
rect 46 46 47 47 
rect 46 47 47 48 
rect 46 58 47 59 
rect 46 59 47 60 
rect 46 60 47 61 
rect 46 61 47 62 
rect 46 62 47 63 
rect 46 63 47 64 
rect 46 74 47 75 
rect 46 75 47 76 
rect 46 76 47 77 
rect 46 77 47 78 
rect 46 78 47 79 
rect 46 79 47 80 
rect 46 90 47 91 
rect 46 91 47 92 
rect 46 92 47 93 
rect 46 93 47 94 
rect 46 94 47 95 
rect 46 95 47 96 
rect 46 106 47 107 
rect 46 107 47 108 
rect 46 108 47 109 
rect 46 109 47 110 
rect 46 110 47 111 
rect 46 111 47 112 
rect 46 122 47 123 
rect 46 123 47 124 
rect 46 124 47 125 
rect 46 125 47 126 
rect 46 126 47 127 
rect 46 127 47 128 
rect 46 138 47 139 
rect 46 139 47 140 
rect 46 140 47 141 
rect 46 141 47 142 
rect 46 142 47 143 
rect 46 143 47 144 
rect 46 154 47 155 
rect 46 155 47 156 
rect 46 156 47 157 
rect 46 157 47 158 
rect 46 158 47 159 
rect 46 159 47 160 
rect 46 170 47 171 
rect 46 171 47 172 
rect 46 172 47 173 
rect 46 173 47 174 
rect 46 174 47 175 
rect 46 175 47 176 
rect 46 186 47 187 
rect 46 187 47 188 
rect 46 188 47 189 
rect 46 189 47 190 
rect 46 190 47 191 
rect 46 191 47 192 
rect 46 202 47 203 
rect 46 203 47 204 
rect 46 204 47 205 
rect 46 205 47 206 
rect 46 206 47 207 
rect 46 207 47 208 
rect 46 218 47 219 
rect 46 219 47 220 
rect 46 220 47 221 
rect 46 221 47 222 
rect 46 222 47 223 
rect 46 223 47 224 
rect 46 234 47 235 
rect 46 235 47 236 
rect 46 236 47 237 
rect 46 237 47 238 
rect 46 238 47 239 
rect 46 239 47 240 
rect 46 250 47 251 
rect 46 251 47 252 
rect 46 252 47 253 
rect 46 253 47 254 
rect 46 254 47 255 
rect 46 255 47 256 
rect 46 266 47 267 
rect 46 267 47 268 
rect 46 268 47 269 
rect 46 269 47 270 
rect 46 270 47 271 
rect 46 271 47 272 
rect 46 282 47 283 
rect 46 283 47 284 
rect 46 284 47 285 
rect 46 285 47 286 
rect 46 286 47 287 
rect 46 287 47 288 
rect 46 298 47 299 
rect 46 299 47 300 
rect 46 300 47 301 
rect 46 301 47 302 
rect 46 302 47 303 
rect 46 303 47 304 
rect 47 10 48 11 
rect 47 11 48 12 
rect 47 12 48 13 
rect 47 13 48 14 
rect 47 14 48 15 
rect 47 15 48 16 
rect 47 26 48 27 
rect 47 28 48 29 
rect 47 29 48 30 
rect 47 30 48 31 
rect 47 31 48 32 
rect 47 42 48 43 
rect 47 43 48 44 
rect 47 44 48 45 
rect 47 45 48 46 
rect 47 47 48 48 
rect 47 58 48 59 
rect 47 60 48 61 
rect 47 61 48 62 
rect 47 63 48 64 
rect 47 74 48 75 
rect 47 76 48 77 
rect 47 77 48 78 
rect 47 78 48 79 
rect 47 79 48 80 
rect 47 90 48 91 
rect 47 92 48 93 
rect 47 93 48 94 
rect 47 95 48 96 
rect 47 106 48 107 
rect 47 108 48 109 
rect 47 109 48 110 
rect 47 110 48 111 
rect 47 111 48 112 
rect 47 122 48 123 
rect 47 123 48 124 
rect 47 124 48 125 
rect 47 125 48 126 
rect 47 127 48 128 
rect 47 138 48 139 
rect 47 140 48 141 
rect 47 141 48 142 
rect 47 143 48 144 
rect 47 154 48 155 
rect 47 155 48 156 
rect 47 156 48 157 
rect 47 157 48 158 
rect 47 159 48 160 
rect 47 170 48 171 
rect 47 172 48 173 
rect 47 173 48 174 
rect 47 174 48 175 
rect 47 175 48 176 
rect 47 186 48 187 
rect 47 188 48 189 
rect 47 189 48 190 
rect 47 191 48 192 
rect 47 202 48 203 
rect 47 204 48 205 
rect 47 205 48 206 
rect 47 206 48 207 
rect 47 207 48 208 
rect 47 218 48 219 
rect 47 220 48 221 
rect 47 221 48 222 
rect 47 222 48 223 
rect 47 223 48 224 
rect 47 234 48 235 
rect 47 236 48 237 
rect 47 237 48 238 
rect 47 238 48 239 
rect 47 239 48 240 
rect 47 250 48 251 
rect 47 251 48 252 
rect 47 252 48 253 
rect 47 253 48 254 
rect 47 254 48 255 
rect 47 255 48 256 
rect 47 266 48 267 
rect 47 267 48 268 
rect 47 268 48 269 
rect 47 269 48 270 
rect 47 271 48 272 
rect 47 282 48 283 
rect 47 284 48 285 
rect 47 285 48 286 
rect 47 286 48 287 
rect 47 287 48 288 
rect 47 298 48 299 
rect 47 300 48 301 
rect 47 301 48 302 
rect 47 303 48 304 
rect 58 10 59 11 
rect 58 11 59 12 
rect 58 12 59 13 
rect 58 13 59 14 
rect 58 14 59 15 
rect 58 15 59 16 
rect 58 26 59 27 
rect 58 28 59 29 
rect 58 29 59 30 
rect 58 31 59 32 
rect 58 42 59 43 
rect 58 43 59 44 
rect 58 44 59 45 
rect 58 45 59 46 
rect 58 46 59 47 
rect 58 47 59 48 
rect 58 58 59 59 
rect 58 59 59 60 
rect 58 60 59 61 
rect 58 61 59 62 
rect 58 62 59 63 
rect 58 63 59 64 
rect 58 74 59 75 
rect 58 75 59 76 
rect 58 76 59 77 
rect 58 77 59 78 
rect 58 79 59 80 
rect 58 90 59 91 
rect 58 92 59 93 
rect 58 93 59 94 
rect 58 94 59 95 
rect 58 95 59 96 
rect 58 106 59 107 
rect 58 107 59 108 
rect 58 108 59 109 
rect 58 109 59 110 
rect 58 110 59 111 
rect 58 111 59 112 
rect 58 122 59 123 
rect 58 124 59 125 
rect 58 125 59 126 
rect 58 127 59 128 
rect 58 138 59 139 
rect 58 139 59 140 
rect 58 140 59 141 
rect 58 141 59 142 
rect 58 142 59 143 
rect 58 143 59 144 
rect 58 154 59 155 
rect 58 156 59 157 
rect 58 157 59 158 
rect 58 159 59 160 
rect 58 170 59 171 
rect 58 172 59 173 
rect 58 173 59 174 
rect 58 174 59 175 
rect 58 175 59 176 
rect 58 186 59 187 
rect 58 187 59 188 
rect 58 188 59 189 
rect 58 189 59 190 
rect 58 191 59 192 
rect 58 202 59 203 
rect 58 204 59 205 
rect 58 205 59 206 
rect 58 206 59 207 
rect 58 207 59 208 
rect 58 218 59 219 
rect 58 219 59 220 
rect 58 220 59 221 
rect 58 221 59 222 
rect 58 223 59 224 
rect 58 234 59 235 
rect 58 236 59 237 
rect 58 237 59 238 
rect 58 239 59 240 
rect 58 250 59 251 
rect 58 252 59 253 
rect 58 253 59 254 
rect 58 254 59 255 
rect 58 255 59 256 
rect 58 266 59 267 
rect 58 267 59 268 
rect 58 268 59 269 
rect 58 269 59 270 
rect 58 271 59 272 
rect 58 282 59 283 
rect 58 283 59 284 
rect 58 284 59 285 
rect 58 285 59 286 
rect 58 287 59 288 
rect 58 298 59 299 
rect 58 299 59 300 
rect 58 300 59 301 
rect 58 301 59 302 
rect 58 303 59 304 
rect 59 10 60 11 
rect 59 11 60 12 
rect 59 12 60 13 
rect 59 13 60 14 
rect 59 14 60 15 
rect 59 15 60 16 
rect 59 26 60 27 
rect 59 27 60 28 
rect 59 28 60 29 
rect 59 29 60 30 
rect 59 30 60 31 
rect 59 31 60 32 
rect 59 42 60 43 
rect 59 43 60 44 
rect 59 44 60 45 
rect 59 45 60 46 
rect 59 46 60 47 
rect 59 47 60 48 
rect 59 58 60 59 
rect 59 59 60 60 
rect 59 60 60 61 
rect 59 61 60 62 
rect 59 62 60 63 
rect 59 63 60 64 
rect 59 74 60 75 
rect 59 75 60 76 
rect 59 76 60 77 
rect 59 77 60 78 
rect 59 78 60 79 
rect 59 79 60 80 
rect 59 90 60 91 
rect 59 91 60 92 
rect 59 92 60 93 
rect 59 93 60 94 
rect 59 94 60 95 
rect 59 95 60 96 
rect 59 106 60 107 
rect 59 107 60 108 
rect 59 108 60 109 
rect 59 109 60 110 
rect 59 110 60 111 
rect 59 111 60 112 
rect 59 122 60 123 
rect 59 123 60 124 
rect 59 124 60 125 
rect 59 125 60 126 
rect 59 126 60 127 
rect 59 127 60 128 
rect 59 138 60 139 
rect 59 139 60 140 
rect 59 140 60 141 
rect 59 141 60 142 
rect 59 142 60 143 
rect 59 143 60 144 
rect 59 154 60 155 
rect 59 155 60 156 
rect 59 156 60 157 
rect 59 157 60 158 
rect 59 158 60 159 
rect 59 159 60 160 
rect 59 170 60 171 
rect 59 171 60 172 
rect 59 172 60 173 
rect 59 173 60 174 
rect 59 174 60 175 
rect 59 175 60 176 
rect 59 186 60 187 
rect 59 187 60 188 
rect 59 188 60 189 
rect 59 189 60 190 
rect 59 190 60 191 
rect 59 191 60 192 
rect 59 202 60 203 
rect 59 203 60 204 
rect 59 204 60 205 
rect 59 205 60 206 
rect 59 206 60 207 
rect 59 207 60 208 
rect 59 218 60 219 
rect 59 219 60 220 
rect 59 220 60 221 
rect 59 221 60 222 
rect 59 222 60 223 
rect 59 223 60 224 
rect 59 234 60 235 
rect 59 235 60 236 
rect 59 236 60 237 
rect 59 237 60 238 
rect 59 238 60 239 
rect 59 239 60 240 
rect 59 250 60 251 
rect 59 251 60 252 
rect 59 252 60 253 
rect 59 253 60 254 
rect 59 254 60 255 
rect 59 255 60 256 
rect 59 266 60 267 
rect 59 267 60 268 
rect 59 268 60 269 
rect 59 269 60 270 
rect 59 270 60 271 
rect 59 271 60 272 
rect 59 282 60 283 
rect 59 283 60 284 
rect 59 284 60 285 
rect 59 285 60 286 
rect 59 286 60 287 
rect 59 287 60 288 
rect 59 298 60 299 
rect 59 299 60 300 
rect 59 300 60 301 
rect 59 301 60 302 
rect 59 302 60 303 
rect 59 303 60 304 
rect 60 10 61 11 
rect 60 11 61 12 
rect 60 12 61 13 
rect 60 13 61 14 
rect 60 14 61 15 
rect 60 15 61 16 
rect 60 26 61 27 
rect 60 27 61 28 
rect 60 28 61 29 
rect 60 29 61 30 
rect 60 30 61 31 
rect 60 31 61 32 
rect 60 42 61 43 
rect 60 43 61 44 
rect 60 44 61 45 
rect 60 45 61 46 
rect 60 46 61 47 
rect 60 47 61 48 
rect 60 58 61 59 
rect 60 59 61 60 
rect 60 60 61 61 
rect 60 61 61 62 
rect 60 62 61 63 
rect 60 63 61 64 
rect 60 74 61 75 
rect 60 75 61 76 
rect 60 76 61 77 
rect 60 77 61 78 
rect 60 78 61 79 
rect 60 79 61 80 
rect 60 90 61 91 
rect 60 91 61 92 
rect 60 92 61 93 
rect 60 93 61 94 
rect 60 94 61 95 
rect 60 95 61 96 
rect 60 106 61 107 
rect 60 107 61 108 
rect 60 108 61 109 
rect 60 109 61 110 
rect 60 110 61 111 
rect 60 111 61 112 
rect 60 122 61 123 
rect 60 123 61 124 
rect 60 124 61 125 
rect 60 125 61 126 
rect 60 126 61 127 
rect 60 127 61 128 
rect 60 138 61 139 
rect 60 139 61 140 
rect 60 140 61 141 
rect 60 141 61 142 
rect 60 142 61 143 
rect 60 143 61 144 
rect 60 154 61 155 
rect 60 155 61 156 
rect 60 156 61 157 
rect 60 157 61 158 
rect 60 158 61 159 
rect 60 159 61 160 
rect 60 170 61 171 
rect 60 171 61 172 
rect 60 172 61 173 
rect 60 173 61 174 
rect 60 174 61 175 
rect 60 175 61 176 
rect 60 186 61 187 
rect 60 187 61 188 
rect 60 188 61 189 
rect 60 189 61 190 
rect 60 190 61 191 
rect 60 191 61 192 
rect 60 202 61 203 
rect 60 203 61 204 
rect 60 204 61 205 
rect 60 205 61 206 
rect 60 206 61 207 
rect 60 207 61 208 
rect 60 218 61 219 
rect 60 219 61 220 
rect 60 220 61 221 
rect 60 221 61 222 
rect 60 222 61 223 
rect 60 223 61 224 
rect 60 234 61 235 
rect 60 235 61 236 
rect 60 236 61 237 
rect 60 237 61 238 
rect 60 238 61 239 
rect 60 239 61 240 
rect 60 250 61 251 
rect 60 251 61 252 
rect 60 252 61 253 
rect 60 253 61 254 
rect 60 254 61 255 
rect 60 255 61 256 
rect 60 266 61 267 
rect 60 267 61 268 
rect 60 268 61 269 
rect 60 269 61 270 
rect 60 270 61 271 
rect 60 271 61 272 
rect 60 282 61 283 
rect 60 283 61 284 
rect 60 284 61 285 
rect 60 285 61 286 
rect 60 286 61 287 
rect 60 287 61 288 
rect 60 298 61 299 
rect 60 299 61 300 
rect 60 300 61 301 
rect 60 301 61 302 
rect 60 302 61 303 
rect 60 303 61 304 
rect 61 10 62 11 
rect 61 11 62 12 
rect 61 12 62 13 
rect 61 13 62 14 
rect 61 14 62 15 
rect 61 15 62 16 
rect 61 26 62 27 
rect 61 27 62 28 
rect 61 28 62 29 
rect 61 29 62 30 
rect 61 30 62 31 
rect 61 31 62 32 
rect 61 42 62 43 
rect 61 43 62 44 
rect 61 44 62 45 
rect 61 45 62 46 
rect 61 46 62 47 
rect 61 47 62 48 
rect 61 58 62 59 
rect 61 59 62 60 
rect 61 60 62 61 
rect 61 61 62 62 
rect 61 62 62 63 
rect 61 63 62 64 
rect 61 74 62 75 
rect 61 75 62 76 
rect 61 76 62 77 
rect 61 77 62 78 
rect 61 78 62 79 
rect 61 79 62 80 
rect 61 90 62 91 
rect 61 91 62 92 
rect 61 92 62 93 
rect 61 93 62 94 
rect 61 94 62 95 
rect 61 95 62 96 
rect 61 106 62 107 
rect 61 107 62 108 
rect 61 108 62 109 
rect 61 109 62 110 
rect 61 110 62 111 
rect 61 111 62 112 
rect 61 122 62 123 
rect 61 123 62 124 
rect 61 124 62 125 
rect 61 125 62 126 
rect 61 126 62 127 
rect 61 127 62 128 
rect 61 138 62 139 
rect 61 139 62 140 
rect 61 140 62 141 
rect 61 141 62 142 
rect 61 142 62 143 
rect 61 143 62 144 
rect 61 154 62 155 
rect 61 155 62 156 
rect 61 156 62 157 
rect 61 157 62 158 
rect 61 158 62 159 
rect 61 159 62 160 
rect 61 170 62 171 
rect 61 171 62 172 
rect 61 172 62 173 
rect 61 173 62 174 
rect 61 174 62 175 
rect 61 175 62 176 
rect 61 186 62 187 
rect 61 187 62 188 
rect 61 188 62 189 
rect 61 189 62 190 
rect 61 190 62 191 
rect 61 191 62 192 
rect 61 202 62 203 
rect 61 203 62 204 
rect 61 204 62 205 
rect 61 205 62 206 
rect 61 206 62 207 
rect 61 207 62 208 
rect 61 218 62 219 
rect 61 219 62 220 
rect 61 220 62 221 
rect 61 221 62 222 
rect 61 222 62 223 
rect 61 223 62 224 
rect 61 234 62 235 
rect 61 235 62 236 
rect 61 236 62 237 
rect 61 237 62 238 
rect 61 238 62 239 
rect 61 239 62 240 
rect 61 250 62 251 
rect 61 251 62 252 
rect 61 252 62 253 
rect 61 253 62 254 
rect 61 254 62 255 
rect 61 255 62 256 
rect 61 266 62 267 
rect 61 267 62 268 
rect 61 268 62 269 
rect 61 269 62 270 
rect 61 270 62 271 
rect 61 271 62 272 
rect 61 282 62 283 
rect 61 283 62 284 
rect 61 284 62 285 
rect 61 285 62 286 
rect 61 286 62 287 
rect 61 287 62 288 
rect 61 298 62 299 
rect 61 299 62 300 
rect 61 300 62 301 
rect 61 301 62 302 
rect 61 302 62 303 
rect 61 303 62 304 
rect 62 10 63 11 
rect 62 11 63 12 
rect 62 12 63 13 
rect 62 13 63 14 
rect 62 14 63 15 
rect 62 15 63 16 
rect 62 26 63 27 
rect 62 27 63 28 
rect 62 28 63 29 
rect 62 29 63 30 
rect 62 30 63 31 
rect 62 31 63 32 
rect 62 42 63 43 
rect 62 43 63 44 
rect 62 44 63 45 
rect 62 45 63 46 
rect 62 46 63 47 
rect 62 47 63 48 
rect 62 58 63 59 
rect 62 59 63 60 
rect 62 60 63 61 
rect 62 61 63 62 
rect 62 62 63 63 
rect 62 63 63 64 
rect 62 74 63 75 
rect 62 75 63 76 
rect 62 76 63 77 
rect 62 77 63 78 
rect 62 78 63 79 
rect 62 79 63 80 
rect 62 90 63 91 
rect 62 91 63 92 
rect 62 92 63 93 
rect 62 93 63 94 
rect 62 94 63 95 
rect 62 95 63 96 
rect 62 106 63 107 
rect 62 107 63 108 
rect 62 108 63 109 
rect 62 109 63 110 
rect 62 110 63 111 
rect 62 111 63 112 
rect 62 122 63 123 
rect 62 123 63 124 
rect 62 124 63 125 
rect 62 125 63 126 
rect 62 126 63 127 
rect 62 127 63 128 
rect 62 138 63 139 
rect 62 139 63 140 
rect 62 140 63 141 
rect 62 141 63 142 
rect 62 142 63 143 
rect 62 143 63 144 
rect 62 154 63 155 
rect 62 155 63 156 
rect 62 156 63 157 
rect 62 157 63 158 
rect 62 158 63 159 
rect 62 159 63 160 
rect 62 170 63 171 
rect 62 171 63 172 
rect 62 172 63 173 
rect 62 173 63 174 
rect 62 174 63 175 
rect 62 175 63 176 
rect 62 186 63 187 
rect 62 187 63 188 
rect 62 188 63 189 
rect 62 189 63 190 
rect 62 190 63 191 
rect 62 191 63 192 
rect 62 202 63 203 
rect 62 203 63 204 
rect 62 204 63 205 
rect 62 205 63 206 
rect 62 206 63 207 
rect 62 207 63 208 
rect 62 218 63 219 
rect 62 219 63 220 
rect 62 220 63 221 
rect 62 221 63 222 
rect 62 222 63 223 
rect 62 223 63 224 
rect 62 234 63 235 
rect 62 235 63 236 
rect 62 236 63 237 
rect 62 237 63 238 
rect 62 238 63 239 
rect 62 239 63 240 
rect 62 250 63 251 
rect 62 251 63 252 
rect 62 252 63 253 
rect 62 253 63 254 
rect 62 254 63 255 
rect 62 255 63 256 
rect 62 266 63 267 
rect 62 267 63 268 
rect 62 268 63 269 
rect 62 269 63 270 
rect 62 270 63 271 
rect 62 271 63 272 
rect 62 282 63 283 
rect 62 283 63 284 
rect 62 284 63 285 
rect 62 285 63 286 
rect 62 286 63 287 
rect 62 287 63 288 
rect 62 298 63 299 
rect 62 299 63 300 
rect 62 300 63 301 
rect 62 301 63 302 
rect 62 302 63 303 
rect 62 303 63 304 
rect 63 10 64 11 
rect 63 12 64 13 
rect 63 13 64 14 
rect 63 14 64 15 
rect 63 15 64 16 
rect 63 26 64 27 
rect 63 27 64 28 
rect 63 28 64 29 
rect 63 29 64 30 
rect 63 30 64 31 
rect 63 31 64 32 
rect 63 42 64 43 
rect 63 44 64 45 
rect 63 45 64 46 
rect 63 46 64 47 
rect 63 47 64 48 
rect 63 58 64 59 
rect 63 59 64 60 
rect 63 60 64 61 
rect 63 61 64 62 
rect 63 63 64 64 
rect 63 74 64 75 
rect 63 75 64 76 
rect 63 76 64 77 
rect 63 77 64 78 
rect 63 78 64 79 
rect 63 79 64 80 
rect 63 90 64 91 
rect 63 91 64 92 
rect 63 92 64 93 
rect 63 93 64 94 
rect 63 94 64 95 
rect 63 95 64 96 
rect 63 106 64 107 
rect 63 108 64 109 
rect 63 109 64 110 
rect 63 111 64 112 
rect 63 122 64 123 
rect 63 124 64 125 
rect 63 125 64 126 
rect 63 126 64 127 
rect 63 127 64 128 
rect 63 138 64 139 
rect 63 140 64 141 
rect 63 141 64 142 
rect 63 143 64 144 
rect 63 154 64 155 
rect 63 155 64 156 
rect 63 156 64 157 
rect 63 157 64 158 
rect 63 158 64 159 
rect 63 159 64 160 
rect 63 170 64 171 
rect 63 171 64 172 
rect 63 172 64 173 
rect 63 173 64 174 
rect 63 175 64 176 
rect 63 186 64 187 
rect 63 188 64 189 
rect 63 189 64 190 
rect 63 190 64 191 
rect 63 191 64 192 
rect 63 202 64 203 
rect 63 203 64 204 
rect 63 204 64 205 
rect 63 205 64 206 
rect 63 207 64 208 
rect 63 218 64 219 
rect 63 220 64 221 
rect 63 221 64 222 
rect 63 223 64 224 
rect 63 234 64 235 
rect 63 235 64 236 
rect 63 236 64 237 
rect 63 237 64 238 
rect 63 238 64 239 
rect 63 239 64 240 
rect 63 250 64 251 
rect 63 252 64 253 
rect 63 253 64 254 
rect 63 254 64 255 
rect 63 255 64 256 
rect 63 266 64 267 
rect 63 268 64 269 
rect 63 269 64 270 
rect 63 270 64 271 
rect 63 271 64 272 
rect 63 282 64 283 
rect 63 284 64 285 
rect 63 285 64 286 
rect 63 286 64 287 
rect 63 287 64 288 
rect 63 298 64 299 
rect 63 299 64 300 
rect 63 300 64 301 
rect 63 301 64 302 
rect 63 302 64 303 
rect 63 303 64 304 
rect 74 10 75 11 
rect 74 11 75 12 
rect 74 12 75 13 
rect 74 13 75 14 
rect 74 15 75 16 
rect 74 26 75 27 
rect 74 27 75 28 
rect 74 28 75 29 
rect 74 29 75 30 
rect 74 30 75 31 
rect 74 31 75 32 
rect 74 42 75 43 
rect 74 43 75 44 
rect 74 44 75 45 
rect 74 45 75 46 
rect 74 46 75 47 
rect 74 47 75 48 
rect 74 58 75 59 
rect 74 60 75 61 
rect 74 61 75 62 
rect 74 62 75 63 
rect 74 63 75 64 
rect 74 74 75 75 
rect 74 75 75 76 
rect 74 76 75 77 
rect 74 77 75 78 
rect 74 79 75 80 
rect 74 90 75 91 
rect 74 91 75 92 
rect 74 92 75 93 
rect 74 93 75 94 
rect 74 95 75 96 
rect 74 106 75 107 
rect 74 108 75 109 
rect 74 109 75 110 
rect 74 111 75 112 
rect 74 122 75 123 
rect 74 124 75 125 
rect 74 125 75 126 
rect 74 127 75 128 
rect 74 138 75 139 
rect 74 140 75 141 
rect 74 141 75 142 
rect 74 143 75 144 
rect 74 154 75 155 
rect 74 155 75 156 
rect 74 156 75 157 
rect 74 157 75 158 
rect 74 159 75 160 
rect 74 170 75 171 
rect 74 171 75 172 
rect 74 172 75 173 
rect 74 173 75 174 
rect 74 175 75 176 
rect 74 186 75 187 
rect 74 188 75 189 
rect 74 189 75 190 
rect 74 191 75 192 
rect 74 202 75 203 
rect 74 203 75 204 
rect 74 204 75 205 
rect 74 205 75 206 
rect 74 206 75 207 
rect 74 207 75 208 
rect 74 218 75 219 
rect 74 220 75 221 
rect 74 221 75 222 
rect 74 223 75 224 
rect 74 234 75 235 
rect 74 235 75 236 
rect 74 236 75 237 
rect 74 237 75 238 
rect 74 239 75 240 
rect 74 250 75 251 
rect 74 252 75 253 
rect 74 253 75 254 
rect 74 254 75 255 
rect 74 255 75 256 
rect 74 266 75 267 
rect 74 268 75 269 
rect 74 269 75 270 
rect 74 271 75 272 
rect 74 282 75 283 
rect 74 284 75 285 
rect 74 285 75 286 
rect 74 286 75 287 
rect 74 287 75 288 
rect 74 298 75 299 
rect 74 299 75 300 
rect 74 300 75 301 
rect 74 301 75 302 
rect 74 303 75 304 
rect 75 10 76 11 
rect 75 11 76 12 
rect 75 12 76 13 
rect 75 13 76 14 
rect 75 14 76 15 
rect 75 15 76 16 
rect 75 26 76 27 
rect 75 27 76 28 
rect 75 28 76 29 
rect 75 29 76 30 
rect 75 30 76 31 
rect 75 31 76 32 
rect 75 42 76 43 
rect 75 43 76 44 
rect 75 44 76 45 
rect 75 45 76 46 
rect 75 46 76 47 
rect 75 47 76 48 
rect 75 58 76 59 
rect 75 59 76 60 
rect 75 60 76 61 
rect 75 61 76 62 
rect 75 62 76 63 
rect 75 63 76 64 
rect 75 74 76 75 
rect 75 75 76 76 
rect 75 76 76 77 
rect 75 77 76 78 
rect 75 78 76 79 
rect 75 79 76 80 
rect 75 90 76 91 
rect 75 91 76 92 
rect 75 92 76 93 
rect 75 93 76 94 
rect 75 94 76 95 
rect 75 95 76 96 
rect 75 106 76 107 
rect 75 107 76 108 
rect 75 108 76 109 
rect 75 109 76 110 
rect 75 110 76 111 
rect 75 111 76 112 
rect 75 122 76 123 
rect 75 123 76 124 
rect 75 124 76 125 
rect 75 125 76 126 
rect 75 126 76 127 
rect 75 127 76 128 
rect 75 138 76 139 
rect 75 139 76 140 
rect 75 140 76 141 
rect 75 141 76 142 
rect 75 142 76 143 
rect 75 143 76 144 
rect 75 154 76 155 
rect 75 155 76 156 
rect 75 156 76 157 
rect 75 157 76 158 
rect 75 158 76 159 
rect 75 159 76 160 
rect 75 170 76 171 
rect 75 171 76 172 
rect 75 172 76 173 
rect 75 173 76 174 
rect 75 174 76 175 
rect 75 175 76 176 
rect 75 186 76 187 
rect 75 187 76 188 
rect 75 188 76 189 
rect 75 189 76 190 
rect 75 190 76 191 
rect 75 191 76 192 
rect 75 202 76 203 
rect 75 203 76 204 
rect 75 204 76 205 
rect 75 205 76 206 
rect 75 206 76 207 
rect 75 207 76 208 
rect 75 218 76 219 
rect 75 219 76 220 
rect 75 220 76 221 
rect 75 221 76 222 
rect 75 222 76 223 
rect 75 223 76 224 
rect 75 234 76 235 
rect 75 235 76 236 
rect 75 236 76 237 
rect 75 237 76 238 
rect 75 238 76 239 
rect 75 239 76 240 
rect 75 250 76 251 
rect 75 251 76 252 
rect 75 252 76 253 
rect 75 253 76 254 
rect 75 254 76 255 
rect 75 255 76 256 
rect 75 266 76 267 
rect 75 267 76 268 
rect 75 268 76 269 
rect 75 269 76 270 
rect 75 270 76 271 
rect 75 271 76 272 
rect 75 282 76 283 
rect 75 283 76 284 
rect 75 284 76 285 
rect 75 285 76 286 
rect 75 286 76 287 
rect 75 287 76 288 
rect 75 298 76 299 
rect 75 299 76 300 
rect 75 300 76 301 
rect 75 301 76 302 
rect 75 302 76 303 
rect 75 303 76 304 
rect 76 10 77 11 
rect 76 11 77 12 
rect 76 12 77 13 
rect 76 13 77 14 
rect 76 14 77 15 
rect 76 15 77 16 
rect 76 26 77 27 
rect 76 27 77 28 
rect 76 28 77 29 
rect 76 29 77 30 
rect 76 30 77 31 
rect 76 31 77 32 
rect 76 42 77 43 
rect 76 43 77 44 
rect 76 44 77 45 
rect 76 45 77 46 
rect 76 46 77 47 
rect 76 47 77 48 
rect 76 58 77 59 
rect 76 59 77 60 
rect 76 60 77 61 
rect 76 61 77 62 
rect 76 62 77 63 
rect 76 63 77 64 
rect 76 74 77 75 
rect 76 75 77 76 
rect 76 76 77 77 
rect 76 77 77 78 
rect 76 78 77 79 
rect 76 79 77 80 
rect 76 90 77 91 
rect 76 91 77 92 
rect 76 92 77 93 
rect 76 93 77 94 
rect 76 94 77 95 
rect 76 95 77 96 
rect 76 106 77 107 
rect 76 107 77 108 
rect 76 108 77 109 
rect 76 109 77 110 
rect 76 110 77 111 
rect 76 111 77 112 
rect 76 122 77 123 
rect 76 123 77 124 
rect 76 124 77 125 
rect 76 125 77 126 
rect 76 126 77 127 
rect 76 127 77 128 
rect 76 138 77 139 
rect 76 139 77 140 
rect 76 140 77 141 
rect 76 141 77 142 
rect 76 142 77 143 
rect 76 143 77 144 
rect 76 154 77 155 
rect 76 155 77 156 
rect 76 156 77 157 
rect 76 157 77 158 
rect 76 158 77 159 
rect 76 159 77 160 
rect 76 170 77 171 
rect 76 171 77 172 
rect 76 172 77 173 
rect 76 173 77 174 
rect 76 174 77 175 
rect 76 175 77 176 
rect 76 186 77 187 
rect 76 187 77 188 
rect 76 188 77 189 
rect 76 189 77 190 
rect 76 190 77 191 
rect 76 191 77 192 
rect 76 202 77 203 
rect 76 203 77 204 
rect 76 204 77 205 
rect 76 205 77 206 
rect 76 206 77 207 
rect 76 207 77 208 
rect 76 218 77 219 
rect 76 219 77 220 
rect 76 220 77 221 
rect 76 221 77 222 
rect 76 222 77 223 
rect 76 223 77 224 
rect 76 234 77 235 
rect 76 235 77 236 
rect 76 236 77 237 
rect 76 237 77 238 
rect 76 238 77 239 
rect 76 239 77 240 
rect 76 250 77 251 
rect 76 251 77 252 
rect 76 252 77 253 
rect 76 253 77 254 
rect 76 254 77 255 
rect 76 255 77 256 
rect 76 266 77 267 
rect 76 267 77 268 
rect 76 268 77 269 
rect 76 269 77 270 
rect 76 270 77 271 
rect 76 271 77 272 
rect 76 282 77 283 
rect 76 283 77 284 
rect 76 284 77 285 
rect 76 285 77 286 
rect 76 286 77 287 
rect 76 287 77 288 
rect 76 298 77 299 
rect 76 299 77 300 
rect 76 300 77 301 
rect 76 301 77 302 
rect 76 302 77 303 
rect 76 303 77 304 
rect 77 10 78 11 
rect 77 11 78 12 
rect 77 12 78 13 
rect 77 13 78 14 
rect 77 14 78 15 
rect 77 15 78 16 
rect 77 26 78 27 
rect 77 27 78 28 
rect 77 28 78 29 
rect 77 29 78 30 
rect 77 30 78 31 
rect 77 31 78 32 
rect 77 42 78 43 
rect 77 43 78 44 
rect 77 44 78 45 
rect 77 45 78 46 
rect 77 46 78 47 
rect 77 47 78 48 
rect 77 58 78 59 
rect 77 59 78 60 
rect 77 60 78 61 
rect 77 61 78 62 
rect 77 62 78 63 
rect 77 63 78 64 
rect 77 74 78 75 
rect 77 75 78 76 
rect 77 76 78 77 
rect 77 77 78 78 
rect 77 78 78 79 
rect 77 79 78 80 
rect 77 90 78 91 
rect 77 91 78 92 
rect 77 92 78 93 
rect 77 93 78 94 
rect 77 94 78 95 
rect 77 95 78 96 
rect 77 106 78 107 
rect 77 107 78 108 
rect 77 108 78 109 
rect 77 109 78 110 
rect 77 110 78 111 
rect 77 111 78 112 
rect 77 122 78 123 
rect 77 123 78 124 
rect 77 124 78 125 
rect 77 125 78 126 
rect 77 126 78 127 
rect 77 127 78 128 
rect 77 138 78 139 
rect 77 139 78 140 
rect 77 140 78 141 
rect 77 141 78 142 
rect 77 142 78 143 
rect 77 143 78 144 
rect 77 154 78 155 
rect 77 155 78 156 
rect 77 156 78 157 
rect 77 157 78 158 
rect 77 158 78 159 
rect 77 159 78 160 
rect 77 170 78 171 
rect 77 171 78 172 
rect 77 172 78 173 
rect 77 173 78 174 
rect 77 174 78 175 
rect 77 175 78 176 
rect 77 186 78 187 
rect 77 187 78 188 
rect 77 188 78 189 
rect 77 189 78 190 
rect 77 190 78 191 
rect 77 191 78 192 
rect 77 202 78 203 
rect 77 203 78 204 
rect 77 204 78 205 
rect 77 205 78 206 
rect 77 206 78 207 
rect 77 207 78 208 
rect 77 218 78 219 
rect 77 219 78 220 
rect 77 220 78 221 
rect 77 221 78 222 
rect 77 222 78 223 
rect 77 223 78 224 
rect 77 234 78 235 
rect 77 235 78 236 
rect 77 236 78 237 
rect 77 237 78 238 
rect 77 238 78 239 
rect 77 239 78 240 
rect 77 250 78 251 
rect 77 251 78 252 
rect 77 252 78 253 
rect 77 253 78 254 
rect 77 254 78 255 
rect 77 255 78 256 
rect 77 266 78 267 
rect 77 267 78 268 
rect 77 268 78 269 
rect 77 269 78 270 
rect 77 270 78 271 
rect 77 271 78 272 
rect 77 282 78 283 
rect 77 283 78 284 
rect 77 284 78 285 
rect 77 285 78 286 
rect 77 286 78 287 
rect 77 287 78 288 
rect 77 298 78 299 
rect 77 299 78 300 
rect 77 300 78 301 
rect 77 301 78 302 
rect 77 302 78 303 
rect 77 303 78 304 
rect 78 10 79 11 
rect 78 11 79 12 
rect 78 12 79 13 
rect 78 13 79 14 
rect 78 14 79 15 
rect 78 15 79 16 
rect 78 26 79 27 
rect 78 27 79 28 
rect 78 28 79 29 
rect 78 29 79 30 
rect 78 30 79 31 
rect 78 31 79 32 
rect 78 42 79 43 
rect 78 43 79 44 
rect 78 44 79 45 
rect 78 45 79 46 
rect 78 46 79 47 
rect 78 47 79 48 
rect 78 58 79 59 
rect 78 59 79 60 
rect 78 60 79 61 
rect 78 61 79 62 
rect 78 62 79 63 
rect 78 63 79 64 
rect 78 74 79 75 
rect 78 75 79 76 
rect 78 76 79 77 
rect 78 77 79 78 
rect 78 78 79 79 
rect 78 79 79 80 
rect 78 90 79 91 
rect 78 91 79 92 
rect 78 92 79 93 
rect 78 93 79 94 
rect 78 94 79 95 
rect 78 95 79 96 
rect 78 106 79 107 
rect 78 107 79 108 
rect 78 108 79 109 
rect 78 109 79 110 
rect 78 110 79 111 
rect 78 111 79 112 
rect 78 122 79 123 
rect 78 123 79 124 
rect 78 124 79 125 
rect 78 125 79 126 
rect 78 126 79 127 
rect 78 127 79 128 
rect 78 138 79 139 
rect 78 139 79 140 
rect 78 140 79 141 
rect 78 141 79 142 
rect 78 142 79 143 
rect 78 143 79 144 
rect 78 154 79 155 
rect 78 155 79 156 
rect 78 156 79 157 
rect 78 157 79 158 
rect 78 158 79 159 
rect 78 159 79 160 
rect 78 170 79 171 
rect 78 171 79 172 
rect 78 172 79 173 
rect 78 173 79 174 
rect 78 174 79 175 
rect 78 175 79 176 
rect 78 186 79 187 
rect 78 187 79 188 
rect 78 188 79 189 
rect 78 189 79 190 
rect 78 190 79 191 
rect 78 191 79 192 
rect 78 202 79 203 
rect 78 203 79 204 
rect 78 204 79 205 
rect 78 205 79 206 
rect 78 206 79 207 
rect 78 207 79 208 
rect 78 218 79 219 
rect 78 219 79 220 
rect 78 220 79 221 
rect 78 221 79 222 
rect 78 222 79 223 
rect 78 223 79 224 
rect 78 234 79 235 
rect 78 235 79 236 
rect 78 236 79 237 
rect 78 237 79 238 
rect 78 238 79 239 
rect 78 239 79 240 
rect 78 250 79 251 
rect 78 251 79 252 
rect 78 252 79 253 
rect 78 253 79 254 
rect 78 254 79 255 
rect 78 255 79 256 
rect 78 266 79 267 
rect 78 267 79 268 
rect 78 268 79 269 
rect 78 269 79 270 
rect 78 270 79 271 
rect 78 271 79 272 
rect 78 282 79 283 
rect 78 283 79 284 
rect 78 284 79 285 
rect 78 285 79 286 
rect 78 286 79 287 
rect 78 287 79 288 
rect 78 298 79 299 
rect 78 299 79 300 
rect 78 300 79 301 
rect 78 301 79 302 
rect 78 302 79 303 
rect 78 303 79 304 
rect 79 10 80 11 
rect 79 11 80 12 
rect 79 12 80 13 
rect 79 13 80 14 
rect 79 14 80 15 
rect 79 15 80 16 
rect 79 26 80 27 
rect 79 28 80 29 
rect 79 29 80 30 
rect 79 30 80 31 
rect 79 31 80 32 
rect 79 42 80 43 
rect 79 43 80 44 
rect 79 44 80 45 
rect 79 45 80 46 
rect 79 47 80 48 
rect 79 58 80 59 
rect 79 59 80 60 
rect 79 60 80 61 
rect 79 61 80 62 
rect 79 63 80 64 
rect 79 74 80 75 
rect 79 76 80 77 
rect 79 77 80 78 
rect 79 78 80 79 
rect 79 79 80 80 
rect 79 90 80 91 
rect 79 92 80 93 
rect 79 93 80 94 
rect 79 95 80 96 
rect 79 106 80 107 
rect 79 107 80 108 
rect 79 108 80 109 
rect 79 109 80 110 
rect 79 110 80 111 
rect 79 111 80 112 
rect 79 122 80 123 
rect 79 123 80 124 
rect 79 124 80 125 
rect 79 125 80 126 
rect 79 127 80 128 
rect 79 138 80 139 
rect 79 140 80 141 
rect 79 141 80 142 
rect 79 143 80 144 
rect 79 154 80 155 
rect 79 156 80 157 
rect 79 157 80 158 
rect 79 159 80 160 
rect 79 170 80 171 
rect 79 172 80 173 
rect 79 173 80 174 
rect 79 174 80 175 
rect 79 175 80 176 
rect 79 186 80 187 
rect 79 188 80 189 
rect 79 189 80 190 
rect 79 190 80 191 
rect 79 191 80 192 
rect 79 202 80 203 
rect 79 203 80 204 
rect 79 204 80 205 
rect 79 205 80 206 
rect 79 207 80 208 
rect 79 218 80 219 
rect 79 219 80 220 
rect 79 220 80 221 
rect 79 221 80 222 
rect 79 222 80 223 
rect 79 223 80 224 
rect 79 234 80 235 
rect 79 235 80 236 
rect 79 236 80 237 
rect 79 237 80 238 
rect 79 239 80 240 
rect 79 250 80 251 
rect 79 251 80 252 
rect 79 252 80 253 
rect 79 253 80 254 
rect 79 255 80 256 
rect 79 266 80 267 
rect 79 267 80 268 
rect 79 268 80 269 
rect 79 269 80 270 
rect 79 270 80 271 
rect 79 271 80 272 
rect 79 282 80 283 
rect 79 284 80 285 
rect 79 285 80 286 
rect 79 287 80 288 
rect 79 298 80 299 
rect 79 299 80 300 
rect 79 300 80 301 
rect 79 301 80 302 
rect 79 303 80 304 
rect 90 10 91 11 
rect 90 11 91 12 
rect 90 12 91 13 
rect 90 13 91 14 
rect 90 14 91 15 
rect 90 15 91 16 
rect 90 26 91 27 
rect 90 27 91 28 
rect 90 28 91 29 
rect 90 29 91 30 
rect 90 30 91 31 
rect 90 31 91 32 
rect 90 42 91 43 
rect 90 44 91 45 
rect 90 45 91 46 
rect 90 47 91 48 
rect 90 58 91 59 
rect 90 60 91 61 
rect 90 61 91 62 
rect 90 63 91 64 
rect 90 74 91 75 
rect 90 76 91 77 
rect 90 77 91 78 
rect 90 79 91 80 
rect 90 90 91 91 
rect 90 92 91 93 
rect 90 93 91 94 
rect 90 95 91 96 
rect 90 106 91 107 
rect 90 107 91 108 
rect 90 108 91 109 
rect 90 109 91 110 
rect 90 111 91 112 
rect 90 122 91 123 
rect 90 123 91 124 
rect 90 124 91 125 
rect 90 125 91 126 
rect 90 127 91 128 
rect 90 138 91 139 
rect 90 140 91 141 
rect 90 141 91 142 
rect 90 143 91 144 
rect 90 154 91 155 
rect 90 156 91 157 
rect 90 157 91 158 
rect 90 159 91 160 
rect 90 170 91 171 
rect 90 171 91 172 
rect 90 172 91 173 
rect 90 173 91 174 
rect 90 175 91 176 
rect 90 186 91 187 
rect 90 188 91 189 
rect 90 189 91 190 
rect 90 190 91 191 
rect 90 191 91 192 
rect 90 202 91 203 
rect 90 203 91 204 
rect 90 204 91 205 
rect 90 205 91 206 
rect 90 206 91 207 
rect 90 207 91 208 
rect 90 218 91 219 
rect 90 219 91 220 
rect 90 220 91 221 
rect 90 221 91 222 
rect 90 223 91 224 
rect 90 234 91 235 
rect 90 236 91 237 
rect 90 237 91 238 
rect 90 239 91 240 
rect 90 250 91 251 
rect 90 251 91 252 
rect 90 252 91 253 
rect 90 253 91 254 
rect 90 255 91 256 
rect 90 266 91 267 
rect 90 268 91 269 
rect 90 269 91 270 
rect 90 270 91 271 
rect 90 271 91 272 
rect 90 282 91 283 
rect 90 283 91 284 
rect 90 284 91 285 
rect 90 285 91 286 
rect 90 286 91 287 
rect 90 287 91 288 
rect 90 298 91 299 
rect 90 299 91 300 
rect 90 300 91 301 
rect 90 301 91 302 
rect 90 302 91 303 
rect 90 303 91 304 
rect 91 10 92 11 
rect 91 11 92 12 
rect 91 12 92 13 
rect 91 13 92 14 
rect 91 14 92 15 
rect 91 15 92 16 
rect 91 26 92 27 
rect 91 27 92 28 
rect 91 28 92 29 
rect 91 29 92 30 
rect 91 30 92 31 
rect 91 31 92 32 
rect 91 42 92 43 
rect 91 43 92 44 
rect 91 44 92 45 
rect 91 45 92 46 
rect 91 46 92 47 
rect 91 47 92 48 
rect 91 58 92 59 
rect 91 59 92 60 
rect 91 60 92 61 
rect 91 61 92 62 
rect 91 62 92 63 
rect 91 63 92 64 
rect 91 74 92 75 
rect 91 75 92 76 
rect 91 76 92 77 
rect 91 77 92 78 
rect 91 78 92 79 
rect 91 79 92 80 
rect 91 90 92 91 
rect 91 91 92 92 
rect 91 92 92 93 
rect 91 93 92 94 
rect 91 94 92 95 
rect 91 95 92 96 
rect 91 106 92 107 
rect 91 107 92 108 
rect 91 108 92 109 
rect 91 109 92 110 
rect 91 110 92 111 
rect 91 111 92 112 
rect 91 122 92 123 
rect 91 123 92 124 
rect 91 124 92 125 
rect 91 125 92 126 
rect 91 126 92 127 
rect 91 127 92 128 
rect 91 138 92 139 
rect 91 139 92 140 
rect 91 140 92 141 
rect 91 141 92 142 
rect 91 142 92 143 
rect 91 143 92 144 
rect 91 154 92 155 
rect 91 155 92 156 
rect 91 156 92 157 
rect 91 157 92 158 
rect 91 158 92 159 
rect 91 159 92 160 
rect 91 170 92 171 
rect 91 171 92 172 
rect 91 172 92 173 
rect 91 173 92 174 
rect 91 174 92 175 
rect 91 175 92 176 
rect 91 186 92 187 
rect 91 187 92 188 
rect 91 188 92 189 
rect 91 189 92 190 
rect 91 190 92 191 
rect 91 191 92 192 
rect 91 202 92 203 
rect 91 203 92 204 
rect 91 204 92 205 
rect 91 205 92 206 
rect 91 206 92 207 
rect 91 207 92 208 
rect 91 218 92 219 
rect 91 219 92 220 
rect 91 220 92 221 
rect 91 221 92 222 
rect 91 222 92 223 
rect 91 223 92 224 
rect 91 234 92 235 
rect 91 235 92 236 
rect 91 236 92 237 
rect 91 237 92 238 
rect 91 238 92 239 
rect 91 239 92 240 
rect 91 250 92 251 
rect 91 251 92 252 
rect 91 252 92 253 
rect 91 253 92 254 
rect 91 254 92 255 
rect 91 255 92 256 
rect 91 266 92 267 
rect 91 267 92 268 
rect 91 268 92 269 
rect 91 269 92 270 
rect 91 270 92 271 
rect 91 271 92 272 
rect 91 282 92 283 
rect 91 283 92 284 
rect 91 284 92 285 
rect 91 285 92 286 
rect 91 286 92 287 
rect 91 287 92 288 
rect 91 298 92 299 
rect 91 299 92 300 
rect 91 300 92 301 
rect 91 301 92 302 
rect 91 302 92 303 
rect 91 303 92 304 
rect 92 10 93 11 
rect 92 11 93 12 
rect 92 12 93 13 
rect 92 13 93 14 
rect 92 14 93 15 
rect 92 15 93 16 
rect 92 26 93 27 
rect 92 27 93 28 
rect 92 28 93 29 
rect 92 29 93 30 
rect 92 30 93 31 
rect 92 31 93 32 
rect 92 42 93 43 
rect 92 43 93 44 
rect 92 44 93 45 
rect 92 45 93 46 
rect 92 46 93 47 
rect 92 47 93 48 
rect 92 58 93 59 
rect 92 59 93 60 
rect 92 60 93 61 
rect 92 61 93 62 
rect 92 62 93 63 
rect 92 63 93 64 
rect 92 74 93 75 
rect 92 75 93 76 
rect 92 76 93 77 
rect 92 77 93 78 
rect 92 78 93 79 
rect 92 79 93 80 
rect 92 90 93 91 
rect 92 91 93 92 
rect 92 92 93 93 
rect 92 93 93 94 
rect 92 94 93 95 
rect 92 95 93 96 
rect 92 106 93 107 
rect 92 107 93 108 
rect 92 108 93 109 
rect 92 109 93 110 
rect 92 110 93 111 
rect 92 111 93 112 
rect 92 122 93 123 
rect 92 123 93 124 
rect 92 124 93 125 
rect 92 125 93 126 
rect 92 126 93 127 
rect 92 127 93 128 
rect 92 138 93 139 
rect 92 139 93 140 
rect 92 140 93 141 
rect 92 141 93 142 
rect 92 142 93 143 
rect 92 143 93 144 
rect 92 154 93 155 
rect 92 155 93 156 
rect 92 156 93 157 
rect 92 157 93 158 
rect 92 158 93 159 
rect 92 159 93 160 
rect 92 170 93 171 
rect 92 171 93 172 
rect 92 172 93 173 
rect 92 173 93 174 
rect 92 174 93 175 
rect 92 175 93 176 
rect 92 186 93 187 
rect 92 187 93 188 
rect 92 188 93 189 
rect 92 189 93 190 
rect 92 190 93 191 
rect 92 191 93 192 
rect 92 202 93 203 
rect 92 203 93 204 
rect 92 204 93 205 
rect 92 205 93 206 
rect 92 206 93 207 
rect 92 207 93 208 
rect 92 218 93 219 
rect 92 219 93 220 
rect 92 220 93 221 
rect 92 221 93 222 
rect 92 222 93 223 
rect 92 223 93 224 
rect 92 234 93 235 
rect 92 235 93 236 
rect 92 236 93 237 
rect 92 237 93 238 
rect 92 238 93 239 
rect 92 239 93 240 
rect 92 250 93 251 
rect 92 251 93 252 
rect 92 252 93 253 
rect 92 253 93 254 
rect 92 254 93 255 
rect 92 255 93 256 
rect 92 266 93 267 
rect 92 267 93 268 
rect 92 268 93 269 
rect 92 269 93 270 
rect 92 270 93 271 
rect 92 271 93 272 
rect 92 282 93 283 
rect 92 283 93 284 
rect 92 284 93 285 
rect 92 285 93 286 
rect 92 286 93 287 
rect 92 287 93 288 
rect 92 298 93 299 
rect 92 299 93 300 
rect 92 300 93 301 
rect 92 301 93 302 
rect 92 302 93 303 
rect 92 303 93 304 
rect 93 10 94 11 
rect 93 11 94 12 
rect 93 12 94 13 
rect 93 13 94 14 
rect 93 14 94 15 
rect 93 15 94 16 
rect 93 26 94 27 
rect 93 27 94 28 
rect 93 28 94 29 
rect 93 29 94 30 
rect 93 30 94 31 
rect 93 31 94 32 
rect 93 42 94 43 
rect 93 43 94 44 
rect 93 44 94 45 
rect 93 45 94 46 
rect 93 46 94 47 
rect 93 47 94 48 
rect 93 58 94 59 
rect 93 59 94 60 
rect 93 60 94 61 
rect 93 61 94 62 
rect 93 62 94 63 
rect 93 63 94 64 
rect 93 74 94 75 
rect 93 75 94 76 
rect 93 76 94 77 
rect 93 77 94 78 
rect 93 78 94 79 
rect 93 79 94 80 
rect 93 90 94 91 
rect 93 91 94 92 
rect 93 92 94 93 
rect 93 93 94 94 
rect 93 94 94 95 
rect 93 95 94 96 
rect 93 106 94 107 
rect 93 107 94 108 
rect 93 108 94 109 
rect 93 109 94 110 
rect 93 110 94 111 
rect 93 111 94 112 
rect 93 122 94 123 
rect 93 123 94 124 
rect 93 124 94 125 
rect 93 125 94 126 
rect 93 126 94 127 
rect 93 127 94 128 
rect 93 138 94 139 
rect 93 139 94 140 
rect 93 140 94 141 
rect 93 141 94 142 
rect 93 142 94 143 
rect 93 143 94 144 
rect 93 154 94 155 
rect 93 155 94 156 
rect 93 156 94 157 
rect 93 157 94 158 
rect 93 158 94 159 
rect 93 159 94 160 
rect 93 170 94 171 
rect 93 171 94 172 
rect 93 172 94 173 
rect 93 173 94 174 
rect 93 174 94 175 
rect 93 175 94 176 
rect 93 186 94 187 
rect 93 187 94 188 
rect 93 188 94 189 
rect 93 189 94 190 
rect 93 190 94 191 
rect 93 191 94 192 
rect 93 202 94 203 
rect 93 203 94 204 
rect 93 204 94 205 
rect 93 205 94 206 
rect 93 206 94 207 
rect 93 207 94 208 
rect 93 218 94 219 
rect 93 219 94 220 
rect 93 220 94 221 
rect 93 221 94 222 
rect 93 222 94 223 
rect 93 223 94 224 
rect 93 234 94 235 
rect 93 235 94 236 
rect 93 236 94 237 
rect 93 237 94 238 
rect 93 238 94 239 
rect 93 239 94 240 
rect 93 250 94 251 
rect 93 251 94 252 
rect 93 252 94 253 
rect 93 253 94 254 
rect 93 254 94 255 
rect 93 255 94 256 
rect 93 266 94 267 
rect 93 267 94 268 
rect 93 268 94 269 
rect 93 269 94 270 
rect 93 270 94 271 
rect 93 271 94 272 
rect 93 282 94 283 
rect 93 283 94 284 
rect 93 284 94 285 
rect 93 285 94 286 
rect 93 286 94 287 
rect 93 287 94 288 
rect 93 298 94 299 
rect 93 299 94 300 
rect 93 300 94 301 
rect 93 301 94 302 
rect 93 302 94 303 
rect 93 303 94 304 
rect 94 10 95 11 
rect 94 11 95 12 
rect 94 12 95 13 
rect 94 13 95 14 
rect 94 14 95 15 
rect 94 15 95 16 
rect 94 26 95 27 
rect 94 27 95 28 
rect 94 28 95 29 
rect 94 29 95 30 
rect 94 30 95 31 
rect 94 31 95 32 
rect 94 42 95 43 
rect 94 43 95 44 
rect 94 44 95 45 
rect 94 45 95 46 
rect 94 46 95 47 
rect 94 47 95 48 
rect 94 58 95 59 
rect 94 59 95 60 
rect 94 60 95 61 
rect 94 61 95 62 
rect 94 62 95 63 
rect 94 63 95 64 
rect 94 74 95 75 
rect 94 75 95 76 
rect 94 76 95 77 
rect 94 77 95 78 
rect 94 78 95 79 
rect 94 79 95 80 
rect 94 90 95 91 
rect 94 91 95 92 
rect 94 92 95 93 
rect 94 93 95 94 
rect 94 94 95 95 
rect 94 95 95 96 
rect 94 106 95 107 
rect 94 107 95 108 
rect 94 108 95 109 
rect 94 109 95 110 
rect 94 110 95 111 
rect 94 111 95 112 
rect 94 122 95 123 
rect 94 123 95 124 
rect 94 124 95 125 
rect 94 125 95 126 
rect 94 126 95 127 
rect 94 127 95 128 
rect 94 138 95 139 
rect 94 139 95 140 
rect 94 140 95 141 
rect 94 141 95 142 
rect 94 142 95 143 
rect 94 143 95 144 
rect 94 154 95 155 
rect 94 155 95 156 
rect 94 156 95 157 
rect 94 157 95 158 
rect 94 158 95 159 
rect 94 159 95 160 
rect 94 170 95 171 
rect 94 171 95 172 
rect 94 172 95 173 
rect 94 173 95 174 
rect 94 174 95 175 
rect 94 175 95 176 
rect 94 186 95 187 
rect 94 187 95 188 
rect 94 188 95 189 
rect 94 189 95 190 
rect 94 190 95 191 
rect 94 191 95 192 
rect 94 202 95 203 
rect 94 203 95 204 
rect 94 204 95 205 
rect 94 205 95 206 
rect 94 206 95 207 
rect 94 207 95 208 
rect 94 218 95 219 
rect 94 219 95 220 
rect 94 220 95 221 
rect 94 221 95 222 
rect 94 222 95 223 
rect 94 223 95 224 
rect 94 234 95 235 
rect 94 235 95 236 
rect 94 236 95 237 
rect 94 237 95 238 
rect 94 238 95 239 
rect 94 239 95 240 
rect 94 250 95 251 
rect 94 251 95 252 
rect 94 252 95 253 
rect 94 253 95 254 
rect 94 254 95 255 
rect 94 255 95 256 
rect 94 266 95 267 
rect 94 267 95 268 
rect 94 268 95 269 
rect 94 269 95 270 
rect 94 270 95 271 
rect 94 271 95 272 
rect 94 282 95 283 
rect 94 283 95 284 
rect 94 284 95 285 
rect 94 285 95 286 
rect 94 286 95 287 
rect 94 287 95 288 
rect 94 298 95 299 
rect 94 299 95 300 
rect 94 300 95 301 
rect 94 301 95 302 
rect 94 302 95 303 
rect 94 303 95 304 
rect 95 10 96 11 
rect 95 11 96 12 
rect 95 12 96 13 
rect 95 13 96 14 
rect 95 14 96 15 
rect 95 15 96 16 
rect 95 26 96 27 
rect 95 28 96 29 
rect 95 29 96 30 
rect 95 30 96 31 
rect 95 31 96 32 
rect 95 42 96 43 
rect 95 43 96 44 
rect 95 44 96 45 
rect 95 45 96 46 
rect 95 47 96 48 
rect 95 58 96 59 
rect 95 59 96 60 
rect 95 60 96 61 
rect 95 61 96 62 
rect 95 62 96 63 
rect 95 63 96 64 
rect 95 74 96 75 
rect 95 76 96 77 
rect 95 77 96 78 
rect 95 78 96 79 
rect 95 79 96 80 
rect 95 90 96 91 
rect 95 92 96 93 
rect 95 93 96 94 
rect 95 94 96 95 
rect 95 95 96 96 
rect 95 106 96 107 
rect 95 108 96 109 
rect 95 109 96 110 
rect 95 111 96 112 
rect 95 122 96 123 
rect 95 124 96 125 
rect 95 125 96 126 
rect 95 127 96 128 
rect 95 138 96 139 
rect 95 140 96 141 
rect 95 141 96 142 
rect 95 142 96 143 
rect 95 143 96 144 
rect 95 154 96 155 
rect 95 156 96 157 
rect 95 157 96 158 
rect 95 159 96 160 
rect 95 170 96 171 
rect 95 171 96 172 
rect 95 172 96 173 
rect 95 173 96 174 
rect 95 175 96 176 
rect 95 186 96 187 
rect 95 188 96 189 
rect 95 189 96 190 
rect 95 191 96 192 
rect 95 202 96 203 
rect 95 203 96 204 
rect 95 204 96 205 
rect 95 205 96 206 
rect 95 207 96 208 
rect 95 218 96 219 
rect 95 219 96 220 
rect 95 220 96 221 
rect 95 221 96 222 
rect 95 223 96 224 
rect 95 234 96 235 
rect 95 235 96 236 
rect 95 236 96 237 
rect 95 237 96 238 
rect 95 239 96 240 
rect 95 250 96 251 
rect 95 252 96 253 
rect 95 253 96 254 
rect 95 254 96 255 
rect 95 255 96 256 
rect 95 266 96 267 
rect 95 268 96 269 
rect 95 269 96 270 
rect 95 270 96 271 
rect 95 271 96 272 
rect 95 282 96 283 
rect 95 283 96 284 
rect 95 284 96 285 
rect 95 285 96 286 
rect 95 287 96 288 
rect 95 298 96 299 
rect 95 299 96 300 
rect 95 300 96 301 
rect 95 301 96 302 
rect 95 302 96 303 
rect 95 303 96 304 
rect 106 10 107 11 
rect 106 11 107 12 
rect 106 12 107 13 
rect 106 13 107 14 
rect 106 15 107 16 
rect 106 26 107 27 
rect 106 28 107 29 
rect 106 29 107 30 
rect 106 30 107 31 
rect 106 31 107 32 
rect 106 58 107 59 
rect 106 60 107 61 
rect 106 61 107 62 
rect 106 62 107 63 
rect 106 63 107 64 
rect 106 74 107 75 
rect 106 75 107 76 
rect 106 76 107 77 
rect 106 77 107 78 
rect 106 78 107 79 
rect 106 79 107 80 
rect 106 90 107 91 
rect 106 91 107 92 
rect 106 92 107 93 
rect 106 93 107 94 
rect 106 95 107 96 
rect 106 106 107 107 
rect 106 108 107 109 
rect 106 109 107 110 
rect 106 110 107 111 
rect 106 111 107 112 
rect 106 122 107 123 
rect 106 123 107 124 
rect 106 124 107 125 
rect 106 125 107 126 
rect 106 127 107 128 
rect 106 138 107 139 
rect 106 139 107 140 
rect 106 140 107 141 
rect 106 141 107 142 
rect 106 143 107 144 
rect 106 154 107 155 
rect 106 155 107 156 
rect 106 156 107 157 
rect 106 157 107 158 
rect 106 158 107 159 
rect 106 159 107 160 
rect 106 170 107 171 
rect 106 171 107 172 
rect 106 172 107 173 
rect 106 173 107 174 
rect 106 174 107 175 
rect 106 175 107 176 
rect 106 186 107 187 
rect 106 188 107 189 
rect 106 189 107 190 
rect 106 190 107 191 
rect 106 191 107 192 
rect 106 202 107 203 
rect 106 204 107 205 
rect 106 205 107 206 
rect 106 206 107 207 
rect 106 207 107 208 
rect 106 218 107 219 
rect 106 220 107 221 
rect 106 221 107 222 
rect 106 223 107 224 
rect 106 234 107 235 
rect 106 236 107 237 
rect 106 237 107 238 
rect 106 239 107 240 
rect 106 250 107 251 
rect 106 251 107 252 
rect 106 252 107 253 
rect 106 253 107 254 
rect 106 254 107 255 
rect 106 255 107 256 
rect 106 266 107 267 
rect 106 268 107 269 
rect 106 269 107 270 
rect 106 270 107 271 
rect 106 271 107 272 
rect 106 282 107 283 
rect 106 283 107 284 
rect 106 284 107 285 
rect 106 285 107 286 
rect 106 286 107 287 
rect 106 287 107 288 
rect 106 298 107 299 
rect 106 300 107 301 
rect 106 301 107 302 
rect 106 303 107 304 
rect 107 10 108 11 
rect 107 11 108 12 
rect 107 12 108 13 
rect 107 13 108 14 
rect 107 14 108 15 
rect 107 15 108 16 
rect 107 26 108 27 
rect 107 27 108 28 
rect 107 28 108 29 
rect 107 29 108 30 
rect 107 30 108 31 
rect 107 31 108 32 
rect 107 58 108 59 
rect 107 59 108 60 
rect 107 60 108 61 
rect 107 61 108 62 
rect 107 62 108 63 
rect 107 63 108 64 
rect 107 74 108 75 
rect 107 75 108 76 
rect 107 76 108 77 
rect 107 77 108 78 
rect 107 78 108 79 
rect 107 79 108 80 
rect 107 90 108 91 
rect 107 91 108 92 
rect 107 92 108 93 
rect 107 93 108 94 
rect 107 94 108 95 
rect 107 95 108 96 
rect 107 106 108 107 
rect 107 107 108 108 
rect 107 108 108 109 
rect 107 109 108 110 
rect 107 110 108 111 
rect 107 111 108 112 
rect 107 122 108 123 
rect 107 123 108 124 
rect 107 124 108 125 
rect 107 125 108 126 
rect 107 126 108 127 
rect 107 127 108 128 
rect 107 138 108 139 
rect 107 139 108 140 
rect 107 140 108 141 
rect 107 141 108 142 
rect 107 142 108 143 
rect 107 143 108 144 
rect 107 154 108 155 
rect 107 155 108 156 
rect 107 156 108 157 
rect 107 157 108 158 
rect 107 158 108 159 
rect 107 159 108 160 
rect 107 170 108 171 
rect 107 171 108 172 
rect 107 172 108 173 
rect 107 173 108 174 
rect 107 174 108 175 
rect 107 175 108 176 
rect 107 186 108 187 
rect 107 187 108 188 
rect 107 188 108 189 
rect 107 189 108 190 
rect 107 190 108 191 
rect 107 191 108 192 
rect 107 202 108 203 
rect 107 203 108 204 
rect 107 204 108 205 
rect 107 205 108 206 
rect 107 206 108 207 
rect 107 207 108 208 
rect 107 218 108 219 
rect 107 219 108 220 
rect 107 220 108 221 
rect 107 221 108 222 
rect 107 222 108 223 
rect 107 223 108 224 
rect 107 234 108 235 
rect 107 235 108 236 
rect 107 236 108 237 
rect 107 237 108 238 
rect 107 238 108 239 
rect 107 239 108 240 
rect 107 250 108 251 
rect 107 251 108 252 
rect 107 252 108 253 
rect 107 253 108 254 
rect 107 254 108 255 
rect 107 255 108 256 
rect 107 266 108 267 
rect 107 267 108 268 
rect 107 268 108 269 
rect 107 269 108 270 
rect 107 270 108 271 
rect 107 271 108 272 
rect 107 282 108 283 
rect 107 283 108 284 
rect 107 284 108 285 
rect 107 285 108 286 
rect 107 286 108 287 
rect 107 287 108 288 
rect 107 298 108 299 
rect 107 299 108 300 
rect 107 300 108 301 
rect 107 301 108 302 
rect 107 302 108 303 
rect 107 303 108 304 
rect 108 10 109 11 
rect 108 11 109 12 
rect 108 12 109 13 
rect 108 13 109 14 
rect 108 14 109 15 
rect 108 15 109 16 
rect 108 26 109 27 
rect 108 27 109 28 
rect 108 28 109 29 
rect 108 29 109 30 
rect 108 30 109 31 
rect 108 31 109 32 
rect 108 58 109 59 
rect 108 59 109 60 
rect 108 60 109 61 
rect 108 61 109 62 
rect 108 62 109 63 
rect 108 63 109 64 
rect 108 74 109 75 
rect 108 75 109 76 
rect 108 76 109 77 
rect 108 77 109 78 
rect 108 78 109 79 
rect 108 79 109 80 
rect 108 90 109 91 
rect 108 91 109 92 
rect 108 92 109 93 
rect 108 93 109 94 
rect 108 94 109 95 
rect 108 95 109 96 
rect 108 106 109 107 
rect 108 107 109 108 
rect 108 108 109 109 
rect 108 109 109 110 
rect 108 110 109 111 
rect 108 111 109 112 
rect 108 122 109 123 
rect 108 123 109 124 
rect 108 124 109 125 
rect 108 125 109 126 
rect 108 126 109 127 
rect 108 127 109 128 
rect 108 138 109 139 
rect 108 139 109 140 
rect 108 140 109 141 
rect 108 141 109 142 
rect 108 142 109 143 
rect 108 143 109 144 
rect 108 154 109 155 
rect 108 155 109 156 
rect 108 156 109 157 
rect 108 157 109 158 
rect 108 158 109 159 
rect 108 159 109 160 
rect 108 170 109 171 
rect 108 171 109 172 
rect 108 172 109 173 
rect 108 173 109 174 
rect 108 174 109 175 
rect 108 175 109 176 
rect 108 186 109 187 
rect 108 187 109 188 
rect 108 188 109 189 
rect 108 189 109 190 
rect 108 190 109 191 
rect 108 191 109 192 
rect 108 202 109 203 
rect 108 203 109 204 
rect 108 204 109 205 
rect 108 205 109 206 
rect 108 206 109 207 
rect 108 207 109 208 
rect 108 218 109 219 
rect 108 219 109 220 
rect 108 220 109 221 
rect 108 221 109 222 
rect 108 222 109 223 
rect 108 223 109 224 
rect 108 234 109 235 
rect 108 235 109 236 
rect 108 236 109 237 
rect 108 237 109 238 
rect 108 238 109 239 
rect 108 239 109 240 
rect 108 250 109 251 
rect 108 251 109 252 
rect 108 252 109 253 
rect 108 253 109 254 
rect 108 254 109 255 
rect 108 255 109 256 
rect 108 266 109 267 
rect 108 267 109 268 
rect 108 268 109 269 
rect 108 269 109 270 
rect 108 270 109 271 
rect 108 271 109 272 
rect 108 282 109 283 
rect 108 283 109 284 
rect 108 284 109 285 
rect 108 285 109 286 
rect 108 286 109 287 
rect 108 287 109 288 
rect 108 298 109 299 
rect 108 299 109 300 
rect 108 300 109 301 
rect 108 301 109 302 
rect 108 302 109 303 
rect 108 303 109 304 
rect 109 10 110 11 
rect 109 11 110 12 
rect 109 12 110 13 
rect 109 13 110 14 
rect 109 14 110 15 
rect 109 15 110 16 
rect 109 26 110 27 
rect 109 27 110 28 
rect 109 28 110 29 
rect 109 29 110 30 
rect 109 30 110 31 
rect 109 31 110 32 
rect 109 58 110 59 
rect 109 59 110 60 
rect 109 60 110 61 
rect 109 61 110 62 
rect 109 62 110 63 
rect 109 63 110 64 
rect 109 74 110 75 
rect 109 75 110 76 
rect 109 76 110 77 
rect 109 77 110 78 
rect 109 78 110 79 
rect 109 79 110 80 
rect 109 90 110 91 
rect 109 91 110 92 
rect 109 92 110 93 
rect 109 93 110 94 
rect 109 94 110 95 
rect 109 95 110 96 
rect 109 106 110 107 
rect 109 107 110 108 
rect 109 108 110 109 
rect 109 109 110 110 
rect 109 110 110 111 
rect 109 111 110 112 
rect 109 122 110 123 
rect 109 123 110 124 
rect 109 124 110 125 
rect 109 125 110 126 
rect 109 126 110 127 
rect 109 127 110 128 
rect 109 138 110 139 
rect 109 139 110 140 
rect 109 140 110 141 
rect 109 141 110 142 
rect 109 142 110 143 
rect 109 143 110 144 
rect 109 154 110 155 
rect 109 155 110 156 
rect 109 156 110 157 
rect 109 157 110 158 
rect 109 158 110 159 
rect 109 159 110 160 
rect 109 170 110 171 
rect 109 171 110 172 
rect 109 172 110 173 
rect 109 173 110 174 
rect 109 174 110 175 
rect 109 175 110 176 
rect 109 186 110 187 
rect 109 187 110 188 
rect 109 188 110 189 
rect 109 189 110 190 
rect 109 190 110 191 
rect 109 191 110 192 
rect 109 202 110 203 
rect 109 203 110 204 
rect 109 204 110 205 
rect 109 205 110 206 
rect 109 206 110 207 
rect 109 207 110 208 
rect 109 218 110 219 
rect 109 219 110 220 
rect 109 220 110 221 
rect 109 221 110 222 
rect 109 222 110 223 
rect 109 223 110 224 
rect 109 234 110 235 
rect 109 235 110 236 
rect 109 236 110 237 
rect 109 237 110 238 
rect 109 238 110 239 
rect 109 239 110 240 
rect 109 250 110 251 
rect 109 251 110 252 
rect 109 252 110 253 
rect 109 253 110 254 
rect 109 254 110 255 
rect 109 255 110 256 
rect 109 266 110 267 
rect 109 267 110 268 
rect 109 268 110 269 
rect 109 269 110 270 
rect 109 270 110 271 
rect 109 271 110 272 
rect 109 282 110 283 
rect 109 283 110 284 
rect 109 284 110 285 
rect 109 285 110 286 
rect 109 286 110 287 
rect 109 287 110 288 
rect 109 298 110 299 
rect 109 299 110 300 
rect 109 300 110 301 
rect 109 301 110 302 
rect 109 302 110 303 
rect 109 303 110 304 
rect 110 10 111 11 
rect 110 11 111 12 
rect 110 12 111 13 
rect 110 13 111 14 
rect 110 14 111 15 
rect 110 15 111 16 
rect 110 26 111 27 
rect 110 27 111 28 
rect 110 28 111 29 
rect 110 29 111 30 
rect 110 30 111 31 
rect 110 31 111 32 
rect 110 58 111 59 
rect 110 59 111 60 
rect 110 60 111 61 
rect 110 61 111 62 
rect 110 62 111 63 
rect 110 63 111 64 
rect 110 74 111 75 
rect 110 75 111 76 
rect 110 76 111 77 
rect 110 77 111 78 
rect 110 78 111 79 
rect 110 79 111 80 
rect 110 90 111 91 
rect 110 91 111 92 
rect 110 92 111 93 
rect 110 93 111 94 
rect 110 94 111 95 
rect 110 95 111 96 
rect 110 106 111 107 
rect 110 107 111 108 
rect 110 108 111 109 
rect 110 109 111 110 
rect 110 110 111 111 
rect 110 111 111 112 
rect 110 122 111 123 
rect 110 123 111 124 
rect 110 124 111 125 
rect 110 125 111 126 
rect 110 126 111 127 
rect 110 127 111 128 
rect 110 138 111 139 
rect 110 139 111 140 
rect 110 140 111 141 
rect 110 141 111 142 
rect 110 142 111 143 
rect 110 143 111 144 
rect 110 154 111 155 
rect 110 155 111 156 
rect 110 156 111 157 
rect 110 157 111 158 
rect 110 158 111 159 
rect 110 159 111 160 
rect 110 170 111 171 
rect 110 171 111 172 
rect 110 172 111 173 
rect 110 173 111 174 
rect 110 174 111 175 
rect 110 175 111 176 
rect 110 186 111 187 
rect 110 187 111 188 
rect 110 188 111 189 
rect 110 189 111 190 
rect 110 190 111 191 
rect 110 191 111 192 
rect 110 202 111 203 
rect 110 203 111 204 
rect 110 204 111 205 
rect 110 205 111 206 
rect 110 206 111 207 
rect 110 207 111 208 
rect 110 218 111 219 
rect 110 219 111 220 
rect 110 220 111 221 
rect 110 221 111 222 
rect 110 222 111 223 
rect 110 223 111 224 
rect 110 234 111 235 
rect 110 235 111 236 
rect 110 236 111 237 
rect 110 237 111 238 
rect 110 238 111 239 
rect 110 239 111 240 
rect 110 250 111 251 
rect 110 251 111 252 
rect 110 252 111 253 
rect 110 253 111 254 
rect 110 254 111 255 
rect 110 255 111 256 
rect 110 266 111 267 
rect 110 267 111 268 
rect 110 268 111 269 
rect 110 269 111 270 
rect 110 270 111 271 
rect 110 271 111 272 
rect 110 282 111 283 
rect 110 283 111 284 
rect 110 284 111 285 
rect 110 285 111 286 
rect 110 286 111 287 
rect 110 287 111 288 
rect 110 298 111 299 
rect 110 299 111 300 
rect 110 300 111 301 
rect 110 301 111 302 
rect 110 302 111 303 
rect 110 303 111 304 
rect 111 10 112 11 
rect 111 11 112 12 
rect 111 12 112 13 
rect 111 13 112 14 
rect 111 14 112 15 
rect 111 15 112 16 
rect 111 26 112 27 
rect 111 28 112 29 
rect 111 29 112 30 
rect 111 31 112 32 
rect 111 58 112 59 
rect 111 59 112 60 
rect 111 60 112 61 
rect 111 61 112 62 
rect 111 63 112 64 
rect 111 74 112 75 
rect 111 76 112 77 
rect 111 77 112 78 
rect 111 79 112 80 
rect 111 90 112 91 
rect 111 91 112 92 
rect 111 92 112 93 
rect 111 93 112 94 
rect 111 95 112 96 
rect 111 106 112 107 
rect 111 107 112 108 
rect 111 108 112 109 
rect 111 109 112 110 
rect 111 111 112 112 
rect 111 122 112 123 
rect 111 123 112 124 
rect 111 124 112 125 
rect 111 125 112 126 
rect 111 126 112 127 
rect 111 127 112 128 
rect 111 138 112 139 
rect 111 140 112 141 
rect 111 141 112 142 
rect 111 142 112 143 
rect 111 143 112 144 
rect 111 154 112 155 
rect 111 156 112 157 
rect 111 157 112 158 
rect 111 159 112 160 
rect 111 170 112 171 
rect 111 172 112 173 
rect 111 173 112 174 
rect 111 175 112 176 
rect 111 186 112 187 
rect 111 187 112 188 
rect 111 188 112 189 
rect 111 189 112 190 
rect 111 191 112 192 
rect 111 202 112 203 
rect 111 204 112 205 
rect 111 205 112 206 
rect 111 207 112 208 
rect 111 218 112 219 
rect 111 219 112 220 
rect 111 220 112 221 
rect 111 221 112 222 
rect 111 223 112 224 
rect 111 234 112 235 
rect 111 235 112 236 
rect 111 236 112 237 
rect 111 237 112 238 
rect 111 239 112 240 
rect 111 250 112 251 
rect 111 252 112 253 
rect 111 253 112 254 
rect 111 254 112 255 
rect 111 255 112 256 
rect 111 266 112 267 
rect 111 268 112 269 
rect 111 269 112 270 
rect 111 271 112 272 
rect 111 282 112 283 
rect 111 284 112 285 
rect 111 285 112 286 
rect 111 286 112 287 
rect 111 287 112 288 
rect 111 298 112 299 
rect 111 300 112 301 
rect 111 301 112 302 
rect 111 303 112 304 
rect 122 10 123 11 
rect 122 12 123 13 
rect 122 13 123 14 
rect 122 14 123 15 
rect 122 15 123 16 
rect 122 26 123 27 
rect 122 27 123 28 
rect 122 28 123 29 
rect 122 29 123 30 
rect 122 31 123 32 
rect 122 42 123 43 
rect 122 44 123 45 
rect 122 45 123 46 
rect 122 46 123 47 
rect 122 47 123 48 
rect 122 58 123 59 
rect 122 59 123 60 
rect 122 60 123 61 
rect 122 61 123 62 
rect 122 63 123 64 
rect 122 74 123 75 
rect 122 76 123 77 
rect 122 77 123 78 
rect 122 79 123 80 
rect 122 90 123 91 
rect 122 91 123 92 
rect 122 92 123 93 
rect 122 93 123 94 
rect 122 95 123 96 
rect 122 106 123 107 
rect 122 107 123 108 
rect 122 108 123 109 
rect 122 109 123 110 
rect 122 111 123 112 
rect 122 122 123 123 
rect 122 124 123 125 
rect 122 125 123 126 
rect 122 126 123 127 
rect 122 127 123 128 
rect 122 138 123 139 
rect 122 140 123 141 
rect 122 141 123 142 
rect 122 143 123 144 
rect 122 154 123 155 
rect 122 155 123 156 
rect 122 156 123 157 
rect 122 157 123 158 
rect 122 158 123 159 
rect 122 159 123 160 
rect 122 170 123 171 
rect 122 172 123 173 
rect 122 173 123 174 
rect 122 174 123 175 
rect 122 175 123 176 
rect 122 186 123 187 
rect 122 188 123 189 
rect 122 189 123 190 
rect 122 190 123 191 
rect 122 191 123 192 
rect 122 202 123 203 
rect 122 204 123 205 
rect 122 205 123 206 
rect 122 206 123 207 
rect 122 207 123 208 
rect 122 218 123 219 
rect 122 220 123 221 
rect 122 221 123 222 
rect 122 222 123 223 
rect 122 223 123 224 
rect 122 234 123 235 
rect 122 236 123 237 
rect 122 237 123 238 
rect 122 239 123 240 
rect 122 250 123 251 
rect 122 251 123 252 
rect 122 252 123 253 
rect 122 253 123 254 
rect 122 255 123 256 
rect 122 266 123 267 
rect 122 267 123 268 
rect 122 268 123 269 
rect 122 269 123 270 
rect 122 270 123 271 
rect 122 271 123 272 
rect 122 282 123 283 
rect 122 284 123 285 
rect 122 285 123 286 
rect 122 287 123 288 
rect 122 298 123 299 
rect 122 299 123 300 
rect 122 300 123 301 
rect 122 301 123 302 
rect 122 302 123 303 
rect 122 303 123 304 
rect 123 10 124 11 
rect 123 11 124 12 
rect 123 12 124 13 
rect 123 13 124 14 
rect 123 14 124 15 
rect 123 15 124 16 
rect 123 26 124 27 
rect 123 27 124 28 
rect 123 28 124 29 
rect 123 29 124 30 
rect 123 30 124 31 
rect 123 31 124 32 
rect 123 42 124 43 
rect 123 43 124 44 
rect 123 44 124 45 
rect 123 45 124 46 
rect 123 46 124 47 
rect 123 47 124 48 
rect 123 58 124 59 
rect 123 59 124 60 
rect 123 60 124 61 
rect 123 61 124 62 
rect 123 62 124 63 
rect 123 63 124 64 
rect 123 74 124 75 
rect 123 75 124 76 
rect 123 76 124 77 
rect 123 77 124 78 
rect 123 78 124 79 
rect 123 79 124 80 
rect 123 90 124 91 
rect 123 91 124 92 
rect 123 92 124 93 
rect 123 93 124 94 
rect 123 94 124 95 
rect 123 95 124 96 
rect 123 106 124 107 
rect 123 107 124 108 
rect 123 108 124 109 
rect 123 109 124 110 
rect 123 110 124 111 
rect 123 111 124 112 
rect 123 122 124 123 
rect 123 123 124 124 
rect 123 124 124 125 
rect 123 125 124 126 
rect 123 126 124 127 
rect 123 127 124 128 
rect 123 138 124 139 
rect 123 139 124 140 
rect 123 140 124 141 
rect 123 141 124 142 
rect 123 142 124 143 
rect 123 143 124 144 
rect 123 154 124 155 
rect 123 155 124 156 
rect 123 156 124 157 
rect 123 157 124 158 
rect 123 158 124 159 
rect 123 159 124 160 
rect 123 170 124 171 
rect 123 171 124 172 
rect 123 172 124 173 
rect 123 173 124 174 
rect 123 174 124 175 
rect 123 175 124 176 
rect 123 186 124 187 
rect 123 187 124 188 
rect 123 188 124 189 
rect 123 189 124 190 
rect 123 190 124 191 
rect 123 191 124 192 
rect 123 202 124 203 
rect 123 203 124 204 
rect 123 204 124 205 
rect 123 205 124 206 
rect 123 206 124 207 
rect 123 207 124 208 
rect 123 218 124 219 
rect 123 219 124 220 
rect 123 220 124 221 
rect 123 221 124 222 
rect 123 222 124 223 
rect 123 223 124 224 
rect 123 234 124 235 
rect 123 235 124 236 
rect 123 236 124 237 
rect 123 237 124 238 
rect 123 238 124 239 
rect 123 239 124 240 
rect 123 250 124 251 
rect 123 251 124 252 
rect 123 252 124 253 
rect 123 253 124 254 
rect 123 254 124 255 
rect 123 255 124 256 
rect 123 266 124 267 
rect 123 267 124 268 
rect 123 268 124 269 
rect 123 269 124 270 
rect 123 270 124 271 
rect 123 271 124 272 
rect 123 282 124 283 
rect 123 283 124 284 
rect 123 284 124 285 
rect 123 285 124 286 
rect 123 286 124 287 
rect 123 287 124 288 
rect 123 298 124 299 
rect 123 299 124 300 
rect 123 300 124 301 
rect 123 301 124 302 
rect 123 302 124 303 
rect 123 303 124 304 
rect 124 10 125 11 
rect 124 11 125 12 
rect 124 12 125 13 
rect 124 13 125 14 
rect 124 14 125 15 
rect 124 15 125 16 
rect 124 26 125 27 
rect 124 27 125 28 
rect 124 28 125 29 
rect 124 29 125 30 
rect 124 30 125 31 
rect 124 31 125 32 
rect 124 42 125 43 
rect 124 43 125 44 
rect 124 44 125 45 
rect 124 45 125 46 
rect 124 46 125 47 
rect 124 47 125 48 
rect 124 58 125 59 
rect 124 59 125 60 
rect 124 60 125 61 
rect 124 61 125 62 
rect 124 62 125 63 
rect 124 63 125 64 
rect 124 74 125 75 
rect 124 75 125 76 
rect 124 76 125 77 
rect 124 77 125 78 
rect 124 78 125 79 
rect 124 79 125 80 
rect 124 90 125 91 
rect 124 91 125 92 
rect 124 92 125 93 
rect 124 93 125 94 
rect 124 94 125 95 
rect 124 95 125 96 
rect 124 106 125 107 
rect 124 107 125 108 
rect 124 108 125 109 
rect 124 109 125 110 
rect 124 110 125 111 
rect 124 111 125 112 
rect 124 122 125 123 
rect 124 123 125 124 
rect 124 124 125 125 
rect 124 125 125 126 
rect 124 126 125 127 
rect 124 127 125 128 
rect 124 138 125 139 
rect 124 139 125 140 
rect 124 140 125 141 
rect 124 141 125 142 
rect 124 142 125 143 
rect 124 143 125 144 
rect 124 154 125 155 
rect 124 155 125 156 
rect 124 156 125 157 
rect 124 157 125 158 
rect 124 158 125 159 
rect 124 159 125 160 
rect 124 170 125 171 
rect 124 171 125 172 
rect 124 172 125 173 
rect 124 173 125 174 
rect 124 174 125 175 
rect 124 175 125 176 
rect 124 186 125 187 
rect 124 187 125 188 
rect 124 188 125 189 
rect 124 189 125 190 
rect 124 190 125 191 
rect 124 191 125 192 
rect 124 202 125 203 
rect 124 203 125 204 
rect 124 204 125 205 
rect 124 205 125 206 
rect 124 206 125 207 
rect 124 207 125 208 
rect 124 218 125 219 
rect 124 219 125 220 
rect 124 220 125 221 
rect 124 221 125 222 
rect 124 222 125 223 
rect 124 223 125 224 
rect 124 234 125 235 
rect 124 235 125 236 
rect 124 236 125 237 
rect 124 237 125 238 
rect 124 238 125 239 
rect 124 239 125 240 
rect 124 250 125 251 
rect 124 251 125 252 
rect 124 252 125 253 
rect 124 253 125 254 
rect 124 254 125 255 
rect 124 255 125 256 
rect 124 266 125 267 
rect 124 267 125 268 
rect 124 268 125 269 
rect 124 269 125 270 
rect 124 270 125 271 
rect 124 271 125 272 
rect 124 282 125 283 
rect 124 283 125 284 
rect 124 284 125 285 
rect 124 285 125 286 
rect 124 286 125 287 
rect 124 287 125 288 
rect 124 298 125 299 
rect 124 299 125 300 
rect 124 300 125 301 
rect 124 301 125 302 
rect 124 302 125 303 
rect 124 303 125 304 
rect 125 10 126 11 
rect 125 11 126 12 
rect 125 12 126 13 
rect 125 13 126 14 
rect 125 14 126 15 
rect 125 15 126 16 
rect 125 26 126 27 
rect 125 27 126 28 
rect 125 28 126 29 
rect 125 29 126 30 
rect 125 30 126 31 
rect 125 31 126 32 
rect 125 42 126 43 
rect 125 43 126 44 
rect 125 44 126 45 
rect 125 45 126 46 
rect 125 46 126 47 
rect 125 47 126 48 
rect 125 58 126 59 
rect 125 59 126 60 
rect 125 60 126 61 
rect 125 61 126 62 
rect 125 62 126 63 
rect 125 63 126 64 
rect 125 74 126 75 
rect 125 75 126 76 
rect 125 76 126 77 
rect 125 77 126 78 
rect 125 78 126 79 
rect 125 79 126 80 
rect 125 90 126 91 
rect 125 91 126 92 
rect 125 92 126 93 
rect 125 93 126 94 
rect 125 94 126 95 
rect 125 95 126 96 
rect 125 106 126 107 
rect 125 107 126 108 
rect 125 108 126 109 
rect 125 109 126 110 
rect 125 110 126 111 
rect 125 111 126 112 
rect 125 122 126 123 
rect 125 123 126 124 
rect 125 124 126 125 
rect 125 125 126 126 
rect 125 126 126 127 
rect 125 127 126 128 
rect 125 138 126 139 
rect 125 139 126 140 
rect 125 140 126 141 
rect 125 141 126 142 
rect 125 142 126 143 
rect 125 143 126 144 
rect 125 154 126 155 
rect 125 155 126 156 
rect 125 156 126 157 
rect 125 157 126 158 
rect 125 158 126 159 
rect 125 159 126 160 
rect 125 170 126 171 
rect 125 171 126 172 
rect 125 172 126 173 
rect 125 173 126 174 
rect 125 174 126 175 
rect 125 175 126 176 
rect 125 186 126 187 
rect 125 187 126 188 
rect 125 188 126 189 
rect 125 189 126 190 
rect 125 190 126 191 
rect 125 191 126 192 
rect 125 202 126 203 
rect 125 203 126 204 
rect 125 204 126 205 
rect 125 205 126 206 
rect 125 206 126 207 
rect 125 207 126 208 
rect 125 218 126 219 
rect 125 219 126 220 
rect 125 220 126 221 
rect 125 221 126 222 
rect 125 222 126 223 
rect 125 223 126 224 
rect 125 234 126 235 
rect 125 235 126 236 
rect 125 236 126 237 
rect 125 237 126 238 
rect 125 238 126 239 
rect 125 239 126 240 
rect 125 250 126 251 
rect 125 251 126 252 
rect 125 252 126 253 
rect 125 253 126 254 
rect 125 254 126 255 
rect 125 255 126 256 
rect 125 266 126 267 
rect 125 267 126 268 
rect 125 268 126 269 
rect 125 269 126 270 
rect 125 270 126 271 
rect 125 271 126 272 
rect 125 282 126 283 
rect 125 283 126 284 
rect 125 284 126 285 
rect 125 285 126 286 
rect 125 286 126 287 
rect 125 287 126 288 
rect 125 298 126 299 
rect 125 299 126 300 
rect 125 300 126 301 
rect 125 301 126 302 
rect 125 302 126 303 
rect 125 303 126 304 
rect 126 10 127 11 
rect 126 11 127 12 
rect 126 12 127 13 
rect 126 13 127 14 
rect 126 14 127 15 
rect 126 15 127 16 
rect 126 26 127 27 
rect 126 27 127 28 
rect 126 28 127 29 
rect 126 29 127 30 
rect 126 30 127 31 
rect 126 31 127 32 
rect 126 42 127 43 
rect 126 43 127 44 
rect 126 44 127 45 
rect 126 45 127 46 
rect 126 46 127 47 
rect 126 47 127 48 
rect 126 58 127 59 
rect 126 59 127 60 
rect 126 60 127 61 
rect 126 61 127 62 
rect 126 62 127 63 
rect 126 63 127 64 
rect 126 74 127 75 
rect 126 75 127 76 
rect 126 76 127 77 
rect 126 77 127 78 
rect 126 78 127 79 
rect 126 79 127 80 
rect 126 90 127 91 
rect 126 91 127 92 
rect 126 92 127 93 
rect 126 93 127 94 
rect 126 94 127 95 
rect 126 95 127 96 
rect 126 106 127 107 
rect 126 107 127 108 
rect 126 108 127 109 
rect 126 109 127 110 
rect 126 110 127 111 
rect 126 111 127 112 
rect 126 122 127 123 
rect 126 123 127 124 
rect 126 124 127 125 
rect 126 125 127 126 
rect 126 126 127 127 
rect 126 127 127 128 
rect 126 138 127 139 
rect 126 139 127 140 
rect 126 140 127 141 
rect 126 141 127 142 
rect 126 142 127 143 
rect 126 143 127 144 
rect 126 154 127 155 
rect 126 155 127 156 
rect 126 156 127 157 
rect 126 157 127 158 
rect 126 158 127 159 
rect 126 159 127 160 
rect 126 170 127 171 
rect 126 171 127 172 
rect 126 172 127 173 
rect 126 173 127 174 
rect 126 174 127 175 
rect 126 175 127 176 
rect 126 186 127 187 
rect 126 187 127 188 
rect 126 188 127 189 
rect 126 189 127 190 
rect 126 190 127 191 
rect 126 191 127 192 
rect 126 202 127 203 
rect 126 203 127 204 
rect 126 204 127 205 
rect 126 205 127 206 
rect 126 206 127 207 
rect 126 207 127 208 
rect 126 218 127 219 
rect 126 219 127 220 
rect 126 220 127 221 
rect 126 221 127 222 
rect 126 222 127 223 
rect 126 223 127 224 
rect 126 234 127 235 
rect 126 235 127 236 
rect 126 236 127 237 
rect 126 237 127 238 
rect 126 238 127 239 
rect 126 239 127 240 
rect 126 250 127 251 
rect 126 251 127 252 
rect 126 252 127 253 
rect 126 253 127 254 
rect 126 254 127 255 
rect 126 255 127 256 
rect 126 266 127 267 
rect 126 267 127 268 
rect 126 268 127 269 
rect 126 269 127 270 
rect 126 270 127 271 
rect 126 271 127 272 
rect 126 282 127 283 
rect 126 283 127 284 
rect 126 284 127 285 
rect 126 285 127 286 
rect 126 286 127 287 
rect 126 287 127 288 
rect 126 298 127 299 
rect 126 299 127 300 
rect 126 300 127 301 
rect 126 301 127 302 
rect 126 302 127 303 
rect 126 303 127 304 
rect 127 10 128 11 
rect 127 12 128 13 
rect 127 13 128 14 
rect 127 15 128 16 
rect 127 26 128 27 
rect 127 27 128 28 
rect 127 28 128 29 
rect 127 29 128 30 
rect 127 30 128 31 
rect 127 31 128 32 
rect 127 42 128 43 
rect 127 44 128 45 
rect 127 45 128 46 
rect 127 47 128 48 
rect 127 58 128 59 
rect 127 60 128 61 
rect 127 61 128 62 
rect 127 63 128 64 
rect 127 74 128 75 
rect 127 75 128 76 
rect 127 76 128 77 
rect 127 77 128 78 
rect 127 79 128 80 
rect 127 90 128 91 
rect 127 92 128 93 
rect 127 93 128 94 
rect 127 94 128 95 
rect 127 95 128 96 
rect 127 106 128 107 
rect 127 108 128 109 
rect 127 109 128 110 
rect 127 111 128 112 
rect 127 122 128 123 
rect 127 123 128 124 
rect 127 124 128 125 
rect 127 125 128 126 
rect 127 127 128 128 
rect 127 138 128 139 
rect 127 140 128 141 
rect 127 141 128 142 
rect 127 142 128 143 
rect 127 143 128 144 
rect 127 154 128 155 
rect 127 155 128 156 
rect 127 156 128 157 
rect 127 157 128 158 
rect 127 158 128 159 
rect 127 159 128 160 
rect 127 170 128 171 
rect 127 171 128 172 
rect 127 172 128 173 
rect 127 173 128 174 
rect 127 174 128 175 
rect 127 175 128 176 
rect 127 186 128 187 
rect 127 188 128 189 
rect 127 189 128 190 
rect 127 191 128 192 
rect 127 202 128 203 
rect 127 203 128 204 
rect 127 204 128 205 
rect 127 205 128 206 
rect 127 207 128 208 
rect 127 218 128 219 
rect 127 220 128 221 
rect 127 221 128 222 
rect 127 222 128 223 
rect 127 223 128 224 
rect 127 234 128 235 
rect 127 235 128 236 
rect 127 236 128 237 
rect 127 237 128 238 
rect 127 239 128 240 
rect 127 250 128 251 
rect 127 251 128 252 
rect 127 252 128 253 
rect 127 253 128 254 
rect 127 255 128 256 
rect 127 266 128 267 
rect 127 267 128 268 
rect 127 268 128 269 
rect 127 269 128 270 
rect 127 271 128 272 
rect 127 282 128 283 
rect 127 283 128 284 
rect 127 284 128 285 
rect 127 285 128 286 
rect 127 286 128 287 
rect 127 287 128 288 
rect 127 298 128 299 
rect 127 299 128 300 
rect 127 300 128 301 
rect 127 301 128 302 
rect 127 302 128 303 
rect 127 303 128 304 
rect 138 10 139 11 
rect 138 12 139 13 
rect 138 13 139 14 
rect 138 14 139 15 
rect 138 15 139 16 
rect 138 26 139 27 
rect 138 27 139 28 
rect 138 28 139 29 
rect 138 29 139 30 
rect 138 30 139 31 
rect 138 31 139 32 
rect 138 42 139 43 
rect 138 44 139 45 
rect 138 45 139 46 
rect 138 46 139 47 
rect 138 47 139 48 
rect 138 58 139 59 
rect 138 59 139 60 
rect 138 60 139 61 
rect 138 61 139 62 
rect 138 63 139 64 
rect 138 74 139 75 
rect 138 75 139 76 
rect 138 76 139 77 
rect 138 77 139 78 
rect 138 78 139 79 
rect 138 79 139 80 
rect 138 90 139 91 
rect 138 92 139 93 
rect 138 93 139 94 
rect 138 95 139 96 
rect 138 106 139 107 
rect 138 108 139 109 
rect 138 109 139 110 
rect 138 111 139 112 
rect 138 122 139 123 
rect 138 123 139 124 
rect 138 124 139 125 
rect 138 125 139 126 
rect 138 127 139 128 
rect 138 138 139 139 
rect 138 140 139 141 
rect 138 141 139 142 
rect 138 142 139 143 
rect 138 143 139 144 
rect 138 154 139 155 
rect 138 156 139 157 
rect 138 157 139 158 
rect 138 159 139 160 
rect 138 170 139 171 
rect 138 171 139 172 
rect 138 172 139 173 
rect 138 173 139 174 
rect 138 175 139 176 
rect 138 186 139 187 
rect 138 188 139 189 
rect 138 189 139 190 
rect 138 191 139 192 
rect 138 202 139 203 
rect 138 204 139 205 
rect 138 205 139 206 
rect 138 207 139 208 
rect 138 218 139 219 
rect 138 219 139 220 
rect 138 220 139 221 
rect 138 221 139 222 
rect 138 223 139 224 
rect 138 234 139 235 
rect 138 236 139 237 
rect 138 237 139 238 
rect 138 238 139 239 
rect 138 239 139 240 
rect 138 250 139 251 
rect 138 252 139 253 
rect 138 253 139 254 
rect 138 254 139 255 
rect 138 255 139 256 
rect 138 266 139 267 
rect 138 268 139 269 
rect 138 269 139 270 
rect 138 270 139 271 
rect 138 271 139 272 
rect 138 282 139 283 
rect 138 284 139 285 
rect 138 285 139 286 
rect 138 287 139 288 
rect 138 298 139 299 
rect 138 300 139 301 
rect 138 301 139 302 
rect 138 302 139 303 
rect 138 303 139 304 
rect 139 10 140 11 
rect 139 11 140 12 
rect 139 12 140 13 
rect 139 13 140 14 
rect 139 14 140 15 
rect 139 15 140 16 
rect 139 26 140 27 
rect 139 27 140 28 
rect 139 28 140 29 
rect 139 29 140 30 
rect 139 30 140 31 
rect 139 31 140 32 
rect 139 42 140 43 
rect 139 43 140 44 
rect 139 44 140 45 
rect 139 45 140 46 
rect 139 46 140 47 
rect 139 47 140 48 
rect 139 58 140 59 
rect 139 59 140 60 
rect 139 60 140 61 
rect 139 61 140 62 
rect 139 62 140 63 
rect 139 63 140 64 
rect 139 74 140 75 
rect 139 75 140 76 
rect 139 76 140 77 
rect 139 77 140 78 
rect 139 78 140 79 
rect 139 79 140 80 
rect 139 90 140 91 
rect 139 91 140 92 
rect 139 92 140 93 
rect 139 93 140 94 
rect 139 94 140 95 
rect 139 95 140 96 
rect 139 106 140 107 
rect 139 107 140 108 
rect 139 108 140 109 
rect 139 109 140 110 
rect 139 110 140 111 
rect 139 111 140 112 
rect 139 122 140 123 
rect 139 123 140 124 
rect 139 124 140 125 
rect 139 125 140 126 
rect 139 126 140 127 
rect 139 127 140 128 
rect 139 138 140 139 
rect 139 139 140 140 
rect 139 140 140 141 
rect 139 141 140 142 
rect 139 142 140 143 
rect 139 143 140 144 
rect 139 154 140 155 
rect 139 155 140 156 
rect 139 156 140 157 
rect 139 157 140 158 
rect 139 158 140 159 
rect 139 159 140 160 
rect 139 170 140 171 
rect 139 171 140 172 
rect 139 172 140 173 
rect 139 173 140 174 
rect 139 174 140 175 
rect 139 175 140 176 
rect 139 186 140 187 
rect 139 187 140 188 
rect 139 188 140 189 
rect 139 189 140 190 
rect 139 190 140 191 
rect 139 191 140 192 
rect 139 202 140 203 
rect 139 203 140 204 
rect 139 204 140 205 
rect 139 205 140 206 
rect 139 206 140 207 
rect 139 207 140 208 
rect 139 218 140 219 
rect 139 219 140 220 
rect 139 220 140 221 
rect 139 221 140 222 
rect 139 222 140 223 
rect 139 223 140 224 
rect 139 234 140 235 
rect 139 235 140 236 
rect 139 236 140 237 
rect 139 237 140 238 
rect 139 238 140 239 
rect 139 239 140 240 
rect 139 250 140 251 
rect 139 251 140 252 
rect 139 252 140 253 
rect 139 253 140 254 
rect 139 254 140 255 
rect 139 255 140 256 
rect 139 266 140 267 
rect 139 267 140 268 
rect 139 268 140 269 
rect 139 269 140 270 
rect 139 270 140 271 
rect 139 271 140 272 
rect 139 282 140 283 
rect 139 283 140 284 
rect 139 284 140 285 
rect 139 285 140 286 
rect 139 286 140 287 
rect 139 287 140 288 
rect 139 298 140 299 
rect 139 299 140 300 
rect 139 300 140 301 
rect 139 301 140 302 
rect 139 302 140 303 
rect 139 303 140 304 
rect 140 10 141 11 
rect 140 11 141 12 
rect 140 12 141 13 
rect 140 13 141 14 
rect 140 14 141 15 
rect 140 15 141 16 
rect 140 26 141 27 
rect 140 27 141 28 
rect 140 28 141 29 
rect 140 29 141 30 
rect 140 30 141 31 
rect 140 31 141 32 
rect 140 42 141 43 
rect 140 43 141 44 
rect 140 44 141 45 
rect 140 45 141 46 
rect 140 46 141 47 
rect 140 47 141 48 
rect 140 58 141 59 
rect 140 59 141 60 
rect 140 60 141 61 
rect 140 61 141 62 
rect 140 62 141 63 
rect 140 63 141 64 
rect 140 74 141 75 
rect 140 75 141 76 
rect 140 76 141 77 
rect 140 77 141 78 
rect 140 78 141 79 
rect 140 79 141 80 
rect 140 90 141 91 
rect 140 91 141 92 
rect 140 92 141 93 
rect 140 93 141 94 
rect 140 94 141 95 
rect 140 95 141 96 
rect 140 106 141 107 
rect 140 107 141 108 
rect 140 108 141 109 
rect 140 109 141 110 
rect 140 110 141 111 
rect 140 111 141 112 
rect 140 122 141 123 
rect 140 123 141 124 
rect 140 124 141 125 
rect 140 125 141 126 
rect 140 126 141 127 
rect 140 127 141 128 
rect 140 138 141 139 
rect 140 139 141 140 
rect 140 140 141 141 
rect 140 141 141 142 
rect 140 142 141 143 
rect 140 143 141 144 
rect 140 154 141 155 
rect 140 155 141 156 
rect 140 156 141 157 
rect 140 157 141 158 
rect 140 158 141 159 
rect 140 159 141 160 
rect 140 170 141 171 
rect 140 171 141 172 
rect 140 172 141 173 
rect 140 173 141 174 
rect 140 174 141 175 
rect 140 175 141 176 
rect 140 186 141 187 
rect 140 187 141 188 
rect 140 188 141 189 
rect 140 189 141 190 
rect 140 190 141 191 
rect 140 191 141 192 
rect 140 202 141 203 
rect 140 203 141 204 
rect 140 204 141 205 
rect 140 205 141 206 
rect 140 206 141 207 
rect 140 207 141 208 
rect 140 218 141 219 
rect 140 219 141 220 
rect 140 220 141 221 
rect 140 221 141 222 
rect 140 222 141 223 
rect 140 223 141 224 
rect 140 234 141 235 
rect 140 235 141 236 
rect 140 236 141 237 
rect 140 237 141 238 
rect 140 238 141 239 
rect 140 239 141 240 
rect 140 250 141 251 
rect 140 251 141 252 
rect 140 252 141 253 
rect 140 253 141 254 
rect 140 254 141 255 
rect 140 255 141 256 
rect 140 266 141 267 
rect 140 267 141 268 
rect 140 268 141 269 
rect 140 269 141 270 
rect 140 270 141 271 
rect 140 271 141 272 
rect 140 282 141 283 
rect 140 283 141 284 
rect 140 284 141 285 
rect 140 285 141 286 
rect 140 286 141 287 
rect 140 287 141 288 
rect 140 298 141 299 
rect 140 299 141 300 
rect 140 300 141 301 
rect 140 301 141 302 
rect 140 302 141 303 
rect 140 303 141 304 
rect 141 10 142 11 
rect 141 11 142 12 
rect 141 12 142 13 
rect 141 13 142 14 
rect 141 14 142 15 
rect 141 15 142 16 
rect 141 26 142 27 
rect 141 27 142 28 
rect 141 28 142 29 
rect 141 29 142 30 
rect 141 30 142 31 
rect 141 31 142 32 
rect 141 42 142 43 
rect 141 43 142 44 
rect 141 44 142 45 
rect 141 45 142 46 
rect 141 46 142 47 
rect 141 47 142 48 
rect 141 58 142 59 
rect 141 59 142 60 
rect 141 60 142 61 
rect 141 61 142 62 
rect 141 62 142 63 
rect 141 63 142 64 
rect 141 74 142 75 
rect 141 75 142 76 
rect 141 76 142 77 
rect 141 77 142 78 
rect 141 78 142 79 
rect 141 79 142 80 
rect 141 90 142 91 
rect 141 91 142 92 
rect 141 92 142 93 
rect 141 93 142 94 
rect 141 94 142 95 
rect 141 95 142 96 
rect 141 106 142 107 
rect 141 107 142 108 
rect 141 108 142 109 
rect 141 109 142 110 
rect 141 110 142 111 
rect 141 111 142 112 
rect 141 122 142 123 
rect 141 123 142 124 
rect 141 124 142 125 
rect 141 125 142 126 
rect 141 126 142 127 
rect 141 127 142 128 
rect 141 138 142 139 
rect 141 139 142 140 
rect 141 140 142 141 
rect 141 141 142 142 
rect 141 142 142 143 
rect 141 143 142 144 
rect 141 154 142 155 
rect 141 155 142 156 
rect 141 156 142 157 
rect 141 157 142 158 
rect 141 158 142 159 
rect 141 159 142 160 
rect 141 170 142 171 
rect 141 171 142 172 
rect 141 172 142 173 
rect 141 173 142 174 
rect 141 174 142 175 
rect 141 175 142 176 
rect 141 186 142 187 
rect 141 187 142 188 
rect 141 188 142 189 
rect 141 189 142 190 
rect 141 190 142 191 
rect 141 191 142 192 
rect 141 202 142 203 
rect 141 203 142 204 
rect 141 204 142 205 
rect 141 205 142 206 
rect 141 206 142 207 
rect 141 207 142 208 
rect 141 218 142 219 
rect 141 219 142 220 
rect 141 220 142 221 
rect 141 221 142 222 
rect 141 222 142 223 
rect 141 223 142 224 
rect 141 234 142 235 
rect 141 235 142 236 
rect 141 236 142 237 
rect 141 237 142 238 
rect 141 238 142 239 
rect 141 239 142 240 
rect 141 250 142 251 
rect 141 251 142 252 
rect 141 252 142 253 
rect 141 253 142 254 
rect 141 254 142 255 
rect 141 255 142 256 
rect 141 266 142 267 
rect 141 267 142 268 
rect 141 268 142 269 
rect 141 269 142 270 
rect 141 270 142 271 
rect 141 271 142 272 
rect 141 282 142 283 
rect 141 283 142 284 
rect 141 284 142 285 
rect 141 285 142 286 
rect 141 286 142 287 
rect 141 287 142 288 
rect 141 298 142 299 
rect 141 299 142 300 
rect 141 300 142 301 
rect 141 301 142 302 
rect 141 302 142 303 
rect 141 303 142 304 
rect 142 10 143 11 
rect 142 11 143 12 
rect 142 12 143 13 
rect 142 13 143 14 
rect 142 14 143 15 
rect 142 15 143 16 
rect 142 26 143 27 
rect 142 27 143 28 
rect 142 28 143 29 
rect 142 29 143 30 
rect 142 30 143 31 
rect 142 31 143 32 
rect 142 42 143 43 
rect 142 43 143 44 
rect 142 44 143 45 
rect 142 45 143 46 
rect 142 46 143 47 
rect 142 47 143 48 
rect 142 58 143 59 
rect 142 59 143 60 
rect 142 60 143 61 
rect 142 61 143 62 
rect 142 62 143 63 
rect 142 63 143 64 
rect 142 74 143 75 
rect 142 75 143 76 
rect 142 76 143 77 
rect 142 77 143 78 
rect 142 78 143 79 
rect 142 79 143 80 
rect 142 90 143 91 
rect 142 91 143 92 
rect 142 92 143 93 
rect 142 93 143 94 
rect 142 94 143 95 
rect 142 95 143 96 
rect 142 106 143 107 
rect 142 107 143 108 
rect 142 108 143 109 
rect 142 109 143 110 
rect 142 110 143 111 
rect 142 111 143 112 
rect 142 122 143 123 
rect 142 123 143 124 
rect 142 124 143 125 
rect 142 125 143 126 
rect 142 126 143 127 
rect 142 127 143 128 
rect 142 138 143 139 
rect 142 139 143 140 
rect 142 140 143 141 
rect 142 141 143 142 
rect 142 142 143 143 
rect 142 143 143 144 
rect 142 154 143 155 
rect 142 155 143 156 
rect 142 156 143 157 
rect 142 157 143 158 
rect 142 158 143 159 
rect 142 159 143 160 
rect 142 170 143 171 
rect 142 171 143 172 
rect 142 172 143 173 
rect 142 173 143 174 
rect 142 174 143 175 
rect 142 175 143 176 
rect 142 186 143 187 
rect 142 187 143 188 
rect 142 188 143 189 
rect 142 189 143 190 
rect 142 190 143 191 
rect 142 191 143 192 
rect 142 202 143 203 
rect 142 203 143 204 
rect 142 204 143 205 
rect 142 205 143 206 
rect 142 206 143 207 
rect 142 207 143 208 
rect 142 218 143 219 
rect 142 219 143 220 
rect 142 220 143 221 
rect 142 221 143 222 
rect 142 222 143 223 
rect 142 223 143 224 
rect 142 234 143 235 
rect 142 235 143 236 
rect 142 236 143 237 
rect 142 237 143 238 
rect 142 238 143 239 
rect 142 239 143 240 
rect 142 250 143 251 
rect 142 251 143 252 
rect 142 252 143 253 
rect 142 253 143 254 
rect 142 254 143 255 
rect 142 255 143 256 
rect 142 266 143 267 
rect 142 267 143 268 
rect 142 268 143 269 
rect 142 269 143 270 
rect 142 270 143 271 
rect 142 271 143 272 
rect 142 282 143 283 
rect 142 283 143 284 
rect 142 284 143 285 
rect 142 285 143 286 
rect 142 286 143 287 
rect 142 287 143 288 
rect 142 298 143 299 
rect 142 299 143 300 
rect 142 300 143 301 
rect 142 301 143 302 
rect 142 302 143 303 
rect 142 303 143 304 
rect 143 10 144 11 
rect 143 11 144 12 
rect 143 12 144 13 
rect 143 13 144 14 
rect 143 15 144 16 
rect 143 26 144 27 
rect 143 28 144 29 
rect 143 29 144 30 
rect 143 30 144 31 
rect 143 31 144 32 
rect 143 42 144 43 
rect 143 43 144 44 
rect 143 44 144 45 
rect 143 45 144 46 
rect 143 46 144 47 
rect 143 47 144 48 
rect 143 58 144 59 
rect 143 59 144 60 
rect 143 60 144 61 
rect 143 61 144 62 
rect 143 63 144 64 
rect 143 74 144 75 
rect 143 76 144 77 
rect 143 77 144 78 
rect 143 78 144 79 
rect 143 79 144 80 
rect 143 90 144 91 
rect 143 91 144 92 
rect 143 92 144 93 
rect 143 93 144 94 
rect 143 94 144 95 
rect 143 95 144 96 
rect 143 106 144 107 
rect 143 108 144 109 
rect 143 109 144 110 
rect 143 110 144 111 
rect 143 111 144 112 
rect 143 122 144 123 
rect 143 123 144 124 
rect 143 124 144 125 
rect 143 125 144 126 
rect 143 126 144 127 
rect 143 127 144 128 
rect 143 138 144 139 
rect 143 140 144 141 
rect 143 141 144 142 
rect 143 142 144 143 
rect 143 143 144 144 
rect 143 154 144 155 
rect 143 155 144 156 
rect 143 156 144 157 
rect 143 157 144 158 
rect 143 158 144 159 
rect 143 159 144 160 
rect 143 170 144 171 
rect 143 171 144 172 
rect 143 172 144 173 
rect 143 173 144 174 
rect 143 174 144 175 
rect 143 175 144 176 
rect 143 186 144 187 
rect 143 187 144 188 
rect 143 188 144 189 
rect 143 189 144 190 
rect 143 191 144 192 
rect 143 202 144 203 
rect 143 204 144 205 
rect 143 205 144 206 
rect 143 207 144 208 
rect 143 218 144 219 
rect 143 220 144 221 
rect 143 221 144 222 
rect 143 222 144 223 
rect 143 223 144 224 
rect 143 234 144 235 
rect 143 235 144 236 
rect 143 236 144 237 
rect 143 237 144 238 
rect 143 238 144 239 
rect 143 239 144 240 
rect 143 250 144 251 
rect 143 252 144 253 
rect 143 253 144 254 
rect 143 254 144 255 
rect 143 255 144 256 
rect 143 266 144 267 
rect 143 267 144 268 
rect 143 268 144 269 
rect 143 269 144 270 
rect 143 270 144 271 
rect 143 271 144 272 
rect 143 282 144 283 
rect 143 283 144 284 
rect 143 284 144 285 
rect 143 285 144 286 
rect 143 286 144 287 
rect 143 287 144 288 
rect 143 298 144 299 
rect 143 299 144 300 
rect 143 300 144 301 
rect 143 301 144 302 
rect 143 303 144 304 
rect 154 10 155 11 
rect 154 11 155 12 
rect 154 12 155 13 
rect 154 13 155 14 
rect 154 15 155 16 
rect 154 26 155 27 
rect 154 27 155 28 
rect 154 28 155 29 
rect 154 29 155 30 
rect 154 31 155 32 
rect 154 42 155 43 
rect 154 43 155 44 
rect 154 44 155 45 
rect 154 45 155 46 
rect 154 46 155 47 
rect 154 47 155 48 
rect 154 58 155 59 
rect 154 59 155 60 
rect 154 60 155 61 
rect 154 61 155 62 
rect 154 63 155 64 
rect 154 74 155 75 
rect 154 76 155 77 
rect 154 77 155 78 
rect 154 79 155 80 
rect 154 90 155 91 
rect 154 91 155 92 
rect 154 92 155 93 
rect 154 93 155 94 
rect 154 95 155 96 
rect 154 106 155 107 
rect 154 108 155 109 
rect 154 109 155 110 
rect 154 110 155 111 
rect 154 111 155 112 
rect 154 122 155 123 
rect 154 123 155 124 
rect 154 124 155 125 
rect 154 125 155 126 
rect 154 127 155 128 
rect 154 138 155 139 
rect 154 139 155 140 
rect 154 140 155 141 
rect 154 141 155 142 
rect 154 142 155 143 
rect 154 143 155 144 
rect 154 154 155 155 
rect 154 156 155 157 
rect 154 157 155 158 
rect 154 159 155 160 
rect 154 170 155 171 
rect 154 172 155 173 
rect 154 173 155 174 
rect 154 175 155 176 
rect 154 186 155 187 
rect 154 187 155 188 
rect 154 188 155 189 
rect 154 189 155 190 
rect 154 191 155 192 
rect 154 202 155 203 
rect 154 204 155 205 
rect 154 205 155 206 
rect 154 206 155 207 
rect 154 207 155 208 
rect 154 218 155 219 
rect 154 220 155 221 
rect 154 221 155 222 
rect 154 223 155 224 
rect 154 234 155 235 
rect 154 236 155 237 
rect 154 237 155 238 
rect 154 239 155 240 
rect 154 250 155 251 
rect 154 251 155 252 
rect 154 252 155 253 
rect 154 253 155 254 
rect 154 254 155 255 
rect 154 255 155 256 
rect 154 266 155 267 
rect 154 268 155 269 
rect 154 269 155 270 
rect 154 270 155 271 
rect 154 271 155 272 
rect 154 282 155 283 
rect 154 283 155 284 
rect 154 284 155 285 
rect 154 285 155 286 
rect 154 287 155 288 
rect 154 298 155 299 
rect 154 299 155 300 
rect 154 300 155 301 
rect 154 301 155 302 
rect 154 302 155 303 
rect 154 303 155 304 
rect 155 10 156 11 
rect 155 11 156 12 
rect 155 12 156 13 
rect 155 13 156 14 
rect 155 14 156 15 
rect 155 15 156 16 
rect 155 26 156 27 
rect 155 27 156 28 
rect 155 28 156 29 
rect 155 29 156 30 
rect 155 30 156 31 
rect 155 31 156 32 
rect 155 42 156 43 
rect 155 43 156 44 
rect 155 44 156 45 
rect 155 45 156 46 
rect 155 46 156 47 
rect 155 47 156 48 
rect 155 58 156 59 
rect 155 59 156 60 
rect 155 60 156 61 
rect 155 61 156 62 
rect 155 62 156 63 
rect 155 63 156 64 
rect 155 74 156 75 
rect 155 75 156 76 
rect 155 76 156 77 
rect 155 77 156 78 
rect 155 78 156 79 
rect 155 79 156 80 
rect 155 90 156 91 
rect 155 91 156 92 
rect 155 92 156 93 
rect 155 93 156 94 
rect 155 94 156 95 
rect 155 95 156 96 
rect 155 106 156 107 
rect 155 107 156 108 
rect 155 108 156 109 
rect 155 109 156 110 
rect 155 110 156 111 
rect 155 111 156 112 
rect 155 122 156 123 
rect 155 123 156 124 
rect 155 124 156 125 
rect 155 125 156 126 
rect 155 126 156 127 
rect 155 127 156 128 
rect 155 138 156 139 
rect 155 139 156 140 
rect 155 140 156 141 
rect 155 141 156 142 
rect 155 142 156 143 
rect 155 143 156 144 
rect 155 154 156 155 
rect 155 155 156 156 
rect 155 156 156 157 
rect 155 157 156 158 
rect 155 158 156 159 
rect 155 159 156 160 
rect 155 170 156 171 
rect 155 171 156 172 
rect 155 172 156 173 
rect 155 173 156 174 
rect 155 174 156 175 
rect 155 175 156 176 
rect 155 186 156 187 
rect 155 187 156 188 
rect 155 188 156 189 
rect 155 189 156 190 
rect 155 190 156 191 
rect 155 191 156 192 
rect 155 202 156 203 
rect 155 203 156 204 
rect 155 204 156 205 
rect 155 205 156 206 
rect 155 206 156 207 
rect 155 207 156 208 
rect 155 218 156 219 
rect 155 219 156 220 
rect 155 220 156 221 
rect 155 221 156 222 
rect 155 222 156 223 
rect 155 223 156 224 
rect 155 234 156 235 
rect 155 235 156 236 
rect 155 236 156 237 
rect 155 237 156 238 
rect 155 238 156 239 
rect 155 239 156 240 
rect 155 250 156 251 
rect 155 251 156 252 
rect 155 252 156 253 
rect 155 253 156 254 
rect 155 254 156 255 
rect 155 255 156 256 
rect 155 266 156 267 
rect 155 267 156 268 
rect 155 268 156 269 
rect 155 269 156 270 
rect 155 270 156 271 
rect 155 271 156 272 
rect 155 282 156 283 
rect 155 283 156 284 
rect 155 284 156 285 
rect 155 285 156 286 
rect 155 286 156 287 
rect 155 287 156 288 
rect 155 298 156 299 
rect 155 299 156 300 
rect 155 300 156 301 
rect 155 301 156 302 
rect 155 302 156 303 
rect 155 303 156 304 
rect 156 10 157 11 
rect 156 11 157 12 
rect 156 12 157 13 
rect 156 13 157 14 
rect 156 14 157 15 
rect 156 15 157 16 
rect 156 26 157 27 
rect 156 27 157 28 
rect 156 28 157 29 
rect 156 29 157 30 
rect 156 30 157 31 
rect 156 31 157 32 
rect 156 42 157 43 
rect 156 43 157 44 
rect 156 44 157 45 
rect 156 45 157 46 
rect 156 46 157 47 
rect 156 47 157 48 
rect 156 58 157 59 
rect 156 59 157 60 
rect 156 60 157 61 
rect 156 61 157 62 
rect 156 62 157 63 
rect 156 63 157 64 
rect 156 74 157 75 
rect 156 75 157 76 
rect 156 76 157 77 
rect 156 77 157 78 
rect 156 78 157 79 
rect 156 79 157 80 
rect 156 90 157 91 
rect 156 91 157 92 
rect 156 92 157 93 
rect 156 93 157 94 
rect 156 94 157 95 
rect 156 95 157 96 
rect 156 106 157 107 
rect 156 107 157 108 
rect 156 108 157 109 
rect 156 109 157 110 
rect 156 110 157 111 
rect 156 111 157 112 
rect 156 122 157 123 
rect 156 123 157 124 
rect 156 124 157 125 
rect 156 125 157 126 
rect 156 126 157 127 
rect 156 127 157 128 
rect 156 138 157 139 
rect 156 139 157 140 
rect 156 140 157 141 
rect 156 141 157 142 
rect 156 142 157 143 
rect 156 143 157 144 
rect 156 154 157 155 
rect 156 155 157 156 
rect 156 156 157 157 
rect 156 157 157 158 
rect 156 158 157 159 
rect 156 159 157 160 
rect 156 170 157 171 
rect 156 171 157 172 
rect 156 172 157 173 
rect 156 173 157 174 
rect 156 174 157 175 
rect 156 175 157 176 
rect 156 186 157 187 
rect 156 187 157 188 
rect 156 188 157 189 
rect 156 189 157 190 
rect 156 190 157 191 
rect 156 191 157 192 
rect 156 202 157 203 
rect 156 203 157 204 
rect 156 204 157 205 
rect 156 205 157 206 
rect 156 206 157 207 
rect 156 207 157 208 
rect 156 218 157 219 
rect 156 219 157 220 
rect 156 220 157 221 
rect 156 221 157 222 
rect 156 222 157 223 
rect 156 223 157 224 
rect 156 234 157 235 
rect 156 235 157 236 
rect 156 236 157 237 
rect 156 237 157 238 
rect 156 238 157 239 
rect 156 239 157 240 
rect 156 250 157 251 
rect 156 251 157 252 
rect 156 252 157 253 
rect 156 253 157 254 
rect 156 254 157 255 
rect 156 255 157 256 
rect 156 266 157 267 
rect 156 267 157 268 
rect 156 268 157 269 
rect 156 269 157 270 
rect 156 270 157 271 
rect 156 271 157 272 
rect 156 282 157 283 
rect 156 283 157 284 
rect 156 284 157 285 
rect 156 285 157 286 
rect 156 286 157 287 
rect 156 287 157 288 
rect 156 298 157 299 
rect 156 299 157 300 
rect 156 300 157 301 
rect 156 301 157 302 
rect 156 302 157 303 
rect 156 303 157 304 
rect 157 10 158 11 
rect 157 11 158 12 
rect 157 12 158 13 
rect 157 13 158 14 
rect 157 14 158 15 
rect 157 15 158 16 
rect 157 26 158 27 
rect 157 27 158 28 
rect 157 28 158 29 
rect 157 29 158 30 
rect 157 30 158 31 
rect 157 31 158 32 
rect 157 42 158 43 
rect 157 43 158 44 
rect 157 44 158 45 
rect 157 45 158 46 
rect 157 46 158 47 
rect 157 47 158 48 
rect 157 58 158 59 
rect 157 59 158 60 
rect 157 60 158 61 
rect 157 61 158 62 
rect 157 62 158 63 
rect 157 63 158 64 
rect 157 74 158 75 
rect 157 75 158 76 
rect 157 76 158 77 
rect 157 77 158 78 
rect 157 78 158 79 
rect 157 79 158 80 
rect 157 90 158 91 
rect 157 91 158 92 
rect 157 92 158 93 
rect 157 93 158 94 
rect 157 94 158 95 
rect 157 95 158 96 
rect 157 106 158 107 
rect 157 107 158 108 
rect 157 108 158 109 
rect 157 109 158 110 
rect 157 110 158 111 
rect 157 111 158 112 
rect 157 122 158 123 
rect 157 123 158 124 
rect 157 124 158 125 
rect 157 125 158 126 
rect 157 126 158 127 
rect 157 127 158 128 
rect 157 138 158 139 
rect 157 139 158 140 
rect 157 140 158 141 
rect 157 141 158 142 
rect 157 142 158 143 
rect 157 143 158 144 
rect 157 154 158 155 
rect 157 155 158 156 
rect 157 156 158 157 
rect 157 157 158 158 
rect 157 158 158 159 
rect 157 159 158 160 
rect 157 170 158 171 
rect 157 171 158 172 
rect 157 172 158 173 
rect 157 173 158 174 
rect 157 174 158 175 
rect 157 175 158 176 
rect 157 186 158 187 
rect 157 187 158 188 
rect 157 188 158 189 
rect 157 189 158 190 
rect 157 190 158 191 
rect 157 191 158 192 
rect 157 202 158 203 
rect 157 203 158 204 
rect 157 204 158 205 
rect 157 205 158 206 
rect 157 206 158 207 
rect 157 207 158 208 
rect 157 218 158 219 
rect 157 219 158 220 
rect 157 220 158 221 
rect 157 221 158 222 
rect 157 222 158 223 
rect 157 223 158 224 
rect 157 234 158 235 
rect 157 235 158 236 
rect 157 236 158 237 
rect 157 237 158 238 
rect 157 238 158 239 
rect 157 239 158 240 
rect 157 250 158 251 
rect 157 251 158 252 
rect 157 252 158 253 
rect 157 253 158 254 
rect 157 254 158 255 
rect 157 255 158 256 
rect 157 266 158 267 
rect 157 267 158 268 
rect 157 268 158 269 
rect 157 269 158 270 
rect 157 270 158 271 
rect 157 271 158 272 
rect 157 282 158 283 
rect 157 283 158 284 
rect 157 284 158 285 
rect 157 285 158 286 
rect 157 286 158 287 
rect 157 287 158 288 
rect 157 298 158 299 
rect 157 299 158 300 
rect 157 300 158 301 
rect 157 301 158 302 
rect 157 302 158 303 
rect 157 303 158 304 
rect 158 10 159 11 
rect 158 11 159 12 
rect 158 12 159 13 
rect 158 13 159 14 
rect 158 14 159 15 
rect 158 15 159 16 
rect 158 26 159 27 
rect 158 27 159 28 
rect 158 28 159 29 
rect 158 29 159 30 
rect 158 30 159 31 
rect 158 31 159 32 
rect 158 42 159 43 
rect 158 43 159 44 
rect 158 44 159 45 
rect 158 45 159 46 
rect 158 46 159 47 
rect 158 47 159 48 
rect 158 58 159 59 
rect 158 59 159 60 
rect 158 60 159 61 
rect 158 61 159 62 
rect 158 62 159 63 
rect 158 63 159 64 
rect 158 74 159 75 
rect 158 75 159 76 
rect 158 76 159 77 
rect 158 77 159 78 
rect 158 78 159 79 
rect 158 79 159 80 
rect 158 90 159 91 
rect 158 91 159 92 
rect 158 92 159 93 
rect 158 93 159 94 
rect 158 94 159 95 
rect 158 95 159 96 
rect 158 106 159 107 
rect 158 107 159 108 
rect 158 108 159 109 
rect 158 109 159 110 
rect 158 110 159 111 
rect 158 111 159 112 
rect 158 122 159 123 
rect 158 123 159 124 
rect 158 124 159 125 
rect 158 125 159 126 
rect 158 126 159 127 
rect 158 127 159 128 
rect 158 138 159 139 
rect 158 139 159 140 
rect 158 140 159 141 
rect 158 141 159 142 
rect 158 142 159 143 
rect 158 143 159 144 
rect 158 154 159 155 
rect 158 155 159 156 
rect 158 156 159 157 
rect 158 157 159 158 
rect 158 158 159 159 
rect 158 159 159 160 
rect 158 170 159 171 
rect 158 171 159 172 
rect 158 172 159 173 
rect 158 173 159 174 
rect 158 174 159 175 
rect 158 175 159 176 
rect 158 186 159 187 
rect 158 187 159 188 
rect 158 188 159 189 
rect 158 189 159 190 
rect 158 190 159 191 
rect 158 191 159 192 
rect 158 202 159 203 
rect 158 203 159 204 
rect 158 204 159 205 
rect 158 205 159 206 
rect 158 206 159 207 
rect 158 207 159 208 
rect 158 218 159 219 
rect 158 219 159 220 
rect 158 220 159 221 
rect 158 221 159 222 
rect 158 222 159 223 
rect 158 223 159 224 
rect 158 234 159 235 
rect 158 235 159 236 
rect 158 236 159 237 
rect 158 237 159 238 
rect 158 238 159 239 
rect 158 239 159 240 
rect 158 250 159 251 
rect 158 251 159 252 
rect 158 252 159 253 
rect 158 253 159 254 
rect 158 254 159 255 
rect 158 255 159 256 
rect 158 266 159 267 
rect 158 267 159 268 
rect 158 268 159 269 
rect 158 269 159 270 
rect 158 270 159 271 
rect 158 271 159 272 
rect 158 282 159 283 
rect 158 283 159 284 
rect 158 284 159 285 
rect 158 285 159 286 
rect 158 286 159 287 
rect 158 287 159 288 
rect 158 298 159 299 
rect 158 299 159 300 
rect 158 300 159 301 
rect 158 301 159 302 
rect 158 302 159 303 
rect 158 303 159 304 
rect 159 10 160 11 
rect 159 12 160 13 
rect 159 13 160 14 
rect 159 14 160 15 
rect 159 15 160 16 
rect 159 26 160 27 
rect 159 27 160 28 
rect 159 28 160 29 
rect 159 29 160 30 
rect 159 30 160 31 
rect 159 31 160 32 
rect 159 42 160 43 
rect 159 43 160 44 
rect 159 44 160 45 
rect 159 45 160 46 
rect 159 47 160 48 
rect 159 58 160 59 
rect 159 59 160 60 
rect 159 60 160 61 
rect 159 61 160 62 
rect 159 62 160 63 
rect 159 63 160 64 
rect 159 74 160 75 
rect 159 76 160 77 
rect 159 77 160 78 
rect 159 78 160 79 
rect 159 79 160 80 
rect 159 90 160 91 
rect 159 91 160 92 
rect 159 92 160 93 
rect 159 93 160 94 
rect 159 94 160 95 
rect 159 95 160 96 
rect 159 106 160 107 
rect 159 108 160 109 
rect 159 109 160 110 
rect 159 110 160 111 
rect 159 111 160 112 
rect 159 122 160 123 
rect 159 124 160 125 
rect 159 125 160 126 
rect 159 127 160 128 
rect 159 138 160 139 
rect 159 140 160 141 
rect 159 141 160 142 
rect 159 142 160 143 
rect 159 143 160 144 
rect 159 154 160 155 
rect 159 155 160 156 
rect 159 156 160 157 
rect 159 157 160 158 
rect 159 159 160 160 
rect 159 170 160 171 
rect 159 171 160 172 
rect 159 172 160 173 
rect 159 173 160 174 
rect 159 175 160 176 
rect 159 186 160 187 
rect 159 188 160 189 
rect 159 189 160 190 
rect 159 191 160 192 
rect 159 202 160 203 
rect 159 204 160 205 
rect 159 205 160 206 
rect 159 206 160 207 
rect 159 207 160 208 
rect 159 218 160 219 
rect 159 220 160 221 
rect 159 221 160 222 
rect 159 222 160 223 
rect 159 223 160 224 
rect 159 234 160 235 
rect 159 235 160 236 
rect 159 236 160 237 
rect 159 237 160 238 
rect 159 239 160 240 
rect 159 250 160 251 
rect 159 252 160 253 
rect 159 253 160 254 
rect 159 255 160 256 
rect 159 266 160 267 
rect 159 267 160 268 
rect 159 268 160 269 
rect 159 269 160 270 
rect 159 271 160 272 
rect 159 282 160 283 
rect 159 283 160 284 
rect 159 284 160 285 
rect 159 285 160 286 
rect 159 287 160 288 
rect 159 298 160 299 
rect 159 299 160 300 
rect 159 300 160 301 
rect 159 301 160 302 
rect 159 302 160 303 
rect 159 303 160 304 
rect 170 10 171 11 
rect 170 12 171 13 
rect 170 13 171 14 
rect 170 14 171 15 
rect 170 15 171 16 
rect 170 26 171 27 
rect 170 27 171 28 
rect 170 28 171 29 
rect 170 29 171 30 
rect 170 31 171 32 
rect 170 42 171 43 
rect 170 44 171 45 
rect 170 45 171 46 
rect 170 46 171 47 
rect 170 47 171 48 
rect 170 58 171 59 
rect 170 60 171 61 
rect 170 61 171 62 
rect 170 62 171 63 
rect 170 63 171 64 
rect 170 74 171 75 
rect 170 76 171 77 
rect 170 77 171 78 
rect 170 79 171 80 
rect 170 90 171 91 
rect 170 92 171 93 
rect 170 93 171 94 
rect 170 94 171 95 
rect 170 95 171 96 
rect 170 106 171 107 
rect 170 108 171 109 
rect 170 109 171 110 
rect 170 110 171 111 
rect 170 111 171 112 
rect 170 122 171 123 
rect 170 124 171 125 
rect 170 125 171 126 
rect 170 127 171 128 
rect 170 138 171 139 
rect 170 140 171 141 
rect 170 141 171 142 
rect 170 143 171 144 
rect 170 154 171 155 
rect 170 156 171 157 
rect 170 157 171 158 
rect 170 159 171 160 
rect 170 170 171 171 
rect 170 171 171 172 
rect 170 172 171 173 
rect 170 173 171 174 
rect 170 175 171 176 
rect 170 186 171 187 
rect 170 188 171 189 
rect 170 189 171 190 
rect 170 190 171 191 
rect 170 191 171 192 
rect 170 202 171 203 
rect 170 203 171 204 
rect 170 204 171 205 
rect 170 205 171 206 
rect 170 206 171 207 
rect 170 207 171 208 
rect 170 218 171 219 
rect 170 219 171 220 
rect 170 220 171 221 
rect 170 221 171 222 
rect 170 223 171 224 
rect 170 234 171 235 
rect 170 236 171 237 
rect 170 237 171 238 
rect 170 239 171 240 
rect 170 250 171 251 
rect 170 251 171 252 
rect 170 252 171 253 
rect 170 253 171 254 
rect 170 255 171 256 
rect 170 266 171 267 
rect 170 268 171 269 
rect 170 269 171 270 
rect 170 270 171 271 
rect 170 271 171 272 
rect 170 282 171 283 
rect 170 284 171 285 
rect 170 285 171 286 
rect 170 286 171 287 
rect 170 287 171 288 
rect 170 298 171 299 
rect 170 299 171 300 
rect 170 300 171 301 
rect 170 301 171 302 
rect 170 302 171 303 
rect 170 303 171 304 
rect 171 10 172 11 
rect 171 11 172 12 
rect 171 12 172 13 
rect 171 13 172 14 
rect 171 14 172 15 
rect 171 15 172 16 
rect 171 26 172 27 
rect 171 27 172 28 
rect 171 28 172 29 
rect 171 29 172 30 
rect 171 30 172 31 
rect 171 31 172 32 
rect 171 42 172 43 
rect 171 43 172 44 
rect 171 44 172 45 
rect 171 45 172 46 
rect 171 46 172 47 
rect 171 47 172 48 
rect 171 58 172 59 
rect 171 59 172 60 
rect 171 60 172 61 
rect 171 61 172 62 
rect 171 62 172 63 
rect 171 63 172 64 
rect 171 74 172 75 
rect 171 75 172 76 
rect 171 76 172 77 
rect 171 77 172 78 
rect 171 78 172 79 
rect 171 79 172 80 
rect 171 90 172 91 
rect 171 91 172 92 
rect 171 92 172 93 
rect 171 93 172 94 
rect 171 94 172 95 
rect 171 95 172 96 
rect 171 106 172 107 
rect 171 107 172 108 
rect 171 108 172 109 
rect 171 109 172 110 
rect 171 110 172 111 
rect 171 111 172 112 
rect 171 122 172 123 
rect 171 123 172 124 
rect 171 124 172 125 
rect 171 125 172 126 
rect 171 126 172 127 
rect 171 127 172 128 
rect 171 138 172 139 
rect 171 139 172 140 
rect 171 140 172 141 
rect 171 141 172 142 
rect 171 142 172 143 
rect 171 143 172 144 
rect 171 154 172 155 
rect 171 155 172 156 
rect 171 156 172 157 
rect 171 157 172 158 
rect 171 158 172 159 
rect 171 159 172 160 
rect 171 170 172 171 
rect 171 171 172 172 
rect 171 172 172 173 
rect 171 173 172 174 
rect 171 174 172 175 
rect 171 175 172 176 
rect 171 186 172 187 
rect 171 187 172 188 
rect 171 188 172 189 
rect 171 189 172 190 
rect 171 190 172 191 
rect 171 191 172 192 
rect 171 202 172 203 
rect 171 203 172 204 
rect 171 204 172 205 
rect 171 205 172 206 
rect 171 206 172 207 
rect 171 207 172 208 
rect 171 218 172 219 
rect 171 219 172 220 
rect 171 220 172 221 
rect 171 221 172 222 
rect 171 222 172 223 
rect 171 223 172 224 
rect 171 234 172 235 
rect 171 235 172 236 
rect 171 236 172 237 
rect 171 237 172 238 
rect 171 238 172 239 
rect 171 239 172 240 
rect 171 250 172 251 
rect 171 251 172 252 
rect 171 252 172 253 
rect 171 253 172 254 
rect 171 254 172 255 
rect 171 255 172 256 
rect 171 266 172 267 
rect 171 267 172 268 
rect 171 268 172 269 
rect 171 269 172 270 
rect 171 270 172 271 
rect 171 271 172 272 
rect 171 282 172 283 
rect 171 283 172 284 
rect 171 284 172 285 
rect 171 285 172 286 
rect 171 286 172 287 
rect 171 287 172 288 
rect 171 298 172 299 
rect 171 299 172 300 
rect 171 300 172 301 
rect 171 301 172 302 
rect 171 302 172 303 
rect 171 303 172 304 
rect 172 10 173 11 
rect 172 11 173 12 
rect 172 12 173 13 
rect 172 13 173 14 
rect 172 14 173 15 
rect 172 15 173 16 
rect 172 26 173 27 
rect 172 27 173 28 
rect 172 28 173 29 
rect 172 29 173 30 
rect 172 30 173 31 
rect 172 31 173 32 
rect 172 42 173 43 
rect 172 43 173 44 
rect 172 44 173 45 
rect 172 45 173 46 
rect 172 46 173 47 
rect 172 47 173 48 
rect 172 58 173 59 
rect 172 59 173 60 
rect 172 60 173 61 
rect 172 61 173 62 
rect 172 62 173 63 
rect 172 63 173 64 
rect 172 74 173 75 
rect 172 75 173 76 
rect 172 76 173 77 
rect 172 77 173 78 
rect 172 78 173 79 
rect 172 79 173 80 
rect 172 90 173 91 
rect 172 91 173 92 
rect 172 92 173 93 
rect 172 93 173 94 
rect 172 94 173 95 
rect 172 95 173 96 
rect 172 106 173 107 
rect 172 107 173 108 
rect 172 108 173 109 
rect 172 109 173 110 
rect 172 110 173 111 
rect 172 111 173 112 
rect 172 122 173 123 
rect 172 123 173 124 
rect 172 124 173 125 
rect 172 125 173 126 
rect 172 126 173 127 
rect 172 127 173 128 
rect 172 138 173 139 
rect 172 139 173 140 
rect 172 140 173 141 
rect 172 141 173 142 
rect 172 142 173 143 
rect 172 143 173 144 
rect 172 154 173 155 
rect 172 155 173 156 
rect 172 156 173 157 
rect 172 157 173 158 
rect 172 158 173 159 
rect 172 159 173 160 
rect 172 170 173 171 
rect 172 171 173 172 
rect 172 172 173 173 
rect 172 173 173 174 
rect 172 174 173 175 
rect 172 175 173 176 
rect 172 186 173 187 
rect 172 187 173 188 
rect 172 188 173 189 
rect 172 189 173 190 
rect 172 190 173 191 
rect 172 191 173 192 
rect 172 202 173 203 
rect 172 203 173 204 
rect 172 204 173 205 
rect 172 205 173 206 
rect 172 206 173 207 
rect 172 207 173 208 
rect 172 218 173 219 
rect 172 219 173 220 
rect 172 220 173 221 
rect 172 221 173 222 
rect 172 222 173 223 
rect 172 223 173 224 
rect 172 234 173 235 
rect 172 235 173 236 
rect 172 236 173 237 
rect 172 237 173 238 
rect 172 238 173 239 
rect 172 239 173 240 
rect 172 250 173 251 
rect 172 251 173 252 
rect 172 252 173 253 
rect 172 253 173 254 
rect 172 254 173 255 
rect 172 255 173 256 
rect 172 266 173 267 
rect 172 267 173 268 
rect 172 268 173 269 
rect 172 269 173 270 
rect 172 270 173 271 
rect 172 271 173 272 
rect 172 282 173 283 
rect 172 283 173 284 
rect 172 284 173 285 
rect 172 285 173 286 
rect 172 286 173 287 
rect 172 287 173 288 
rect 172 298 173 299 
rect 172 299 173 300 
rect 172 300 173 301 
rect 172 301 173 302 
rect 172 302 173 303 
rect 172 303 173 304 
rect 173 10 174 11 
rect 173 11 174 12 
rect 173 12 174 13 
rect 173 13 174 14 
rect 173 14 174 15 
rect 173 15 174 16 
rect 173 26 174 27 
rect 173 27 174 28 
rect 173 28 174 29 
rect 173 29 174 30 
rect 173 30 174 31 
rect 173 31 174 32 
rect 173 42 174 43 
rect 173 43 174 44 
rect 173 44 174 45 
rect 173 45 174 46 
rect 173 46 174 47 
rect 173 47 174 48 
rect 173 58 174 59 
rect 173 59 174 60 
rect 173 60 174 61 
rect 173 61 174 62 
rect 173 62 174 63 
rect 173 63 174 64 
rect 173 74 174 75 
rect 173 75 174 76 
rect 173 76 174 77 
rect 173 77 174 78 
rect 173 78 174 79 
rect 173 79 174 80 
rect 173 90 174 91 
rect 173 91 174 92 
rect 173 92 174 93 
rect 173 93 174 94 
rect 173 94 174 95 
rect 173 95 174 96 
rect 173 106 174 107 
rect 173 107 174 108 
rect 173 108 174 109 
rect 173 109 174 110 
rect 173 110 174 111 
rect 173 111 174 112 
rect 173 122 174 123 
rect 173 123 174 124 
rect 173 124 174 125 
rect 173 125 174 126 
rect 173 126 174 127 
rect 173 127 174 128 
rect 173 138 174 139 
rect 173 139 174 140 
rect 173 140 174 141 
rect 173 141 174 142 
rect 173 142 174 143 
rect 173 143 174 144 
rect 173 154 174 155 
rect 173 155 174 156 
rect 173 156 174 157 
rect 173 157 174 158 
rect 173 158 174 159 
rect 173 159 174 160 
rect 173 170 174 171 
rect 173 171 174 172 
rect 173 172 174 173 
rect 173 173 174 174 
rect 173 174 174 175 
rect 173 175 174 176 
rect 173 186 174 187 
rect 173 187 174 188 
rect 173 188 174 189 
rect 173 189 174 190 
rect 173 190 174 191 
rect 173 191 174 192 
rect 173 202 174 203 
rect 173 203 174 204 
rect 173 204 174 205 
rect 173 205 174 206 
rect 173 206 174 207 
rect 173 207 174 208 
rect 173 218 174 219 
rect 173 219 174 220 
rect 173 220 174 221 
rect 173 221 174 222 
rect 173 222 174 223 
rect 173 223 174 224 
rect 173 234 174 235 
rect 173 235 174 236 
rect 173 236 174 237 
rect 173 237 174 238 
rect 173 238 174 239 
rect 173 239 174 240 
rect 173 250 174 251 
rect 173 251 174 252 
rect 173 252 174 253 
rect 173 253 174 254 
rect 173 254 174 255 
rect 173 255 174 256 
rect 173 266 174 267 
rect 173 267 174 268 
rect 173 268 174 269 
rect 173 269 174 270 
rect 173 270 174 271 
rect 173 271 174 272 
rect 173 282 174 283 
rect 173 283 174 284 
rect 173 284 174 285 
rect 173 285 174 286 
rect 173 286 174 287 
rect 173 287 174 288 
rect 173 298 174 299 
rect 173 299 174 300 
rect 173 300 174 301 
rect 173 301 174 302 
rect 173 302 174 303 
rect 173 303 174 304 
rect 174 10 175 11 
rect 174 11 175 12 
rect 174 12 175 13 
rect 174 13 175 14 
rect 174 14 175 15 
rect 174 15 175 16 
rect 174 26 175 27 
rect 174 27 175 28 
rect 174 28 175 29 
rect 174 29 175 30 
rect 174 30 175 31 
rect 174 31 175 32 
rect 174 42 175 43 
rect 174 43 175 44 
rect 174 44 175 45 
rect 174 45 175 46 
rect 174 46 175 47 
rect 174 47 175 48 
rect 174 58 175 59 
rect 174 59 175 60 
rect 174 60 175 61 
rect 174 61 175 62 
rect 174 62 175 63 
rect 174 63 175 64 
rect 174 74 175 75 
rect 174 75 175 76 
rect 174 76 175 77 
rect 174 77 175 78 
rect 174 78 175 79 
rect 174 79 175 80 
rect 174 90 175 91 
rect 174 91 175 92 
rect 174 92 175 93 
rect 174 93 175 94 
rect 174 94 175 95 
rect 174 95 175 96 
rect 174 106 175 107 
rect 174 107 175 108 
rect 174 108 175 109 
rect 174 109 175 110 
rect 174 110 175 111 
rect 174 111 175 112 
rect 174 122 175 123 
rect 174 123 175 124 
rect 174 124 175 125 
rect 174 125 175 126 
rect 174 126 175 127 
rect 174 127 175 128 
rect 174 138 175 139 
rect 174 139 175 140 
rect 174 140 175 141 
rect 174 141 175 142 
rect 174 142 175 143 
rect 174 143 175 144 
rect 174 154 175 155 
rect 174 155 175 156 
rect 174 156 175 157 
rect 174 157 175 158 
rect 174 158 175 159 
rect 174 159 175 160 
rect 174 170 175 171 
rect 174 171 175 172 
rect 174 172 175 173 
rect 174 173 175 174 
rect 174 174 175 175 
rect 174 175 175 176 
rect 174 186 175 187 
rect 174 187 175 188 
rect 174 188 175 189 
rect 174 189 175 190 
rect 174 190 175 191 
rect 174 191 175 192 
rect 174 202 175 203 
rect 174 203 175 204 
rect 174 204 175 205 
rect 174 205 175 206 
rect 174 206 175 207 
rect 174 207 175 208 
rect 174 218 175 219 
rect 174 219 175 220 
rect 174 220 175 221 
rect 174 221 175 222 
rect 174 222 175 223 
rect 174 223 175 224 
rect 174 234 175 235 
rect 174 235 175 236 
rect 174 236 175 237 
rect 174 237 175 238 
rect 174 238 175 239 
rect 174 239 175 240 
rect 174 250 175 251 
rect 174 251 175 252 
rect 174 252 175 253 
rect 174 253 175 254 
rect 174 254 175 255 
rect 174 255 175 256 
rect 174 266 175 267 
rect 174 267 175 268 
rect 174 268 175 269 
rect 174 269 175 270 
rect 174 270 175 271 
rect 174 271 175 272 
rect 174 282 175 283 
rect 174 283 175 284 
rect 174 284 175 285 
rect 174 285 175 286 
rect 174 286 175 287 
rect 174 287 175 288 
rect 174 298 175 299 
rect 174 299 175 300 
rect 174 300 175 301 
rect 174 301 175 302 
rect 174 302 175 303 
rect 174 303 175 304 
rect 175 10 176 11 
rect 175 12 176 13 
rect 175 13 176 14 
rect 175 14 176 15 
rect 175 15 176 16 
rect 175 26 176 27 
rect 175 28 176 29 
rect 175 29 176 30 
rect 175 31 176 32 
rect 175 42 176 43 
rect 175 43 176 44 
rect 175 44 176 45 
rect 175 45 176 46 
rect 175 47 176 48 
rect 175 58 176 59 
rect 175 60 176 61 
rect 175 61 176 62 
rect 175 63 176 64 
rect 175 74 176 75 
rect 175 76 176 77 
rect 175 77 176 78 
rect 175 78 176 79 
rect 175 79 176 80 
rect 175 90 176 91 
rect 175 92 176 93 
rect 175 93 176 94 
rect 175 94 176 95 
rect 175 95 176 96 
rect 175 106 176 107 
rect 175 108 176 109 
rect 175 109 176 110 
rect 175 111 176 112 
rect 175 122 176 123 
rect 175 123 176 124 
rect 175 124 176 125 
rect 175 125 176 126 
rect 175 127 176 128 
rect 175 138 176 139 
rect 175 139 176 140 
rect 175 140 176 141 
rect 175 141 176 142 
rect 175 143 176 144 
rect 175 154 176 155 
rect 175 156 176 157 
rect 175 157 176 158 
rect 175 159 176 160 
rect 175 170 176 171 
rect 175 172 176 173 
rect 175 173 176 174 
rect 175 175 176 176 
rect 175 186 176 187 
rect 175 187 176 188 
rect 175 188 176 189 
rect 175 189 176 190 
rect 175 191 176 192 
rect 175 202 176 203 
rect 175 203 176 204 
rect 175 204 176 205 
rect 175 205 176 206 
rect 175 206 176 207 
rect 175 207 176 208 
rect 175 218 176 219 
rect 175 219 176 220 
rect 175 220 176 221 
rect 175 221 176 222 
rect 175 223 176 224 
rect 175 234 176 235 
rect 175 235 176 236 
rect 175 236 176 237 
rect 175 237 176 238 
rect 175 239 176 240 
rect 175 250 176 251 
rect 175 251 176 252 
rect 175 252 176 253 
rect 175 253 176 254 
rect 175 254 176 255 
rect 175 255 176 256 
rect 175 266 176 267 
rect 175 267 176 268 
rect 175 268 176 269 
rect 175 269 176 270 
rect 175 271 176 272 
rect 175 282 176 283 
rect 175 283 176 284 
rect 175 284 176 285 
rect 175 285 176 286 
rect 175 287 176 288 
rect 175 298 176 299 
rect 175 300 176 301 
rect 175 301 176 302 
rect 175 302 176 303 
rect 175 303 176 304 
rect 186 10 187 11 
rect 186 12 187 13 
rect 186 13 187 14 
rect 186 15 187 16 
rect 186 26 187 27 
rect 186 28 187 29 
rect 186 29 187 30 
rect 186 31 187 32 
rect 186 42 187 43 
rect 186 43 187 44 
rect 186 44 187 45 
rect 186 45 187 46 
rect 186 47 187 48 
rect 186 58 187 59 
rect 186 59 187 60 
rect 186 60 187 61 
rect 186 61 187 62 
rect 186 63 187 64 
rect 186 74 187 75 
rect 186 76 187 77 
rect 186 77 187 78 
rect 186 79 187 80 
rect 186 90 187 91 
rect 186 92 187 93 
rect 186 93 187 94 
rect 186 94 187 95 
rect 186 95 187 96 
rect 186 106 187 107 
rect 186 108 187 109 
rect 186 109 187 110 
rect 186 111 187 112 
rect 186 122 187 123 
rect 186 124 187 125 
rect 186 125 187 126 
rect 186 126 187 127 
rect 186 127 187 128 
rect 186 138 187 139 
rect 186 139 187 140 
rect 186 140 187 141 
rect 186 141 187 142 
rect 186 143 187 144 
rect 186 154 187 155 
rect 186 156 187 157 
rect 186 157 187 158 
rect 186 159 187 160 
rect 186 170 187 171 
rect 186 171 187 172 
rect 186 172 187 173 
rect 186 173 187 174 
rect 186 174 187 175 
rect 186 175 187 176 
rect 186 186 187 187 
rect 186 187 187 188 
rect 186 188 187 189 
rect 186 189 187 190 
rect 186 190 187 191 
rect 186 191 187 192 
rect 186 202 187 203 
rect 186 204 187 205 
rect 186 205 187 206 
rect 186 206 187 207 
rect 186 207 187 208 
rect 186 218 187 219 
rect 186 219 187 220 
rect 186 220 187 221 
rect 186 221 187 222 
rect 186 223 187 224 
rect 186 234 187 235 
rect 186 235 187 236 
rect 186 236 187 237 
rect 186 237 187 238 
rect 186 238 187 239 
rect 186 239 187 240 
rect 186 250 187 251 
rect 186 252 187 253 
rect 186 253 187 254 
rect 186 254 187 255 
rect 186 255 187 256 
rect 186 266 187 267 
rect 186 268 187 269 
rect 186 269 187 270 
rect 186 270 187 271 
rect 186 271 187 272 
rect 186 282 187 283 
rect 186 283 187 284 
rect 186 284 187 285 
rect 186 285 187 286 
rect 186 287 187 288 
rect 186 298 187 299 
rect 186 300 187 301 
rect 186 301 187 302 
rect 186 302 187 303 
rect 186 303 187 304 
rect 187 10 188 11 
rect 187 11 188 12 
rect 187 12 188 13 
rect 187 13 188 14 
rect 187 14 188 15 
rect 187 15 188 16 
rect 187 26 188 27 
rect 187 27 188 28 
rect 187 28 188 29 
rect 187 29 188 30 
rect 187 30 188 31 
rect 187 31 188 32 
rect 187 42 188 43 
rect 187 43 188 44 
rect 187 44 188 45 
rect 187 45 188 46 
rect 187 46 188 47 
rect 187 47 188 48 
rect 187 58 188 59 
rect 187 59 188 60 
rect 187 60 188 61 
rect 187 61 188 62 
rect 187 62 188 63 
rect 187 63 188 64 
rect 187 74 188 75 
rect 187 75 188 76 
rect 187 76 188 77 
rect 187 77 188 78 
rect 187 78 188 79 
rect 187 79 188 80 
rect 187 90 188 91 
rect 187 91 188 92 
rect 187 92 188 93 
rect 187 93 188 94 
rect 187 94 188 95 
rect 187 95 188 96 
rect 187 106 188 107 
rect 187 107 188 108 
rect 187 108 188 109 
rect 187 109 188 110 
rect 187 110 188 111 
rect 187 111 188 112 
rect 187 122 188 123 
rect 187 123 188 124 
rect 187 124 188 125 
rect 187 125 188 126 
rect 187 126 188 127 
rect 187 127 188 128 
rect 187 138 188 139 
rect 187 139 188 140 
rect 187 140 188 141 
rect 187 141 188 142 
rect 187 142 188 143 
rect 187 143 188 144 
rect 187 154 188 155 
rect 187 155 188 156 
rect 187 156 188 157 
rect 187 157 188 158 
rect 187 158 188 159 
rect 187 159 188 160 
rect 187 170 188 171 
rect 187 171 188 172 
rect 187 172 188 173 
rect 187 173 188 174 
rect 187 174 188 175 
rect 187 175 188 176 
rect 187 186 188 187 
rect 187 187 188 188 
rect 187 188 188 189 
rect 187 189 188 190 
rect 187 190 188 191 
rect 187 191 188 192 
rect 187 202 188 203 
rect 187 203 188 204 
rect 187 204 188 205 
rect 187 205 188 206 
rect 187 206 188 207 
rect 187 207 188 208 
rect 187 218 188 219 
rect 187 219 188 220 
rect 187 220 188 221 
rect 187 221 188 222 
rect 187 222 188 223 
rect 187 223 188 224 
rect 187 234 188 235 
rect 187 235 188 236 
rect 187 236 188 237 
rect 187 237 188 238 
rect 187 238 188 239 
rect 187 239 188 240 
rect 187 250 188 251 
rect 187 251 188 252 
rect 187 252 188 253 
rect 187 253 188 254 
rect 187 254 188 255 
rect 187 255 188 256 
rect 187 266 188 267 
rect 187 267 188 268 
rect 187 268 188 269 
rect 187 269 188 270 
rect 187 270 188 271 
rect 187 271 188 272 
rect 187 282 188 283 
rect 187 283 188 284 
rect 187 284 188 285 
rect 187 285 188 286 
rect 187 286 188 287 
rect 187 287 188 288 
rect 187 298 188 299 
rect 187 299 188 300 
rect 187 300 188 301 
rect 187 301 188 302 
rect 187 302 188 303 
rect 187 303 188 304 
rect 188 10 189 11 
rect 188 11 189 12 
rect 188 12 189 13 
rect 188 13 189 14 
rect 188 14 189 15 
rect 188 15 189 16 
rect 188 26 189 27 
rect 188 27 189 28 
rect 188 28 189 29 
rect 188 29 189 30 
rect 188 30 189 31 
rect 188 31 189 32 
rect 188 42 189 43 
rect 188 43 189 44 
rect 188 44 189 45 
rect 188 45 189 46 
rect 188 46 189 47 
rect 188 47 189 48 
rect 188 58 189 59 
rect 188 59 189 60 
rect 188 60 189 61 
rect 188 61 189 62 
rect 188 62 189 63 
rect 188 63 189 64 
rect 188 74 189 75 
rect 188 75 189 76 
rect 188 76 189 77 
rect 188 77 189 78 
rect 188 78 189 79 
rect 188 79 189 80 
rect 188 90 189 91 
rect 188 91 189 92 
rect 188 92 189 93 
rect 188 93 189 94 
rect 188 94 189 95 
rect 188 95 189 96 
rect 188 106 189 107 
rect 188 107 189 108 
rect 188 108 189 109 
rect 188 109 189 110 
rect 188 110 189 111 
rect 188 111 189 112 
rect 188 122 189 123 
rect 188 123 189 124 
rect 188 124 189 125 
rect 188 125 189 126 
rect 188 126 189 127 
rect 188 127 189 128 
rect 188 138 189 139 
rect 188 139 189 140 
rect 188 140 189 141 
rect 188 141 189 142 
rect 188 142 189 143 
rect 188 143 189 144 
rect 188 154 189 155 
rect 188 155 189 156 
rect 188 156 189 157 
rect 188 157 189 158 
rect 188 158 189 159 
rect 188 159 189 160 
rect 188 170 189 171 
rect 188 171 189 172 
rect 188 172 189 173 
rect 188 173 189 174 
rect 188 174 189 175 
rect 188 175 189 176 
rect 188 186 189 187 
rect 188 187 189 188 
rect 188 188 189 189 
rect 188 189 189 190 
rect 188 190 189 191 
rect 188 191 189 192 
rect 188 202 189 203 
rect 188 203 189 204 
rect 188 204 189 205 
rect 188 205 189 206 
rect 188 206 189 207 
rect 188 207 189 208 
rect 188 218 189 219 
rect 188 219 189 220 
rect 188 220 189 221 
rect 188 221 189 222 
rect 188 222 189 223 
rect 188 223 189 224 
rect 188 234 189 235 
rect 188 235 189 236 
rect 188 236 189 237 
rect 188 237 189 238 
rect 188 238 189 239 
rect 188 239 189 240 
rect 188 250 189 251 
rect 188 251 189 252 
rect 188 252 189 253 
rect 188 253 189 254 
rect 188 254 189 255 
rect 188 255 189 256 
rect 188 266 189 267 
rect 188 267 189 268 
rect 188 268 189 269 
rect 188 269 189 270 
rect 188 270 189 271 
rect 188 271 189 272 
rect 188 282 189 283 
rect 188 283 189 284 
rect 188 284 189 285 
rect 188 285 189 286 
rect 188 286 189 287 
rect 188 287 189 288 
rect 188 298 189 299 
rect 188 299 189 300 
rect 188 300 189 301 
rect 188 301 189 302 
rect 188 302 189 303 
rect 188 303 189 304 
rect 189 10 190 11 
rect 189 11 190 12 
rect 189 12 190 13 
rect 189 13 190 14 
rect 189 14 190 15 
rect 189 15 190 16 
rect 189 26 190 27 
rect 189 27 190 28 
rect 189 28 190 29 
rect 189 29 190 30 
rect 189 30 190 31 
rect 189 31 190 32 
rect 189 42 190 43 
rect 189 43 190 44 
rect 189 44 190 45 
rect 189 45 190 46 
rect 189 46 190 47 
rect 189 47 190 48 
rect 189 58 190 59 
rect 189 59 190 60 
rect 189 60 190 61 
rect 189 61 190 62 
rect 189 62 190 63 
rect 189 63 190 64 
rect 189 74 190 75 
rect 189 75 190 76 
rect 189 76 190 77 
rect 189 77 190 78 
rect 189 78 190 79 
rect 189 79 190 80 
rect 189 90 190 91 
rect 189 91 190 92 
rect 189 92 190 93 
rect 189 93 190 94 
rect 189 94 190 95 
rect 189 95 190 96 
rect 189 106 190 107 
rect 189 107 190 108 
rect 189 108 190 109 
rect 189 109 190 110 
rect 189 110 190 111 
rect 189 111 190 112 
rect 189 122 190 123 
rect 189 123 190 124 
rect 189 124 190 125 
rect 189 125 190 126 
rect 189 126 190 127 
rect 189 127 190 128 
rect 189 138 190 139 
rect 189 139 190 140 
rect 189 140 190 141 
rect 189 141 190 142 
rect 189 142 190 143 
rect 189 143 190 144 
rect 189 154 190 155 
rect 189 155 190 156 
rect 189 156 190 157 
rect 189 157 190 158 
rect 189 158 190 159 
rect 189 159 190 160 
rect 189 170 190 171 
rect 189 171 190 172 
rect 189 172 190 173 
rect 189 173 190 174 
rect 189 174 190 175 
rect 189 175 190 176 
rect 189 186 190 187 
rect 189 187 190 188 
rect 189 188 190 189 
rect 189 189 190 190 
rect 189 190 190 191 
rect 189 191 190 192 
rect 189 202 190 203 
rect 189 203 190 204 
rect 189 204 190 205 
rect 189 205 190 206 
rect 189 206 190 207 
rect 189 207 190 208 
rect 189 218 190 219 
rect 189 219 190 220 
rect 189 220 190 221 
rect 189 221 190 222 
rect 189 222 190 223 
rect 189 223 190 224 
rect 189 234 190 235 
rect 189 235 190 236 
rect 189 236 190 237 
rect 189 237 190 238 
rect 189 238 190 239 
rect 189 239 190 240 
rect 189 250 190 251 
rect 189 251 190 252 
rect 189 252 190 253 
rect 189 253 190 254 
rect 189 254 190 255 
rect 189 255 190 256 
rect 189 266 190 267 
rect 189 267 190 268 
rect 189 268 190 269 
rect 189 269 190 270 
rect 189 270 190 271 
rect 189 271 190 272 
rect 189 282 190 283 
rect 189 283 190 284 
rect 189 284 190 285 
rect 189 285 190 286 
rect 189 286 190 287 
rect 189 287 190 288 
rect 189 298 190 299 
rect 189 299 190 300 
rect 189 300 190 301 
rect 189 301 190 302 
rect 189 302 190 303 
rect 189 303 190 304 
rect 190 10 191 11 
rect 190 11 191 12 
rect 190 12 191 13 
rect 190 13 191 14 
rect 190 14 191 15 
rect 190 15 191 16 
rect 190 26 191 27 
rect 190 27 191 28 
rect 190 28 191 29 
rect 190 29 191 30 
rect 190 30 191 31 
rect 190 31 191 32 
rect 190 42 191 43 
rect 190 43 191 44 
rect 190 44 191 45 
rect 190 45 191 46 
rect 190 46 191 47 
rect 190 47 191 48 
rect 190 58 191 59 
rect 190 59 191 60 
rect 190 60 191 61 
rect 190 61 191 62 
rect 190 62 191 63 
rect 190 63 191 64 
rect 190 74 191 75 
rect 190 75 191 76 
rect 190 76 191 77 
rect 190 77 191 78 
rect 190 78 191 79 
rect 190 79 191 80 
rect 190 90 191 91 
rect 190 91 191 92 
rect 190 92 191 93 
rect 190 93 191 94 
rect 190 94 191 95 
rect 190 95 191 96 
rect 190 106 191 107 
rect 190 107 191 108 
rect 190 108 191 109 
rect 190 109 191 110 
rect 190 110 191 111 
rect 190 111 191 112 
rect 190 122 191 123 
rect 190 123 191 124 
rect 190 124 191 125 
rect 190 125 191 126 
rect 190 126 191 127 
rect 190 127 191 128 
rect 190 138 191 139 
rect 190 139 191 140 
rect 190 140 191 141 
rect 190 141 191 142 
rect 190 142 191 143 
rect 190 143 191 144 
rect 190 154 191 155 
rect 190 155 191 156 
rect 190 156 191 157 
rect 190 157 191 158 
rect 190 158 191 159 
rect 190 159 191 160 
rect 190 170 191 171 
rect 190 171 191 172 
rect 190 172 191 173 
rect 190 173 191 174 
rect 190 174 191 175 
rect 190 175 191 176 
rect 190 186 191 187 
rect 190 187 191 188 
rect 190 188 191 189 
rect 190 189 191 190 
rect 190 190 191 191 
rect 190 191 191 192 
rect 190 202 191 203 
rect 190 203 191 204 
rect 190 204 191 205 
rect 190 205 191 206 
rect 190 206 191 207 
rect 190 207 191 208 
rect 190 218 191 219 
rect 190 219 191 220 
rect 190 220 191 221 
rect 190 221 191 222 
rect 190 222 191 223 
rect 190 223 191 224 
rect 190 234 191 235 
rect 190 235 191 236 
rect 190 236 191 237 
rect 190 237 191 238 
rect 190 238 191 239 
rect 190 239 191 240 
rect 190 250 191 251 
rect 190 251 191 252 
rect 190 252 191 253 
rect 190 253 191 254 
rect 190 254 191 255 
rect 190 255 191 256 
rect 190 266 191 267 
rect 190 267 191 268 
rect 190 268 191 269 
rect 190 269 191 270 
rect 190 270 191 271 
rect 190 271 191 272 
rect 190 282 191 283 
rect 190 283 191 284 
rect 190 284 191 285 
rect 190 285 191 286 
rect 190 286 191 287 
rect 190 287 191 288 
rect 190 298 191 299 
rect 190 299 191 300 
rect 190 300 191 301 
rect 190 301 191 302 
rect 190 302 191 303 
rect 190 303 191 304 
rect 191 10 192 11 
rect 191 11 192 12 
rect 191 12 192 13 
rect 191 13 192 14 
rect 191 14 192 15 
rect 191 15 192 16 
rect 191 26 192 27 
rect 191 28 192 29 
rect 191 29 192 30 
rect 191 30 192 31 
rect 191 31 192 32 
rect 191 42 192 43 
rect 191 44 192 45 
rect 191 45 192 46 
rect 191 47 192 48 
rect 191 58 192 59 
rect 191 60 192 61 
rect 191 61 192 62 
rect 191 63 192 64 
rect 191 74 192 75 
rect 191 76 192 77 
rect 191 77 192 78 
rect 191 79 192 80 
rect 191 90 192 91 
rect 191 91 192 92 
rect 191 92 192 93 
rect 191 93 192 94 
rect 191 95 192 96 
rect 191 106 192 107 
rect 191 107 192 108 
rect 191 108 192 109 
rect 191 109 192 110 
rect 191 111 192 112 
rect 191 122 192 123 
rect 191 123 192 124 
rect 191 124 192 125 
rect 191 125 192 126 
rect 191 126 192 127 
rect 191 127 192 128 
rect 191 138 192 139 
rect 191 139 192 140 
rect 191 140 192 141 
rect 191 141 192 142 
rect 191 142 192 143 
rect 191 143 192 144 
rect 191 154 192 155 
rect 191 155 192 156 
rect 191 156 192 157 
rect 191 157 192 158 
rect 191 159 192 160 
rect 191 170 192 171 
rect 191 172 192 173 
rect 191 173 192 174 
rect 191 175 192 176 
rect 191 186 192 187 
rect 191 188 192 189 
rect 191 189 192 190 
rect 191 191 192 192 
rect 191 202 192 203 
rect 191 204 192 205 
rect 191 205 192 206 
rect 191 207 192 208 
rect 191 218 192 219 
rect 191 220 192 221 
rect 191 221 192 222 
rect 191 222 192 223 
rect 191 223 192 224 
rect 191 234 192 235 
rect 191 235 192 236 
rect 191 236 192 237 
rect 191 237 192 238 
rect 191 239 192 240 
rect 191 250 192 251 
rect 191 251 192 252 
rect 191 252 192 253 
rect 191 253 192 254 
rect 191 255 192 256 
rect 191 266 192 267 
rect 191 267 192 268 
rect 191 268 192 269 
rect 191 269 192 270 
rect 191 270 192 271 
rect 191 271 192 272 
rect 191 282 192 283 
rect 191 284 192 285 
rect 191 285 192 286 
rect 191 286 192 287 
rect 191 287 192 288 
rect 191 298 192 299 
rect 191 300 192 301 
rect 191 301 192 302 
rect 191 302 192 303 
rect 191 303 192 304 
rect 202 10 203 11 
rect 202 12 203 13 
rect 202 13 203 14 
rect 202 14 203 15 
rect 202 15 203 16 
rect 202 26 203 27 
rect 202 28 203 29 
rect 202 29 203 30 
rect 202 31 203 32 
rect 202 42 203 43 
rect 202 43 203 44 
rect 202 44 203 45 
rect 202 45 203 46 
rect 202 46 203 47 
rect 202 47 203 48 
rect 202 58 203 59 
rect 202 59 203 60 
rect 202 60 203 61 
rect 202 61 203 62 
rect 202 62 203 63 
rect 202 63 203 64 
rect 202 74 203 75 
rect 202 76 203 77 
rect 202 77 203 78 
rect 202 79 203 80 
rect 202 90 203 91 
rect 202 91 203 92 
rect 202 92 203 93 
rect 202 93 203 94 
rect 202 95 203 96 
rect 202 106 203 107 
rect 202 107 203 108 
rect 202 108 203 109 
rect 202 109 203 110 
rect 202 110 203 111 
rect 202 111 203 112 
rect 202 122 203 123 
rect 202 124 203 125 
rect 202 125 203 126 
rect 202 127 203 128 
rect 202 138 203 139 
rect 202 140 203 141 
rect 202 141 203 142 
rect 202 143 203 144 
rect 202 154 203 155 
rect 202 156 203 157 
rect 202 157 203 158 
rect 202 159 203 160 
rect 202 170 203 171 
rect 202 172 203 173 
rect 202 173 203 174 
rect 202 174 203 175 
rect 202 175 203 176 
rect 202 186 203 187 
rect 202 187 203 188 
rect 202 188 203 189 
rect 202 189 203 190 
rect 202 190 203 191 
rect 202 191 203 192 
rect 202 202 203 203 
rect 202 204 203 205 
rect 202 205 203 206 
rect 202 207 203 208 
rect 202 218 203 219 
rect 202 220 203 221 
rect 202 221 203 222 
rect 202 223 203 224 
rect 202 234 203 235 
rect 202 235 203 236 
rect 202 236 203 237 
rect 202 237 203 238 
rect 202 239 203 240 
rect 202 250 203 251 
rect 202 251 203 252 
rect 202 252 203 253 
rect 202 253 203 254 
rect 202 255 203 256 
rect 202 266 203 267 
rect 202 267 203 268 
rect 202 268 203 269 
rect 202 269 203 270 
rect 202 271 203 272 
rect 202 282 203 283 
rect 202 284 203 285 
rect 202 285 203 286 
rect 202 287 203 288 
rect 202 298 203 299 
rect 202 300 203 301 
rect 202 301 203 302 
rect 202 303 203 304 
rect 203 10 204 11 
rect 203 11 204 12 
rect 203 12 204 13 
rect 203 13 204 14 
rect 203 14 204 15 
rect 203 15 204 16 
rect 203 26 204 27 
rect 203 27 204 28 
rect 203 28 204 29 
rect 203 29 204 30 
rect 203 30 204 31 
rect 203 31 204 32 
rect 203 42 204 43 
rect 203 43 204 44 
rect 203 44 204 45 
rect 203 45 204 46 
rect 203 46 204 47 
rect 203 47 204 48 
rect 203 58 204 59 
rect 203 59 204 60 
rect 203 60 204 61 
rect 203 61 204 62 
rect 203 62 204 63 
rect 203 63 204 64 
rect 203 74 204 75 
rect 203 75 204 76 
rect 203 76 204 77 
rect 203 77 204 78 
rect 203 78 204 79 
rect 203 79 204 80 
rect 203 90 204 91 
rect 203 91 204 92 
rect 203 92 204 93 
rect 203 93 204 94 
rect 203 94 204 95 
rect 203 95 204 96 
rect 203 106 204 107 
rect 203 107 204 108 
rect 203 108 204 109 
rect 203 109 204 110 
rect 203 110 204 111 
rect 203 111 204 112 
rect 203 122 204 123 
rect 203 123 204 124 
rect 203 124 204 125 
rect 203 125 204 126 
rect 203 126 204 127 
rect 203 127 204 128 
rect 203 138 204 139 
rect 203 139 204 140 
rect 203 140 204 141 
rect 203 141 204 142 
rect 203 142 204 143 
rect 203 143 204 144 
rect 203 154 204 155 
rect 203 155 204 156 
rect 203 156 204 157 
rect 203 157 204 158 
rect 203 158 204 159 
rect 203 159 204 160 
rect 203 170 204 171 
rect 203 171 204 172 
rect 203 172 204 173 
rect 203 173 204 174 
rect 203 174 204 175 
rect 203 175 204 176 
rect 203 186 204 187 
rect 203 187 204 188 
rect 203 188 204 189 
rect 203 189 204 190 
rect 203 190 204 191 
rect 203 191 204 192 
rect 203 202 204 203 
rect 203 203 204 204 
rect 203 204 204 205 
rect 203 205 204 206 
rect 203 206 204 207 
rect 203 207 204 208 
rect 203 218 204 219 
rect 203 219 204 220 
rect 203 220 204 221 
rect 203 221 204 222 
rect 203 222 204 223 
rect 203 223 204 224 
rect 203 234 204 235 
rect 203 235 204 236 
rect 203 236 204 237 
rect 203 237 204 238 
rect 203 238 204 239 
rect 203 239 204 240 
rect 203 250 204 251 
rect 203 251 204 252 
rect 203 252 204 253 
rect 203 253 204 254 
rect 203 254 204 255 
rect 203 255 204 256 
rect 203 266 204 267 
rect 203 267 204 268 
rect 203 268 204 269 
rect 203 269 204 270 
rect 203 270 204 271 
rect 203 271 204 272 
rect 203 282 204 283 
rect 203 283 204 284 
rect 203 284 204 285 
rect 203 285 204 286 
rect 203 286 204 287 
rect 203 287 204 288 
rect 203 298 204 299 
rect 203 299 204 300 
rect 203 300 204 301 
rect 203 301 204 302 
rect 203 302 204 303 
rect 203 303 204 304 
rect 204 10 205 11 
rect 204 11 205 12 
rect 204 12 205 13 
rect 204 13 205 14 
rect 204 14 205 15 
rect 204 15 205 16 
rect 204 26 205 27 
rect 204 27 205 28 
rect 204 28 205 29 
rect 204 29 205 30 
rect 204 30 205 31 
rect 204 31 205 32 
rect 204 42 205 43 
rect 204 43 205 44 
rect 204 44 205 45 
rect 204 45 205 46 
rect 204 46 205 47 
rect 204 47 205 48 
rect 204 58 205 59 
rect 204 59 205 60 
rect 204 60 205 61 
rect 204 61 205 62 
rect 204 62 205 63 
rect 204 63 205 64 
rect 204 74 205 75 
rect 204 75 205 76 
rect 204 76 205 77 
rect 204 77 205 78 
rect 204 78 205 79 
rect 204 79 205 80 
rect 204 90 205 91 
rect 204 91 205 92 
rect 204 92 205 93 
rect 204 93 205 94 
rect 204 94 205 95 
rect 204 95 205 96 
rect 204 106 205 107 
rect 204 107 205 108 
rect 204 108 205 109 
rect 204 109 205 110 
rect 204 110 205 111 
rect 204 111 205 112 
rect 204 122 205 123 
rect 204 123 205 124 
rect 204 124 205 125 
rect 204 125 205 126 
rect 204 126 205 127 
rect 204 127 205 128 
rect 204 138 205 139 
rect 204 139 205 140 
rect 204 140 205 141 
rect 204 141 205 142 
rect 204 142 205 143 
rect 204 143 205 144 
rect 204 154 205 155 
rect 204 155 205 156 
rect 204 156 205 157 
rect 204 157 205 158 
rect 204 158 205 159 
rect 204 159 205 160 
rect 204 170 205 171 
rect 204 171 205 172 
rect 204 172 205 173 
rect 204 173 205 174 
rect 204 174 205 175 
rect 204 175 205 176 
rect 204 186 205 187 
rect 204 187 205 188 
rect 204 188 205 189 
rect 204 189 205 190 
rect 204 190 205 191 
rect 204 191 205 192 
rect 204 202 205 203 
rect 204 203 205 204 
rect 204 204 205 205 
rect 204 205 205 206 
rect 204 206 205 207 
rect 204 207 205 208 
rect 204 218 205 219 
rect 204 219 205 220 
rect 204 220 205 221 
rect 204 221 205 222 
rect 204 222 205 223 
rect 204 223 205 224 
rect 204 234 205 235 
rect 204 235 205 236 
rect 204 236 205 237 
rect 204 237 205 238 
rect 204 238 205 239 
rect 204 239 205 240 
rect 204 250 205 251 
rect 204 251 205 252 
rect 204 252 205 253 
rect 204 253 205 254 
rect 204 254 205 255 
rect 204 255 205 256 
rect 204 266 205 267 
rect 204 267 205 268 
rect 204 268 205 269 
rect 204 269 205 270 
rect 204 270 205 271 
rect 204 271 205 272 
rect 204 282 205 283 
rect 204 283 205 284 
rect 204 284 205 285 
rect 204 285 205 286 
rect 204 286 205 287 
rect 204 287 205 288 
rect 204 298 205 299 
rect 204 299 205 300 
rect 204 300 205 301 
rect 204 301 205 302 
rect 204 302 205 303 
rect 204 303 205 304 
rect 205 10 206 11 
rect 205 11 206 12 
rect 205 12 206 13 
rect 205 13 206 14 
rect 205 14 206 15 
rect 205 15 206 16 
rect 205 26 206 27 
rect 205 27 206 28 
rect 205 28 206 29 
rect 205 29 206 30 
rect 205 30 206 31 
rect 205 31 206 32 
rect 205 42 206 43 
rect 205 43 206 44 
rect 205 44 206 45 
rect 205 45 206 46 
rect 205 46 206 47 
rect 205 47 206 48 
rect 205 58 206 59 
rect 205 59 206 60 
rect 205 60 206 61 
rect 205 61 206 62 
rect 205 62 206 63 
rect 205 63 206 64 
rect 205 74 206 75 
rect 205 75 206 76 
rect 205 76 206 77 
rect 205 77 206 78 
rect 205 78 206 79 
rect 205 79 206 80 
rect 205 90 206 91 
rect 205 91 206 92 
rect 205 92 206 93 
rect 205 93 206 94 
rect 205 94 206 95 
rect 205 95 206 96 
rect 205 106 206 107 
rect 205 107 206 108 
rect 205 108 206 109 
rect 205 109 206 110 
rect 205 110 206 111 
rect 205 111 206 112 
rect 205 122 206 123 
rect 205 123 206 124 
rect 205 124 206 125 
rect 205 125 206 126 
rect 205 126 206 127 
rect 205 127 206 128 
rect 205 138 206 139 
rect 205 139 206 140 
rect 205 140 206 141 
rect 205 141 206 142 
rect 205 142 206 143 
rect 205 143 206 144 
rect 205 154 206 155 
rect 205 155 206 156 
rect 205 156 206 157 
rect 205 157 206 158 
rect 205 158 206 159 
rect 205 159 206 160 
rect 205 170 206 171 
rect 205 171 206 172 
rect 205 172 206 173 
rect 205 173 206 174 
rect 205 174 206 175 
rect 205 175 206 176 
rect 205 186 206 187 
rect 205 187 206 188 
rect 205 188 206 189 
rect 205 189 206 190 
rect 205 190 206 191 
rect 205 191 206 192 
rect 205 202 206 203 
rect 205 203 206 204 
rect 205 204 206 205 
rect 205 205 206 206 
rect 205 206 206 207 
rect 205 207 206 208 
rect 205 218 206 219 
rect 205 219 206 220 
rect 205 220 206 221 
rect 205 221 206 222 
rect 205 222 206 223 
rect 205 223 206 224 
rect 205 234 206 235 
rect 205 235 206 236 
rect 205 236 206 237 
rect 205 237 206 238 
rect 205 238 206 239 
rect 205 239 206 240 
rect 205 250 206 251 
rect 205 251 206 252 
rect 205 252 206 253 
rect 205 253 206 254 
rect 205 254 206 255 
rect 205 255 206 256 
rect 205 266 206 267 
rect 205 267 206 268 
rect 205 268 206 269 
rect 205 269 206 270 
rect 205 270 206 271 
rect 205 271 206 272 
rect 205 282 206 283 
rect 205 283 206 284 
rect 205 284 206 285 
rect 205 285 206 286 
rect 205 286 206 287 
rect 205 287 206 288 
rect 205 298 206 299 
rect 205 299 206 300 
rect 205 300 206 301 
rect 205 301 206 302 
rect 205 302 206 303 
rect 205 303 206 304 
rect 206 10 207 11 
rect 206 11 207 12 
rect 206 12 207 13 
rect 206 13 207 14 
rect 206 14 207 15 
rect 206 15 207 16 
rect 206 26 207 27 
rect 206 27 207 28 
rect 206 28 207 29 
rect 206 29 207 30 
rect 206 30 207 31 
rect 206 31 207 32 
rect 206 42 207 43 
rect 206 43 207 44 
rect 206 44 207 45 
rect 206 45 207 46 
rect 206 46 207 47 
rect 206 47 207 48 
rect 206 58 207 59 
rect 206 59 207 60 
rect 206 60 207 61 
rect 206 61 207 62 
rect 206 62 207 63 
rect 206 63 207 64 
rect 206 74 207 75 
rect 206 75 207 76 
rect 206 76 207 77 
rect 206 77 207 78 
rect 206 78 207 79 
rect 206 79 207 80 
rect 206 90 207 91 
rect 206 91 207 92 
rect 206 92 207 93 
rect 206 93 207 94 
rect 206 94 207 95 
rect 206 95 207 96 
rect 206 106 207 107 
rect 206 107 207 108 
rect 206 108 207 109 
rect 206 109 207 110 
rect 206 110 207 111 
rect 206 111 207 112 
rect 206 122 207 123 
rect 206 123 207 124 
rect 206 124 207 125 
rect 206 125 207 126 
rect 206 126 207 127 
rect 206 127 207 128 
rect 206 138 207 139 
rect 206 139 207 140 
rect 206 140 207 141 
rect 206 141 207 142 
rect 206 142 207 143 
rect 206 143 207 144 
rect 206 154 207 155 
rect 206 155 207 156 
rect 206 156 207 157 
rect 206 157 207 158 
rect 206 158 207 159 
rect 206 159 207 160 
rect 206 170 207 171 
rect 206 171 207 172 
rect 206 172 207 173 
rect 206 173 207 174 
rect 206 174 207 175 
rect 206 175 207 176 
rect 206 186 207 187 
rect 206 187 207 188 
rect 206 188 207 189 
rect 206 189 207 190 
rect 206 190 207 191 
rect 206 191 207 192 
rect 206 202 207 203 
rect 206 203 207 204 
rect 206 204 207 205 
rect 206 205 207 206 
rect 206 206 207 207 
rect 206 207 207 208 
rect 206 218 207 219 
rect 206 219 207 220 
rect 206 220 207 221 
rect 206 221 207 222 
rect 206 222 207 223 
rect 206 223 207 224 
rect 206 234 207 235 
rect 206 235 207 236 
rect 206 236 207 237 
rect 206 237 207 238 
rect 206 238 207 239 
rect 206 239 207 240 
rect 206 250 207 251 
rect 206 251 207 252 
rect 206 252 207 253 
rect 206 253 207 254 
rect 206 254 207 255 
rect 206 255 207 256 
rect 206 266 207 267 
rect 206 267 207 268 
rect 206 268 207 269 
rect 206 269 207 270 
rect 206 270 207 271 
rect 206 271 207 272 
rect 206 282 207 283 
rect 206 283 207 284 
rect 206 284 207 285 
rect 206 285 207 286 
rect 206 286 207 287 
rect 206 287 207 288 
rect 206 298 207 299 
rect 206 299 207 300 
rect 206 300 207 301 
rect 206 301 207 302 
rect 206 302 207 303 
rect 206 303 207 304 
rect 207 10 208 11 
rect 207 11 208 12 
rect 207 12 208 13 
rect 207 13 208 14 
rect 207 14 208 15 
rect 207 15 208 16 
rect 207 26 208 27 
rect 207 27 208 28 
rect 207 28 208 29 
rect 207 29 208 30 
rect 207 31 208 32 
rect 207 42 208 43 
rect 207 44 208 45 
rect 207 45 208 46 
rect 207 46 208 47 
rect 207 47 208 48 
rect 207 58 208 59 
rect 207 60 208 61 
rect 207 61 208 62 
rect 207 63 208 64 
rect 207 74 208 75 
rect 207 75 208 76 
rect 207 76 208 77 
rect 207 77 208 78 
rect 207 79 208 80 
rect 207 90 208 91 
rect 207 92 208 93 
rect 207 93 208 94 
rect 207 94 208 95 
rect 207 95 208 96 
rect 207 106 208 107 
rect 207 108 208 109 
rect 207 109 208 110 
rect 207 110 208 111 
rect 207 111 208 112 
rect 207 122 208 123 
rect 207 123 208 124 
rect 207 124 208 125 
rect 207 125 208 126 
rect 207 127 208 128 
rect 207 138 208 139 
rect 207 140 208 141 
rect 207 141 208 142 
rect 207 142 208 143 
rect 207 143 208 144 
rect 207 154 208 155 
rect 207 155 208 156 
rect 207 156 208 157 
rect 207 157 208 158 
rect 207 159 208 160 
rect 207 170 208 171 
rect 207 171 208 172 
rect 207 172 208 173 
rect 207 173 208 174 
rect 207 174 208 175 
rect 207 175 208 176 
rect 207 186 208 187 
rect 207 187 208 188 
rect 207 188 208 189 
rect 207 189 208 190 
rect 207 191 208 192 
rect 207 202 208 203 
rect 207 203 208 204 
rect 207 204 208 205 
rect 207 205 208 206 
rect 207 207 208 208 
rect 207 218 208 219 
rect 207 219 208 220 
rect 207 220 208 221 
rect 207 221 208 222 
rect 207 223 208 224 
rect 207 234 208 235 
rect 207 236 208 237 
rect 207 237 208 238 
rect 207 238 208 239 
rect 207 239 208 240 
rect 207 250 208 251 
rect 207 251 208 252 
rect 207 252 208 253 
rect 207 253 208 254 
rect 207 254 208 255 
rect 207 255 208 256 
rect 207 266 208 267 
rect 207 267 208 268 
rect 207 268 208 269 
rect 207 269 208 270 
rect 207 271 208 272 
rect 207 282 208 283 
rect 207 284 208 285 
rect 207 285 208 286 
rect 207 286 208 287 
rect 207 287 208 288 
rect 207 298 208 299 
rect 207 300 208 301 
rect 207 301 208 302 
rect 207 302 208 303 
rect 207 303 208 304 
rect 218 10 219 11 
rect 218 11 219 12 
rect 218 12 219 13 
rect 218 13 219 14 
rect 218 15 219 16 
rect 218 26 219 27 
rect 218 27 219 28 
rect 218 28 219 29 
rect 218 29 219 30 
rect 218 30 219 31 
rect 218 31 219 32 
rect 218 42 219 43 
rect 218 44 219 45 
rect 218 45 219 46 
rect 218 47 219 48 
rect 218 58 219 59 
rect 218 60 219 61 
rect 218 61 219 62 
rect 218 63 219 64 
rect 218 74 219 75 
rect 218 75 219 76 
rect 218 76 219 77 
rect 218 77 219 78 
rect 218 79 219 80 
rect 218 90 219 91 
rect 218 91 219 92 
rect 218 92 219 93 
rect 218 93 219 94 
rect 218 94 219 95 
rect 218 95 219 96 
rect 218 106 219 107 
rect 218 107 219 108 
rect 218 108 219 109 
rect 218 109 219 110 
rect 218 110 219 111 
rect 218 111 219 112 
rect 218 122 219 123 
rect 218 123 219 124 
rect 218 124 219 125 
rect 218 125 219 126 
rect 218 126 219 127 
rect 218 127 219 128 
rect 218 138 219 139 
rect 218 140 219 141 
rect 218 141 219 142 
rect 218 143 219 144 
rect 218 154 219 155 
rect 218 156 219 157 
rect 218 157 219 158 
rect 218 158 219 159 
rect 218 159 219 160 
rect 218 170 219 171 
rect 218 171 219 172 
rect 218 172 219 173 
rect 218 173 219 174 
rect 218 175 219 176 
rect 218 186 219 187 
rect 218 187 219 188 
rect 218 188 219 189 
rect 218 189 219 190 
rect 218 190 219 191 
rect 218 191 219 192 
rect 218 202 219 203 
rect 218 204 219 205 
rect 218 205 219 206 
rect 218 207 219 208 
rect 218 218 219 219 
rect 218 219 219 220 
rect 218 220 219 221 
rect 218 221 219 222 
rect 218 222 219 223 
rect 218 223 219 224 
rect 218 234 219 235 
rect 218 235 219 236 
rect 218 236 219 237 
rect 218 237 219 238 
rect 218 239 219 240 
rect 218 250 219 251 
rect 218 252 219 253 
rect 218 253 219 254 
rect 218 254 219 255 
rect 218 255 219 256 
rect 218 266 219 267 
rect 218 267 219 268 
rect 218 268 219 269 
rect 218 269 219 270 
rect 218 271 219 272 
rect 218 282 219 283 
rect 218 284 219 285 
rect 218 285 219 286 
rect 218 287 219 288 
rect 218 298 219 299 
rect 218 300 219 301 
rect 218 301 219 302 
rect 218 302 219 303 
rect 218 303 219 304 
rect 219 10 220 11 
rect 219 11 220 12 
rect 219 12 220 13 
rect 219 13 220 14 
rect 219 14 220 15 
rect 219 15 220 16 
rect 219 26 220 27 
rect 219 27 220 28 
rect 219 28 220 29 
rect 219 29 220 30 
rect 219 30 220 31 
rect 219 31 220 32 
rect 219 42 220 43 
rect 219 43 220 44 
rect 219 44 220 45 
rect 219 45 220 46 
rect 219 46 220 47 
rect 219 47 220 48 
rect 219 58 220 59 
rect 219 59 220 60 
rect 219 60 220 61 
rect 219 61 220 62 
rect 219 62 220 63 
rect 219 63 220 64 
rect 219 74 220 75 
rect 219 75 220 76 
rect 219 76 220 77 
rect 219 77 220 78 
rect 219 78 220 79 
rect 219 79 220 80 
rect 219 90 220 91 
rect 219 91 220 92 
rect 219 92 220 93 
rect 219 93 220 94 
rect 219 94 220 95 
rect 219 95 220 96 
rect 219 106 220 107 
rect 219 107 220 108 
rect 219 108 220 109 
rect 219 109 220 110 
rect 219 110 220 111 
rect 219 111 220 112 
rect 219 122 220 123 
rect 219 123 220 124 
rect 219 124 220 125 
rect 219 125 220 126 
rect 219 126 220 127 
rect 219 127 220 128 
rect 219 138 220 139 
rect 219 139 220 140 
rect 219 140 220 141 
rect 219 141 220 142 
rect 219 142 220 143 
rect 219 143 220 144 
rect 219 154 220 155 
rect 219 155 220 156 
rect 219 156 220 157 
rect 219 157 220 158 
rect 219 158 220 159 
rect 219 159 220 160 
rect 219 170 220 171 
rect 219 171 220 172 
rect 219 172 220 173 
rect 219 173 220 174 
rect 219 174 220 175 
rect 219 175 220 176 
rect 219 186 220 187 
rect 219 187 220 188 
rect 219 188 220 189 
rect 219 189 220 190 
rect 219 190 220 191 
rect 219 191 220 192 
rect 219 202 220 203 
rect 219 203 220 204 
rect 219 204 220 205 
rect 219 205 220 206 
rect 219 206 220 207 
rect 219 207 220 208 
rect 219 218 220 219 
rect 219 219 220 220 
rect 219 220 220 221 
rect 219 221 220 222 
rect 219 222 220 223 
rect 219 223 220 224 
rect 219 234 220 235 
rect 219 235 220 236 
rect 219 236 220 237 
rect 219 237 220 238 
rect 219 238 220 239 
rect 219 239 220 240 
rect 219 250 220 251 
rect 219 251 220 252 
rect 219 252 220 253 
rect 219 253 220 254 
rect 219 254 220 255 
rect 219 255 220 256 
rect 219 266 220 267 
rect 219 267 220 268 
rect 219 268 220 269 
rect 219 269 220 270 
rect 219 270 220 271 
rect 219 271 220 272 
rect 219 282 220 283 
rect 219 283 220 284 
rect 219 284 220 285 
rect 219 285 220 286 
rect 219 286 220 287 
rect 219 287 220 288 
rect 219 298 220 299 
rect 219 299 220 300 
rect 219 300 220 301 
rect 219 301 220 302 
rect 219 302 220 303 
rect 219 303 220 304 
rect 220 10 221 11 
rect 220 11 221 12 
rect 220 12 221 13 
rect 220 13 221 14 
rect 220 14 221 15 
rect 220 15 221 16 
rect 220 26 221 27 
rect 220 27 221 28 
rect 220 28 221 29 
rect 220 29 221 30 
rect 220 30 221 31 
rect 220 31 221 32 
rect 220 42 221 43 
rect 220 43 221 44 
rect 220 44 221 45 
rect 220 45 221 46 
rect 220 46 221 47 
rect 220 47 221 48 
rect 220 58 221 59 
rect 220 59 221 60 
rect 220 60 221 61 
rect 220 61 221 62 
rect 220 62 221 63 
rect 220 63 221 64 
rect 220 74 221 75 
rect 220 75 221 76 
rect 220 76 221 77 
rect 220 77 221 78 
rect 220 78 221 79 
rect 220 79 221 80 
rect 220 90 221 91 
rect 220 91 221 92 
rect 220 92 221 93 
rect 220 93 221 94 
rect 220 94 221 95 
rect 220 95 221 96 
rect 220 106 221 107 
rect 220 107 221 108 
rect 220 108 221 109 
rect 220 109 221 110 
rect 220 110 221 111 
rect 220 111 221 112 
rect 220 122 221 123 
rect 220 123 221 124 
rect 220 124 221 125 
rect 220 125 221 126 
rect 220 126 221 127 
rect 220 127 221 128 
rect 220 138 221 139 
rect 220 139 221 140 
rect 220 140 221 141 
rect 220 141 221 142 
rect 220 142 221 143 
rect 220 143 221 144 
rect 220 154 221 155 
rect 220 155 221 156 
rect 220 156 221 157 
rect 220 157 221 158 
rect 220 158 221 159 
rect 220 159 221 160 
rect 220 170 221 171 
rect 220 171 221 172 
rect 220 172 221 173 
rect 220 173 221 174 
rect 220 174 221 175 
rect 220 175 221 176 
rect 220 186 221 187 
rect 220 187 221 188 
rect 220 188 221 189 
rect 220 189 221 190 
rect 220 190 221 191 
rect 220 191 221 192 
rect 220 202 221 203 
rect 220 203 221 204 
rect 220 204 221 205 
rect 220 205 221 206 
rect 220 206 221 207 
rect 220 207 221 208 
rect 220 218 221 219 
rect 220 219 221 220 
rect 220 220 221 221 
rect 220 221 221 222 
rect 220 222 221 223 
rect 220 223 221 224 
rect 220 234 221 235 
rect 220 235 221 236 
rect 220 236 221 237 
rect 220 237 221 238 
rect 220 238 221 239 
rect 220 239 221 240 
rect 220 250 221 251 
rect 220 251 221 252 
rect 220 252 221 253 
rect 220 253 221 254 
rect 220 254 221 255 
rect 220 255 221 256 
rect 220 266 221 267 
rect 220 267 221 268 
rect 220 268 221 269 
rect 220 269 221 270 
rect 220 270 221 271 
rect 220 271 221 272 
rect 220 282 221 283 
rect 220 283 221 284 
rect 220 284 221 285 
rect 220 285 221 286 
rect 220 286 221 287 
rect 220 287 221 288 
rect 220 298 221 299 
rect 220 299 221 300 
rect 220 300 221 301 
rect 220 301 221 302 
rect 220 302 221 303 
rect 220 303 221 304 
rect 221 10 222 11 
rect 221 11 222 12 
rect 221 12 222 13 
rect 221 13 222 14 
rect 221 14 222 15 
rect 221 15 222 16 
rect 221 26 222 27 
rect 221 27 222 28 
rect 221 28 222 29 
rect 221 29 222 30 
rect 221 30 222 31 
rect 221 31 222 32 
rect 221 42 222 43 
rect 221 43 222 44 
rect 221 44 222 45 
rect 221 45 222 46 
rect 221 46 222 47 
rect 221 47 222 48 
rect 221 58 222 59 
rect 221 59 222 60 
rect 221 60 222 61 
rect 221 61 222 62 
rect 221 62 222 63 
rect 221 63 222 64 
rect 221 74 222 75 
rect 221 75 222 76 
rect 221 76 222 77 
rect 221 77 222 78 
rect 221 78 222 79 
rect 221 79 222 80 
rect 221 90 222 91 
rect 221 91 222 92 
rect 221 92 222 93 
rect 221 93 222 94 
rect 221 94 222 95 
rect 221 95 222 96 
rect 221 106 222 107 
rect 221 107 222 108 
rect 221 108 222 109 
rect 221 109 222 110 
rect 221 110 222 111 
rect 221 111 222 112 
rect 221 122 222 123 
rect 221 123 222 124 
rect 221 124 222 125 
rect 221 125 222 126 
rect 221 126 222 127 
rect 221 127 222 128 
rect 221 138 222 139 
rect 221 139 222 140 
rect 221 140 222 141 
rect 221 141 222 142 
rect 221 142 222 143 
rect 221 143 222 144 
rect 221 154 222 155 
rect 221 155 222 156 
rect 221 156 222 157 
rect 221 157 222 158 
rect 221 158 222 159 
rect 221 159 222 160 
rect 221 170 222 171 
rect 221 171 222 172 
rect 221 172 222 173 
rect 221 173 222 174 
rect 221 174 222 175 
rect 221 175 222 176 
rect 221 186 222 187 
rect 221 187 222 188 
rect 221 188 222 189 
rect 221 189 222 190 
rect 221 190 222 191 
rect 221 191 222 192 
rect 221 202 222 203 
rect 221 203 222 204 
rect 221 204 222 205 
rect 221 205 222 206 
rect 221 206 222 207 
rect 221 207 222 208 
rect 221 218 222 219 
rect 221 219 222 220 
rect 221 220 222 221 
rect 221 221 222 222 
rect 221 222 222 223 
rect 221 223 222 224 
rect 221 234 222 235 
rect 221 235 222 236 
rect 221 236 222 237 
rect 221 237 222 238 
rect 221 238 222 239 
rect 221 239 222 240 
rect 221 250 222 251 
rect 221 251 222 252 
rect 221 252 222 253 
rect 221 253 222 254 
rect 221 254 222 255 
rect 221 255 222 256 
rect 221 266 222 267 
rect 221 267 222 268 
rect 221 268 222 269 
rect 221 269 222 270 
rect 221 270 222 271 
rect 221 271 222 272 
rect 221 282 222 283 
rect 221 283 222 284 
rect 221 284 222 285 
rect 221 285 222 286 
rect 221 286 222 287 
rect 221 287 222 288 
rect 221 298 222 299 
rect 221 299 222 300 
rect 221 300 222 301 
rect 221 301 222 302 
rect 221 302 222 303 
rect 221 303 222 304 
rect 222 10 223 11 
rect 222 11 223 12 
rect 222 12 223 13 
rect 222 13 223 14 
rect 222 14 223 15 
rect 222 15 223 16 
rect 222 26 223 27 
rect 222 27 223 28 
rect 222 28 223 29 
rect 222 29 223 30 
rect 222 30 223 31 
rect 222 31 223 32 
rect 222 42 223 43 
rect 222 43 223 44 
rect 222 44 223 45 
rect 222 45 223 46 
rect 222 46 223 47 
rect 222 47 223 48 
rect 222 58 223 59 
rect 222 59 223 60 
rect 222 60 223 61 
rect 222 61 223 62 
rect 222 62 223 63 
rect 222 63 223 64 
rect 222 74 223 75 
rect 222 75 223 76 
rect 222 76 223 77 
rect 222 77 223 78 
rect 222 78 223 79 
rect 222 79 223 80 
rect 222 90 223 91 
rect 222 91 223 92 
rect 222 92 223 93 
rect 222 93 223 94 
rect 222 94 223 95 
rect 222 95 223 96 
rect 222 106 223 107 
rect 222 107 223 108 
rect 222 108 223 109 
rect 222 109 223 110 
rect 222 110 223 111 
rect 222 111 223 112 
rect 222 122 223 123 
rect 222 123 223 124 
rect 222 124 223 125 
rect 222 125 223 126 
rect 222 126 223 127 
rect 222 127 223 128 
rect 222 138 223 139 
rect 222 139 223 140 
rect 222 140 223 141 
rect 222 141 223 142 
rect 222 142 223 143 
rect 222 143 223 144 
rect 222 154 223 155 
rect 222 155 223 156 
rect 222 156 223 157 
rect 222 157 223 158 
rect 222 158 223 159 
rect 222 159 223 160 
rect 222 170 223 171 
rect 222 171 223 172 
rect 222 172 223 173 
rect 222 173 223 174 
rect 222 174 223 175 
rect 222 175 223 176 
rect 222 186 223 187 
rect 222 187 223 188 
rect 222 188 223 189 
rect 222 189 223 190 
rect 222 190 223 191 
rect 222 191 223 192 
rect 222 202 223 203 
rect 222 203 223 204 
rect 222 204 223 205 
rect 222 205 223 206 
rect 222 206 223 207 
rect 222 207 223 208 
rect 222 218 223 219 
rect 222 219 223 220 
rect 222 220 223 221 
rect 222 221 223 222 
rect 222 222 223 223 
rect 222 223 223 224 
rect 222 234 223 235 
rect 222 235 223 236 
rect 222 236 223 237 
rect 222 237 223 238 
rect 222 238 223 239 
rect 222 239 223 240 
rect 222 250 223 251 
rect 222 251 223 252 
rect 222 252 223 253 
rect 222 253 223 254 
rect 222 254 223 255 
rect 222 255 223 256 
rect 222 266 223 267 
rect 222 267 223 268 
rect 222 268 223 269 
rect 222 269 223 270 
rect 222 270 223 271 
rect 222 271 223 272 
rect 222 282 223 283 
rect 222 283 223 284 
rect 222 284 223 285 
rect 222 285 223 286 
rect 222 286 223 287 
rect 222 287 223 288 
rect 222 298 223 299 
rect 222 299 223 300 
rect 222 300 223 301 
rect 222 301 223 302 
rect 222 302 223 303 
rect 222 303 223 304 
rect 223 10 224 11 
rect 223 11 224 12 
rect 223 12 224 13 
rect 223 13 224 14 
rect 223 14 224 15 
rect 223 15 224 16 
rect 223 26 224 27 
rect 223 28 224 29 
rect 223 29 224 30 
rect 223 30 224 31 
rect 223 31 224 32 
rect 223 42 224 43 
rect 223 44 224 45 
rect 223 45 224 46 
rect 223 47 224 48 
rect 223 58 224 59 
rect 223 59 224 60 
rect 223 60 224 61 
rect 223 61 224 62 
rect 223 63 224 64 
rect 223 74 224 75 
rect 223 76 224 77 
rect 223 77 224 78 
rect 223 78 224 79 
rect 223 79 224 80 
rect 223 90 224 91 
rect 223 92 224 93 
rect 223 93 224 94 
rect 223 95 224 96 
rect 223 106 224 107 
rect 223 108 224 109 
rect 223 109 224 110 
rect 223 111 224 112 
rect 223 122 224 123 
rect 223 124 224 125 
rect 223 125 224 126 
rect 223 127 224 128 
rect 223 138 224 139 
rect 223 140 224 141 
rect 223 141 224 142 
rect 223 142 224 143 
rect 223 143 224 144 
rect 223 154 224 155 
rect 223 156 224 157 
rect 223 157 224 158 
rect 223 159 224 160 
rect 223 170 224 171 
rect 223 171 224 172 
rect 223 172 224 173 
rect 223 173 224 174 
rect 223 174 224 175 
rect 223 175 224 176 
rect 223 186 224 187 
rect 223 188 224 189 
rect 223 189 224 190 
rect 223 190 224 191 
rect 223 191 224 192 
rect 223 202 224 203 
rect 223 204 224 205 
rect 223 205 224 206 
rect 223 206 224 207 
rect 223 207 224 208 
rect 223 218 224 219 
rect 223 220 224 221 
rect 223 221 224 222 
rect 223 223 224 224 
rect 223 234 224 235 
rect 223 236 224 237 
rect 223 237 224 238 
rect 223 238 224 239 
rect 223 239 224 240 
rect 223 250 224 251 
rect 223 252 224 253 
rect 223 253 224 254 
rect 223 254 224 255 
rect 223 255 224 256 
rect 223 266 224 267 
rect 223 267 224 268 
rect 223 268 224 269 
rect 223 269 224 270 
rect 223 271 224 272 
rect 223 282 224 283 
rect 223 284 224 285 
rect 223 285 224 286 
rect 223 286 224 287 
rect 223 287 224 288 
rect 223 298 224 299 
rect 223 300 224 301 
rect 223 301 224 302 
rect 223 303 224 304 
rect 234 10 235 11 
rect 234 11 235 12 
rect 234 12 235 13 
rect 234 13 235 14 
rect 234 14 235 15 
rect 234 15 235 16 
rect 234 26 235 27 
rect 234 28 235 29 
rect 234 29 235 30 
rect 234 31 235 32 
rect 234 42 235 43 
rect 234 43 235 44 
rect 234 44 235 45 
rect 234 45 235 46 
rect 234 47 235 48 
rect 234 58 235 59 
rect 234 60 235 61 
rect 234 61 235 62 
rect 234 62 235 63 
rect 234 63 235 64 
rect 234 74 235 75 
rect 234 76 235 77 
rect 234 77 235 78 
rect 234 79 235 80 
rect 234 90 235 91 
rect 234 92 235 93 
rect 234 93 235 94 
rect 234 94 235 95 
rect 234 95 235 96 
rect 234 106 235 107 
rect 234 108 235 109 
rect 234 109 235 110 
rect 234 110 235 111 
rect 234 111 235 112 
rect 234 122 235 123 
rect 234 124 235 125 
rect 234 125 235 126 
rect 234 126 235 127 
rect 234 127 235 128 
rect 234 138 235 139 
rect 234 139 235 140 
rect 234 140 235 141 
rect 234 141 235 142 
rect 234 143 235 144 
rect 234 154 235 155 
rect 234 156 235 157 
rect 234 157 235 158 
rect 234 159 235 160 
rect 234 170 235 171 
rect 234 172 235 173 
rect 234 173 235 174 
rect 234 175 235 176 
rect 234 186 235 187 
rect 234 188 235 189 
rect 234 189 235 190 
rect 234 191 235 192 
rect 234 202 235 203 
rect 234 204 235 205 
rect 234 205 235 206 
rect 234 207 235 208 
rect 234 218 235 219 
rect 234 220 235 221 
rect 234 221 235 222 
rect 234 222 235 223 
rect 234 223 235 224 
rect 234 234 235 235 
rect 234 236 235 237 
rect 234 237 235 238 
rect 234 238 235 239 
rect 234 239 235 240 
rect 234 250 235 251 
rect 234 252 235 253 
rect 234 253 235 254 
rect 234 254 235 255 
rect 234 255 235 256 
rect 234 266 235 267 
rect 234 268 235 269 
rect 234 269 235 270 
rect 234 271 235 272 
rect 234 282 235 283 
rect 234 283 235 284 
rect 234 284 235 285 
rect 234 285 235 286 
rect 234 287 235 288 
rect 234 298 235 299 
rect 234 299 235 300 
rect 234 300 235 301 
rect 234 301 235 302 
rect 234 303 235 304 
rect 235 10 236 11 
rect 235 11 236 12 
rect 235 12 236 13 
rect 235 13 236 14 
rect 235 14 236 15 
rect 235 15 236 16 
rect 235 26 236 27 
rect 235 27 236 28 
rect 235 28 236 29 
rect 235 29 236 30 
rect 235 30 236 31 
rect 235 31 236 32 
rect 235 42 236 43 
rect 235 43 236 44 
rect 235 44 236 45 
rect 235 45 236 46 
rect 235 46 236 47 
rect 235 47 236 48 
rect 235 58 236 59 
rect 235 59 236 60 
rect 235 60 236 61 
rect 235 61 236 62 
rect 235 62 236 63 
rect 235 63 236 64 
rect 235 74 236 75 
rect 235 75 236 76 
rect 235 76 236 77 
rect 235 77 236 78 
rect 235 78 236 79 
rect 235 79 236 80 
rect 235 90 236 91 
rect 235 91 236 92 
rect 235 92 236 93 
rect 235 93 236 94 
rect 235 94 236 95 
rect 235 95 236 96 
rect 235 106 236 107 
rect 235 107 236 108 
rect 235 108 236 109 
rect 235 109 236 110 
rect 235 110 236 111 
rect 235 111 236 112 
rect 235 122 236 123 
rect 235 123 236 124 
rect 235 124 236 125 
rect 235 125 236 126 
rect 235 126 236 127 
rect 235 127 236 128 
rect 235 138 236 139 
rect 235 139 236 140 
rect 235 140 236 141 
rect 235 141 236 142 
rect 235 142 236 143 
rect 235 143 236 144 
rect 235 154 236 155 
rect 235 155 236 156 
rect 235 156 236 157 
rect 235 157 236 158 
rect 235 158 236 159 
rect 235 159 236 160 
rect 235 170 236 171 
rect 235 171 236 172 
rect 235 172 236 173 
rect 235 173 236 174 
rect 235 174 236 175 
rect 235 175 236 176 
rect 235 186 236 187 
rect 235 187 236 188 
rect 235 188 236 189 
rect 235 189 236 190 
rect 235 190 236 191 
rect 235 191 236 192 
rect 235 202 236 203 
rect 235 203 236 204 
rect 235 204 236 205 
rect 235 205 236 206 
rect 235 206 236 207 
rect 235 207 236 208 
rect 235 218 236 219 
rect 235 219 236 220 
rect 235 220 236 221 
rect 235 221 236 222 
rect 235 222 236 223 
rect 235 223 236 224 
rect 235 234 236 235 
rect 235 235 236 236 
rect 235 236 236 237 
rect 235 237 236 238 
rect 235 238 236 239 
rect 235 239 236 240 
rect 235 250 236 251 
rect 235 251 236 252 
rect 235 252 236 253 
rect 235 253 236 254 
rect 235 254 236 255 
rect 235 255 236 256 
rect 235 266 236 267 
rect 235 267 236 268 
rect 235 268 236 269 
rect 235 269 236 270 
rect 235 270 236 271 
rect 235 271 236 272 
rect 235 282 236 283 
rect 235 283 236 284 
rect 235 284 236 285 
rect 235 285 236 286 
rect 235 286 236 287 
rect 235 287 236 288 
rect 235 298 236 299 
rect 235 299 236 300 
rect 235 300 236 301 
rect 235 301 236 302 
rect 235 302 236 303 
rect 235 303 236 304 
rect 236 10 237 11 
rect 236 11 237 12 
rect 236 12 237 13 
rect 236 13 237 14 
rect 236 14 237 15 
rect 236 15 237 16 
rect 236 26 237 27 
rect 236 27 237 28 
rect 236 28 237 29 
rect 236 29 237 30 
rect 236 30 237 31 
rect 236 31 237 32 
rect 236 42 237 43 
rect 236 43 237 44 
rect 236 44 237 45 
rect 236 45 237 46 
rect 236 46 237 47 
rect 236 47 237 48 
rect 236 58 237 59 
rect 236 59 237 60 
rect 236 60 237 61 
rect 236 61 237 62 
rect 236 62 237 63 
rect 236 63 237 64 
rect 236 74 237 75 
rect 236 75 237 76 
rect 236 76 237 77 
rect 236 77 237 78 
rect 236 78 237 79 
rect 236 79 237 80 
rect 236 90 237 91 
rect 236 91 237 92 
rect 236 92 237 93 
rect 236 93 237 94 
rect 236 94 237 95 
rect 236 95 237 96 
rect 236 106 237 107 
rect 236 107 237 108 
rect 236 108 237 109 
rect 236 109 237 110 
rect 236 110 237 111 
rect 236 111 237 112 
rect 236 122 237 123 
rect 236 123 237 124 
rect 236 124 237 125 
rect 236 125 237 126 
rect 236 126 237 127 
rect 236 127 237 128 
rect 236 138 237 139 
rect 236 139 237 140 
rect 236 140 237 141 
rect 236 141 237 142 
rect 236 142 237 143 
rect 236 143 237 144 
rect 236 154 237 155 
rect 236 155 237 156 
rect 236 156 237 157 
rect 236 157 237 158 
rect 236 158 237 159 
rect 236 159 237 160 
rect 236 170 237 171 
rect 236 171 237 172 
rect 236 172 237 173 
rect 236 173 237 174 
rect 236 174 237 175 
rect 236 175 237 176 
rect 236 186 237 187 
rect 236 187 237 188 
rect 236 188 237 189 
rect 236 189 237 190 
rect 236 190 237 191 
rect 236 191 237 192 
rect 236 202 237 203 
rect 236 203 237 204 
rect 236 204 237 205 
rect 236 205 237 206 
rect 236 206 237 207 
rect 236 207 237 208 
rect 236 218 237 219 
rect 236 219 237 220 
rect 236 220 237 221 
rect 236 221 237 222 
rect 236 222 237 223 
rect 236 223 237 224 
rect 236 234 237 235 
rect 236 235 237 236 
rect 236 236 237 237 
rect 236 237 237 238 
rect 236 238 237 239 
rect 236 239 237 240 
rect 236 250 237 251 
rect 236 251 237 252 
rect 236 252 237 253 
rect 236 253 237 254 
rect 236 254 237 255 
rect 236 255 237 256 
rect 236 266 237 267 
rect 236 267 237 268 
rect 236 268 237 269 
rect 236 269 237 270 
rect 236 270 237 271 
rect 236 271 237 272 
rect 236 282 237 283 
rect 236 283 237 284 
rect 236 284 237 285 
rect 236 285 237 286 
rect 236 286 237 287 
rect 236 287 237 288 
rect 236 298 237 299 
rect 236 299 237 300 
rect 236 300 237 301 
rect 236 301 237 302 
rect 236 302 237 303 
rect 236 303 237 304 
rect 237 10 238 11 
rect 237 11 238 12 
rect 237 12 238 13 
rect 237 13 238 14 
rect 237 14 238 15 
rect 237 15 238 16 
rect 237 26 238 27 
rect 237 27 238 28 
rect 237 28 238 29 
rect 237 29 238 30 
rect 237 30 238 31 
rect 237 31 238 32 
rect 237 42 238 43 
rect 237 43 238 44 
rect 237 44 238 45 
rect 237 45 238 46 
rect 237 46 238 47 
rect 237 47 238 48 
rect 237 58 238 59 
rect 237 59 238 60 
rect 237 60 238 61 
rect 237 61 238 62 
rect 237 62 238 63 
rect 237 63 238 64 
rect 237 74 238 75 
rect 237 75 238 76 
rect 237 76 238 77 
rect 237 77 238 78 
rect 237 78 238 79 
rect 237 79 238 80 
rect 237 90 238 91 
rect 237 91 238 92 
rect 237 92 238 93 
rect 237 93 238 94 
rect 237 94 238 95 
rect 237 95 238 96 
rect 237 106 238 107 
rect 237 107 238 108 
rect 237 108 238 109 
rect 237 109 238 110 
rect 237 110 238 111 
rect 237 111 238 112 
rect 237 122 238 123 
rect 237 123 238 124 
rect 237 124 238 125 
rect 237 125 238 126 
rect 237 126 238 127 
rect 237 127 238 128 
rect 237 138 238 139 
rect 237 139 238 140 
rect 237 140 238 141 
rect 237 141 238 142 
rect 237 142 238 143 
rect 237 143 238 144 
rect 237 154 238 155 
rect 237 155 238 156 
rect 237 156 238 157 
rect 237 157 238 158 
rect 237 158 238 159 
rect 237 159 238 160 
rect 237 170 238 171 
rect 237 171 238 172 
rect 237 172 238 173 
rect 237 173 238 174 
rect 237 174 238 175 
rect 237 175 238 176 
rect 237 186 238 187 
rect 237 187 238 188 
rect 237 188 238 189 
rect 237 189 238 190 
rect 237 190 238 191 
rect 237 191 238 192 
rect 237 202 238 203 
rect 237 203 238 204 
rect 237 204 238 205 
rect 237 205 238 206 
rect 237 206 238 207 
rect 237 207 238 208 
rect 237 218 238 219 
rect 237 219 238 220 
rect 237 220 238 221 
rect 237 221 238 222 
rect 237 222 238 223 
rect 237 223 238 224 
rect 237 234 238 235 
rect 237 235 238 236 
rect 237 236 238 237 
rect 237 237 238 238 
rect 237 238 238 239 
rect 237 239 238 240 
rect 237 250 238 251 
rect 237 251 238 252 
rect 237 252 238 253 
rect 237 253 238 254 
rect 237 254 238 255 
rect 237 255 238 256 
rect 237 266 238 267 
rect 237 267 238 268 
rect 237 268 238 269 
rect 237 269 238 270 
rect 237 270 238 271 
rect 237 271 238 272 
rect 237 282 238 283 
rect 237 283 238 284 
rect 237 284 238 285 
rect 237 285 238 286 
rect 237 286 238 287 
rect 237 287 238 288 
rect 237 298 238 299 
rect 237 299 238 300 
rect 237 300 238 301 
rect 237 301 238 302 
rect 237 302 238 303 
rect 237 303 238 304 
rect 238 10 239 11 
rect 238 11 239 12 
rect 238 12 239 13 
rect 238 13 239 14 
rect 238 14 239 15 
rect 238 15 239 16 
rect 238 26 239 27 
rect 238 27 239 28 
rect 238 28 239 29 
rect 238 29 239 30 
rect 238 30 239 31 
rect 238 31 239 32 
rect 238 42 239 43 
rect 238 43 239 44 
rect 238 44 239 45 
rect 238 45 239 46 
rect 238 46 239 47 
rect 238 47 239 48 
rect 238 58 239 59 
rect 238 59 239 60 
rect 238 60 239 61 
rect 238 61 239 62 
rect 238 62 239 63 
rect 238 63 239 64 
rect 238 74 239 75 
rect 238 75 239 76 
rect 238 76 239 77 
rect 238 77 239 78 
rect 238 78 239 79 
rect 238 79 239 80 
rect 238 90 239 91 
rect 238 91 239 92 
rect 238 92 239 93 
rect 238 93 239 94 
rect 238 94 239 95 
rect 238 95 239 96 
rect 238 106 239 107 
rect 238 107 239 108 
rect 238 108 239 109 
rect 238 109 239 110 
rect 238 110 239 111 
rect 238 111 239 112 
rect 238 122 239 123 
rect 238 123 239 124 
rect 238 124 239 125 
rect 238 125 239 126 
rect 238 126 239 127 
rect 238 127 239 128 
rect 238 138 239 139 
rect 238 139 239 140 
rect 238 140 239 141 
rect 238 141 239 142 
rect 238 142 239 143 
rect 238 143 239 144 
rect 238 154 239 155 
rect 238 155 239 156 
rect 238 156 239 157 
rect 238 157 239 158 
rect 238 158 239 159 
rect 238 159 239 160 
rect 238 170 239 171 
rect 238 171 239 172 
rect 238 172 239 173 
rect 238 173 239 174 
rect 238 174 239 175 
rect 238 175 239 176 
rect 238 186 239 187 
rect 238 187 239 188 
rect 238 188 239 189 
rect 238 189 239 190 
rect 238 190 239 191 
rect 238 191 239 192 
rect 238 202 239 203 
rect 238 203 239 204 
rect 238 204 239 205 
rect 238 205 239 206 
rect 238 206 239 207 
rect 238 207 239 208 
rect 238 218 239 219 
rect 238 219 239 220 
rect 238 220 239 221 
rect 238 221 239 222 
rect 238 222 239 223 
rect 238 223 239 224 
rect 238 234 239 235 
rect 238 235 239 236 
rect 238 236 239 237 
rect 238 237 239 238 
rect 238 238 239 239 
rect 238 239 239 240 
rect 238 250 239 251 
rect 238 251 239 252 
rect 238 252 239 253 
rect 238 253 239 254 
rect 238 254 239 255 
rect 238 255 239 256 
rect 238 266 239 267 
rect 238 267 239 268 
rect 238 268 239 269 
rect 238 269 239 270 
rect 238 270 239 271 
rect 238 271 239 272 
rect 238 282 239 283 
rect 238 283 239 284 
rect 238 284 239 285 
rect 238 285 239 286 
rect 238 286 239 287 
rect 238 287 239 288 
rect 238 298 239 299 
rect 238 299 239 300 
rect 238 300 239 301 
rect 238 301 239 302 
rect 238 302 239 303 
rect 238 303 239 304 
rect 239 10 240 11 
rect 239 11 240 12 
rect 239 12 240 13 
rect 239 13 240 14 
rect 239 15 240 16 
rect 239 26 240 27 
rect 239 28 240 29 
rect 239 29 240 30 
rect 239 30 240 31 
rect 239 31 240 32 
rect 239 42 240 43 
rect 239 43 240 44 
rect 239 44 240 45 
rect 239 45 240 46 
rect 239 46 240 47 
rect 239 47 240 48 
rect 239 58 240 59 
rect 239 59 240 60 
rect 239 60 240 61 
rect 239 61 240 62 
rect 239 63 240 64 
rect 239 74 240 75 
rect 239 75 240 76 
rect 239 76 240 77 
rect 239 77 240 78 
rect 239 78 240 79 
rect 239 79 240 80 
rect 239 90 240 91 
rect 239 91 240 92 
rect 239 92 240 93 
rect 239 93 240 94 
rect 239 94 240 95 
rect 239 95 240 96 
rect 239 106 240 107 
rect 239 108 240 109 
rect 239 109 240 110 
rect 239 111 240 112 
rect 239 122 240 123 
rect 239 124 240 125 
rect 239 125 240 126 
rect 239 126 240 127 
rect 239 127 240 128 
rect 239 138 240 139 
rect 239 139 240 140 
rect 239 140 240 141 
rect 239 141 240 142 
rect 239 142 240 143 
rect 239 143 240 144 
rect 239 154 240 155 
rect 239 155 240 156 
rect 239 156 240 157 
rect 239 157 240 158 
rect 239 159 240 160 
rect 239 170 240 171 
rect 239 171 240 172 
rect 239 172 240 173 
rect 239 173 240 174 
rect 239 175 240 176 
rect 239 186 240 187 
rect 239 188 240 189 
rect 239 189 240 190 
rect 239 190 240 191 
rect 239 191 240 192 
rect 239 202 240 203 
rect 239 203 240 204 
rect 239 204 240 205 
rect 239 205 240 206 
rect 239 207 240 208 
rect 239 218 240 219 
rect 239 220 240 221 
rect 239 221 240 222 
rect 239 223 240 224 
rect 239 234 240 235 
rect 239 235 240 236 
rect 239 236 240 237 
rect 239 237 240 238 
rect 239 239 240 240 
rect 239 250 240 251 
rect 239 252 240 253 
rect 239 253 240 254 
rect 239 255 240 256 
rect 239 266 240 267 
rect 239 267 240 268 
rect 239 268 240 269 
rect 239 269 240 270 
rect 239 270 240 271 
rect 239 271 240 272 
rect 239 282 240 283 
rect 239 283 240 284 
rect 239 284 240 285 
rect 239 285 240 286 
rect 239 287 240 288 
rect 239 298 240 299 
rect 239 299 240 300 
rect 239 300 240 301 
rect 239 301 240 302 
rect 239 302 240 303 
rect 239 303 240 304 
rect 250 10 251 11 
rect 250 11 251 12 
rect 250 12 251 13 
rect 250 13 251 14 
rect 250 15 251 16 
rect 250 26 251 27 
rect 250 28 251 29 
rect 250 29 251 30 
rect 250 30 251 31 
rect 250 31 251 32 
rect 250 42 251 43 
rect 250 44 251 45 
rect 250 45 251 46 
rect 250 46 251 47 
rect 250 47 251 48 
rect 250 58 251 59 
rect 250 59 251 60 
rect 250 60 251 61 
rect 250 61 251 62 
rect 250 62 251 63 
rect 250 63 251 64 
rect 250 74 251 75 
rect 250 76 251 77 
rect 250 77 251 78 
rect 250 78 251 79 
rect 250 79 251 80 
rect 250 90 251 91 
rect 250 92 251 93 
rect 250 93 251 94 
rect 250 95 251 96 
rect 250 106 251 107 
rect 250 108 251 109 
rect 250 109 251 110 
rect 250 110 251 111 
rect 250 111 251 112 
rect 250 122 251 123 
rect 250 124 251 125 
rect 250 125 251 126 
rect 250 127 251 128 
rect 250 138 251 139 
rect 250 140 251 141 
rect 250 141 251 142 
rect 250 142 251 143 
rect 250 143 251 144 
rect 250 154 251 155 
rect 250 155 251 156 
rect 250 156 251 157 
rect 250 157 251 158 
rect 250 159 251 160 
rect 250 170 251 171 
rect 250 171 251 172 
rect 250 172 251 173 
rect 250 173 251 174 
rect 250 174 251 175 
rect 250 175 251 176 
rect 250 186 251 187 
rect 250 188 251 189 
rect 250 189 251 190 
rect 250 190 251 191 
rect 250 191 251 192 
rect 250 202 251 203 
rect 250 204 251 205 
rect 250 205 251 206 
rect 250 207 251 208 
rect 250 218 251 219 
rect 250 219 251 220 
rect 250 220 251 221 
rect 250 221 251 222 
rect 250 222 251 223 
rect 250 223 251 224 
rect 250 234 251 235 
rect 250 235 251 236 
rect 250 236 251 237 
rect 250 237 251 238 
rect 250 239 251 240 
rect 250 250 251 251 
rect 250 251 251 252 
rect 250 252 251 253 
rect 250 253 251 254 
rect 250 255 251 256 
rect 250 266 251 267 
rect 250 268 251 269 
rect 250 269 251 270 
rect 250 271 251 272 
rect 250 282 251 283 
rect 250 284 251 285 
rect 250 285 251 286 
rect 250 286 251 287 
rect 250 287 251 288 
rect 250 298 251 299 
rect 250 300 251 301 
rect 250 301 251 302 
rect 250 302 251 303 
rect 250 303 251 304 
rect 251 10 252 11 
rect 251 11 252 12 
rect 251 12 252 13 
rect 251 13 252 14 
rect 251 14 252 15 
rect 251 15 252 16 
rect 251 26 252 27 
rect 251 27 252 28 
rect 251 28 252 29 
rect 251 29 252 30 
rect 251 30 252 31 
rect 251 31 252 32 
rect 251 42 252 43 
rect 251 43 252 44 
rect 251 44 252 45 
rect 251 45 252 46 
rect 251 46 252 47 
rect 251 47 252 48 
rect 251 58 252 59 
rect 251 59 252 60 
rect 251 60 252 61 
rect 251 61 252 62 
rect 251 62 252 63 
rect 251 63 252 64 
rect 251 74 252 75 
rect 251 75 252 76 
rect 251 76 252 77 
rect 251 77 252 78 
rect 251 78 252 79 
rect 251 79 252 80 
rect 251 90 252 91 
rect 251 91 252 92 
rect 251 92 252 93 
rect 251 93 252 94 
rect 251 94 252 95 
rect 251 95 252 96 
rect 251 106 252 107 
rect 251 107 252 108 
rect 251 108 252 109 
rect 251 109 252 110 
rect 251 110 252 111 
rect 251 111 252 112 
rect 251 122 252 123 
rect 251 123 252 124 
rect 251 124 252 125 
rect 251 125 252 126 
rect 251 126 252 127 
rect 251 127 252 128 
rect 251 138 252 139 
rect 251 139 252 140 
rect 251 140 252 141 
rect 251 141 252 142 
rect 251 142 252 143 
rect 251 143 252 144 
rect 251 154 252 155 
rect 251 155 252 156 
rect 251 156 252 157 
rect 251 157 252 158 
rect 251 158 252 159 
rect 251 159 252 160 
rect 251 170 252 171 
rect 251 171 252 172 
rect 251 172 252 173 
rect 251 173 252 174 
rect 251 174 252 175 
rect 251 175 252 176 
rect 251 186 252 187 
rect 251 187 252 188 
rect 251 188 252 189 
rect 251 189 252 190 
rect 251 190 252 191 
rect 251 191 252 192 
rect 251 202 252 203 
rect 251 203 252 204 
rect 251 204 252 205 
rect 251 205 252 206 
rect 251 206 252 207 
rect 251 207 252 208 
rect 251 218 252 219 
rect 251 219 252 220 
rect 251 220 252 221 
rect 251 221 252 222 
rect 251 222 252 223 
rect 251 223 252 224 
rect 251 234 252 235 
rect 251 235 252 236 
rect 251 236 252 237 
rect 251 237 252 238 
rect 251 238 252 239 
rect 251 239 252 240 
rect 251 250 252 251 
rect 251 251 252 252 
rect 251 252 252 253 
rect 251 253 252 254 
rect 251 254 252 255 
rect 251 255 252 256 
rect 251 266 252 267 
rect 251 267 252 268 
rect 251 268 252 269 
rect 251 269 252 270 
rect 251 270 252 271 
rect 251 271 252 272 
rect 251 282 252 283 
rect 251 283 252 284 
rect 251 284 252 285 
rect 251 285 252 286 
rect 251 286 252 287 
rect 251 287 252 288 
rect 251 298 252 299 
rect 251 299 252 300 
rect 251 300 252 301 
rect 251 301 252 302 
rect 251 302 252 303 
rect 251 303 252 304 
rect 252 10 253 11 
rect 252 11 253 12 
rect 252 12 253 13 
rect 252 13 253 14 
rect 252 14 253 15 
rect 252 15 253 16 
rect 252 26 253 27 
rect 252 27 253 28 
rect 252 28 253 29 
rect 252 29 253 30 
rect 252 30 253 31 
rect 252 31 253 32 
rect 252 42 253 43 
rect 252 43 253 44 
rect 252 44 253 45 
rect 252 45 253 46 
rect 252 46 253 47 
rect 252 47 253 48 
rect 252 58 253 59 
rect 252 59 253 60 
rect 252 60 253 61 
rect 252 61 253 62 
rect 252 62 253 63 
rect 252 63 253 64 
rect 252 74 253 75 
rect 252 75 253 76 
rect 252 76 253 77 
rect 252 77 253 78 
rect 252 78 253 79 
rect 252 79 253 80 
rect 252 90 253 91 
rect 252 91 253 92 
rect 252 92 253 93 
rect 252 93 253 94 
rect 252 94 253 95 
rect 252 95 253 96 
rect 252 106 253 107 
rect 252 107 253 108 
rect 252 108 253 109 
rect 252 109 253 110 
rect 252 110 253 111 
rect 252 111 253 112 
rect 252 122 253 123 
rect 252 123 253 124 
rect 252 124 253 125 
rect 252 125 253 126 
rect 252 126 253 127 
rect 252 127 253 128 
rect 252 138 253 139 
rect 252 139 253 140 
rect 252 140 253 141 
rect 252 141 253 142 
rect 252 142 253 143 
rect 252 143 253 144 
rect 252 154 253 155 
rect 252 155 253 156 
rect 252 156 253 157 
rect 252 157 253 158 
rect 252 158 253 159 
rect 252 159 253 160 
rect 252 170 253 171 
rect 252 171 253 172 
rect 252 172 253 173 
rect 252 173 253 174 
rect 252 174 253 175 
rect 252 175 253 176 
rect 252 186 253 187 
rect 252 187 253 188 
rect 252 188 253 189 
rect 252 189 253 190 
rect 252 190 253 191 
rect 252 191 253 192 
rect 252 202 253 203 
rect 252 203 253 204 
rect 252 204 253 205 
rect 252 205 253 206 
rect 252 206 253 207 
rect 252 207 253 208 
rect 252 218 253 219 
rect 252 219 253 220 
rect 252 220 253 221 
rect 252 221 253 222 
rect 252 222 253 223 
rect 252 223 253 224 
rect 252 234 253 235 
rect 252 235 253 236 
rect 252 236 253 237 
rect 252 237 253 238 
rect 252 238 253 239 
rect 252 239 253 240 
rect 252 250 253 251 
rect 252 251 253 252 
rect 252 252 253 253 
rect 252 253 253 254 
rect 252 254 253 255 
rect 252 255 253 256 
rect 252 266 253 267 
rect 252 267 253 268 
rect 252 268 253 269 
rect 252 269 253 270 
rect 252 270 253 271 
rect 252 271 253 272 
rect 252 282 253 283 
rect 252 283 253 284 
rect 252 284 253 285 
rect 252 285 253 286 
rect 252 286 253 287 
rect 252 287 253 288 
rect 252 298 253 299 
rect 252 299 253 300 
rect 252 300 253 301 
rect 252 301 253 302 
rect 252 302 253 303 
rect 252 303 253 304 
rect 253 10 254 11 
rect 253 11 254 12 
rect 253 12 254 13 
rect 253 13 254 14 
rect 253 14 254 15 
rect 253 15 254 16 
rect 253 26 254 27 
rect 253 27 254 28 
rect 253 28 254 29 
rect 253 29 254 30 
rect 253 30 254 31 
rect 253 31 254 32 
rect 253 42 254 43 
rect 253 43 254 44 
rect 253 44 254 45 
rect 253 45 254 46 
rect 253 46 254 47 
rect 253 47 254 48 
rect 253 58 254 59 
rect 253 59 254 60 
rect 253 60 254 61 
rect 253 61 254 62 
rect 253 62 254 63 
rect 253 63 254 64 
rect 253 74 254 75 
rect 253 75 254 76 
rect 253 76 254 77 
rect 253 77 254 78 
rect 253 78 254 79 
rect 253 79 254 80 
rect 253 90 254 91 
rect 253 91 254 92 
rect 253 92 254 93 
rect 253 93 254 94 
rect 253 94 254 95 
rect 253 95 254 96 
rect 253 106 254 107 
rect 253 107 254 108 
rect 253 108 254 109 
rect 253 109 254 110 
rect 253 110 254 111 
rect 253 111 254 112 
rect 253 122 254 123 
rect 253 123 254 124 
rect 253 124 254 125 
rect 253 125 254 126 
rect 253 126 254 127 
rect 253 127 254 128 
rect 253 138 254 139 
rect 253 139 254 140 
rect 253 140 254 141 
rect 253 141 254 142 
rect 253 142 254 143 
rect 253 143 254 144 
rect 253 154 254 155 
rect 253 155 254 156 
rect 253 156 254 157 
rect 253 157 254 158 
rect 253 158 254 159 
rect 253 159 254 160 
rect 253 170 254 171 
rect 253 171 254 172 
rect 253 172 254 173 
rect 253 173 254 174 
rect 253 174 254 175 
rect 253 175 254 176 
rect 253 186 254 187 
rect 253 187 254 188 
rect 253 188 254 189 
rect 253 189 254 190 
rect 253 190 254 191 
rect 253 191 254 192 
rect 253 202 254 203 
rect 253 203 254 204 
rect 253 204 254 205 
rect 253 205 254 206 
rect 253 206 254 207 
rect 253 207 254 208 
rect 253 218 254 219 
rect 253 219 254 220 
rect 253 220 254 221 
rect 253 221 254 222 
rect 253 222 254 223 
rect 253 223 254 224 
rect 253 234 254 235 
rect 253 235 254 236 
rect 253 236 254 237 
rect 253 237 254 238 
rect 253 238 254 239 
rect 253 239 254 240 
rect 253 250 254 251 
rect 253 251 254 252 
rect 253 252 254 253 
rect 253 253 254 254 
rect 253 254 254 255 
rect 253 255 254 256 
rect 253 266 254 267 
rect 253 267 254 268 
rect 253 268 254 269 
rect 253 269 254 270 
rect 253 270 254 271 
rect 253 271 254 272 
rect 253 282 254 283 
rect 253 283 254 284 
rect 253 284 254 285 
rect 253 285 254 286 
rect 253 286 254 287 
rect 253 287 254 288 
rect 253 298 254 299 
rect 253 299 254 300 
rect 253 300 254 301 
rect 253 301 254 302 
rect 253 302 254 303 
rect 253 303 254 304 
rect 254 10 255 11 
rect 254 11 255 12 
rect 254 12 255 13 
rect 254 13 255 14 
rect 254 14 255 15 
rect 254 15 255 16 
rect 254 26 255 27 
rect 254 27 255 28 
rect 254 28 255 29 
rect 254 29 255 30 
rect 254 30 255 31 
rect 254 31 255 32 
rect 254 42 255 43 
rect 254 43 255 44 
rect 254 44 255 45 
rect 254 45 255 46 
rect 254 46 255 47 
rect 254 47 255 48 
rect 254 58 255 59 
rect 254 59 255 60 
rect 254 60 255 61 
rect 254 61 255 62 
rect 254 62 255 63 
rect 254 63 255 64 
rect 254 74 255 75 
rect 254 75 255 76 
rect 254 76 255 77 
rect 254 77 255 78 
rect 254 78 255 79 
rect 254 79 255 80 
rect 254 90 255 91 
rect 254 91 255 92 
rect 254 92 255 93 
rect 254 93 255 94 
rect 254 94 255 95 
rect 254 95 255 96 
rect 254 106 255 107 
rect 254 107 255 108 
rect 254 108 255 109 
rect 254 109 255 110 
rect 254 110 255 111 
rect 254 111 255 112 
rect 254 122 255 123 
rect 254 123 255 124 
rect 254 124 255 125 
rect 254 125 255 126 
rect 254 126 255 127 
rect 254 127 255 128 
rect 254 138 255 139 
rect 254 139 255 140 
rect 254 140 255 141 
rect 254 141 255 142 
rect 254 142 255 143 
rect 254 143 255 144 
rect 254 154 255 155 
rect 254 155 255 156 
rect 254 156 255 157 
rect 254 157 255 158 
rect 254 158 255 159 
rect 254 159 255 160 
rect 254 170 255 171 
rect 254 171 255 172 
rect 254 172 255 173 
rect 254 173 255 174 
rect 254 174 255 175 
rect 254 175 255 176 
rect 254 186 255 187 
rect 254 187 255 188 
rect 254 188 255 189 
rect 254 189 255 190 
rect 254 190 255 191 
rect 254 191 255 192 
rect 254 202 255 203 
rect 254 203 255 204 
rect 254 204 255 205 
rect 254 205 255 206 
rect 254 206 255 207 
rect 254 207 255 208 
rect 254 218 255 219 
rect 254 219 255 220 
rect 254 220 255 221 
rect 254 221 255 222 
rect 254 222 255 223 
rect 254 223 255 224 
rect 254 234 255 235 
rect 254 235 255 236 
rect 254 236 255 237 
rect 254 237 255 238 
rect 254 238 255 239 
rect 254 239 255 240 
rect 254 250 255 251 
rect 254 251 255 252 
rect 254 252 255 253 
rect 254 253 255 254 
rect 254 254 255 255 
rect 254 255 255 256 
rect 254 266 255 267 
rect 254 267 255 268 
rect 254 268 255 269 
rect 254 269 255 270 
rect 254 270 255 271 
rect 254 271 255 272 
rect 254 282 255 283 
rect 254 283 255 284 
rect 254 284 255 285 
rect 254 285 255 286 
rect 254 286 255 287 
rect 254 287 255 288 
rect 254 298 255 299 
rect 254 299 255 300 
rect 254 300 255 301 
rect 254 301 255 302 
rect 254 302 255 303 
rect 254 303 255 304 
rect 255 10 256 11 
rect 255 11 256 12 
rect 255 12 256 13 
rect 255 13 256 14 
rect 255 14 256 15 
rect 255 15 256 16 
rect 255 26 256 27 
rect 255 27 256 28 
rect 255 28 256 29 
rect 255 29 256 30 
rect 255 30 256 31 
rect 255 31 256 32 
rect 255 42 256 43 
rect 255 44 256 45 
rect 255 45 256 46 
rect 255 46 256 47 
rect 255 47 256 48 
rect 255 58 256 59 
rect 255 60 256 61 
rect 255 61 256 62 
rect 255 62 256 63 
rect 255 63 256 64 
rect 255 74 256 75 
rect 255 75 256 76 
rect 255 76 256 77 
rect 255 77 256 78 
rect 255 78 256 79 
rect 255 79 256 80 
rect 255 90 256 91 
rect 255 91 256 92 
rect 255 92 256 93 
rect 255 93 256 94 
rect 255 94 256 95 
rect 255 95 256 96 
rect 255 106 256 107 
rect 255 108 256 109 
rect 255 109 256 110 
rect 255 111 256 112 
rect 255 122 256 123 
rect 255 123 256 124 
rect 255 124 256 125 
rect 255 125 256 126 
rect 255 127 256 128 
rect 255 138 256 139 
rect 255 140 256 141 
rect 255 141 256 142 
rect 255 142 256 143 
rect 255 143 256 144 
rect 255 154 256 155 
rect 255 155 256 156 
rect 255 156 256 157 
rect 255 157 256 158 
rect 255 158 256 159 
rect 255 159 256 160 
rect 255 170 256 171 
rect 255 172 256 173 
rect 255 173 256 174 
rect 255 174 256 175 
rect 255 175 256 176 
rect 255 186 256 187 
rect 255 188 256 189 
rect 255 189 256 190 
rect 255 190 256 191 
rect 255 191 256 192 
rect 255 202 256 203 
rect 255 204 256 205 
rect 255 205 256 206 
rect 255 207 256 208 
rect 255 218 256 219 
rect 255 220 256 221 
rect 255 221 256 222 
rect 255 222 256 223 
rect 255 223 256 224 
rect 255 234 256 235 
rect 255 235 256 236 
rect 255 236 256 237 
rect 255 237 256 238 
rect 255 238 256 239 
rect 255 239 256 240 
rect 255 250 256 251 
rect 255 252 256 253 
rect 255 253 256 254 
rect 255 254 256 255 
rect 255 255 256 256 
rect 255 266 256 267 
rect 255 268 256 269 
rect 255 269 256 270 
rect 255 270 256 271 
rect 255 271 256 272 
rect 255 282 256 283 
rect 255 283 256 284 
rect 255 284 256 285 
rect 255 285 256 286 
rect 255 286 256 287 
rect 255 287 256 288 
rect 255 298 256 299 
rect 255 299 256 300 
rect 255 300 256 301 
rect 255 301 256 302 
rect 255 302 256 303 
rect 255 303 256 304 
rect 266 10 267 11 
rect 266 12 267 13 
rect 266 13 267 14 
rect 266 14 267 15 
rect 266 15 267 16 
rect 266 26 267 27 
rect 266 28 267 29 
rect 266 29 267 30 
rect 266 30 267 31 
rect 266 31 267 32 
rect 266 42 267 43 
rect 266 44 267 45 
rect 266 45 267 46 
rect 266 47 267 48 
rect 266 58 267 59 
rect 266 59 267 60 
rect 266 60 267 61 
rect 266 61 267 62 
rect 266 63 267 64 
rect 266 74 267 75 
rect 266 75 267 76 
rect 266 76 267 77 
rect 266 77 267 78 
rect 266 78 267 79 
rect 266 79 267 80 
rect 266 90 267 91 
rect 266 92 267 93 
rect 266 93 267 94 
rect 266 94 267 95 
rect 266 95 267 96 
rect 266 106 267 107 
rect 266 108 267 109 
rect 266 109 267 110 
rect 266 110 267 111 
rect 266 111 267 112 
rect 266 122 267 123 
rect 266 124 267 125 
rect 266 125 267 126 
rect 266 126 267 127 
rect 266 127 267 128 
rect 266 138 267 139 
rect 266 140 267 141 
rect 266 141 267 142 
rect 266 142 267 143 
rect 266 143 267 144 
rect 266 154 267 155 
rect 266 155 267 156 
rect 266 156 267 157 
rect 266 157 267 158 
rect 266 158 267 159 
rect 266 159 267 160 
rect 266 170 267 171 
rect 266 171 267 172 
rect 266 172 267 173 
rect 266 173 267 174 
rect 266 175 267 176 
rect 266 186 267 187 
rect 266 188 267 189 
rect 266 189 267 190 
rect 266 191 267 192 
rect 266 202 267 203 
rect 266 204 267 205 
rect 266 205 267 206 
rect 266 207 267 208 
rect 266 218 267 219 
rect 266 219 267 220 
rect 266 220 267 221 
rect 266 221 267 222 
rect 266 222 267 223 
rect 266 223 267 224 
rect 266 234 267 235 
rect 266 236 267 237 
rect 266 237 267 238 
rect 266 239 267 240 
rect 266 250 267 251 
rect 266 251 267 252 
rect 266 252 267 253 
rect 266 253 267 254 
rect 266 255 267 256 
rect 266 266 267 267 
rect 266 268 267 269 
rect 266 269 267 270 
rect 266 270 267 271 
rect 266 271 267 272 
rect 266 282 267 283 
rect 266 284 267 285 
rect 266 285 267 286 
rect 266 286 267 287 
rect 266 287 267 288 
rect 266 298 267 299 
rect 266 300 267 301 
rect 266 301 267 302 
rect 266 303 267 304 
rect 267 10 268 11 
rect 267 11 268 12 
rect 267 12 268 13 
rect 267 13 268 14 
rect 267 14 268 15 
rect 267 15 268 16 
rect 267 26 268 27 
rect 267 27 268 28 
rect 267 28 268 29 
rect 267 29 268 30 
rect 267 30 268 31 
rect 267 31 268 32 
rect 267 42 268 43 
rect 267 43 268 44 
rect 267 44 268 45 
rect 267 45 268 46 
rect 267 46 268 47 
rect 267 47 268 48 
rect 267 58 268 59 
rect 267 59 268 60 
rect 267 60 268 61 
rect 267 61 268 62 
rect 267 62 268 63 
rect 267 63 268 64 
rect 267 74 268 75 
rect 267 75 268 76 
rect 267 76 268 77 
rect 267 77 268 78 
rect 267 78 268 79 
rect 267 79 268 80 
rect 267 90 268 91 
rect 267 91 268 92 
rect 267 92 268 93 
rect 267 93 268 94 
rect 267 94 268 95 
rect 267 95 268 96 
rect 267 106 268 107 
rect 267 107 268 108 
rect 267 108 268 109 
rect 267 109 268 110 
rect 267 110 268 111 
rect 267 111 268 112 
rect 267 122 268 123 
rect 267 123 268 124 
rect 267 124 268 125 
rect 267 125 268 126 
rect 267 126 268 127 
rect 267 127 268 128 
rect 267 138 268 139 
rect 267 139 268 140 
rect 267 140 268 141 
rect 267 141 268 142 
rect 267 142 268 143 
rect 267 143 268 144 
rect 267 154 268 155 
rect 267 155 268 156 
rect 267 156 268 157 
rect 267 157 268 158 
rect 267 158 268 159 
rect 267 159 268 160 
rect 267 170 268 171 
rect 267 171 268 172 
rect 267 172 268 173 
rect 267 173 268 174 
rect 267 174 268 175 
rect 267 175 268 176 
rect 267 186 268 187 
rect 267 187 268 188 
rect 267 188 268 189 
rect 267 189 268 190 
rect 267 190 268 191 
rect 267 191 268 192 
rect 267 202 268 203 
rect 267 203 268 204 
rect 267 204 268 205 
rect 267 205 268 206 
rect 267 206 268 207 
rect 267 207 268 208 
rect 267 218 268 219 
rect 267 219 268 220 
rect 267 220 268 221 
rect 267 221 268 222 
rect 267 222 268 223 
rect 267 223 268 224 
rect 267 234 268 235 
rect 267 235 268 236 
rect 267 236 268 237 
rect 267 237 268 238 
rect 267 238 268 239 
rect 267 239 268 240 
rect 267 250 268 251 
rect 267 251 268 252 
rect 267 252 268 253 
rect 267 253 268 254 
rect 267 254 268 255 
rect 267 255 268 256 
rect 267 266 268 267 
rect 267 267 268 268 
rect 267 268 268 269 
rect 267 269 268 270 
rect 267 270 268 271 
rect 267 271 268 272 
rect 267 282 268 283 
rect 267 283 268 284 
rect 267 284 268 285 
rect 267 285 268 286 
rect 267 286 268 287 
rect 267 287 268 288 
rect 267 298 268 299 
rect 267 299 268 300 
rect 267 300 268 301 
rect 267 301 268 302 
rect 267 302 268 303 
rect 267 303 268 304 
rect 268 10 269 11 
rect 268 11 269 12 
rect 268 12 269 13 
rect 268 13 269 14 
rect 268 14 269 15 
rect 268 15 269 16 
rect 268 26 269 27 
rect 268 27 269 28 
rect 268 28 269 29 
rect 268 29 269 30 
rect 268 30 269 31 
rect 268 31 269 32 
rect 268 42 269 43 
rect 268 43 269 44 
rect 268 44 269 45 
rect 268 45 269 46 
rect 268 46 269 47 
rect 268 47 269 48 
rect 268 58 269 59 
rect 268 59 269 60 
rect 268 60 269 61 
rect 268 61 269 62 
rect 268 62 269 63 
rect 268 63 269 64 
rect 268 74 269 75 
rect 268 75 269 76 
rect 268 76 269 77 
rect 268 77 269 78 
rect 268 78 269 79 
rect 268 79 269 80 
rect 268 90 269 91 
rect 268 91 269 92 
rect 268 92 269 93 
rect 268 93 269 94 
rect 268 94 269 95 
rect 268 95 269 96 
rect 268 106 269 107 
rect 268 107 269 108 
rect 268 108 269 109 
rect 268 109 269 110 
rect 268 110 269 111 
rect 268 111 269 112 
rect 268 122 269 123 
rect 268 123 269 124 
rect 268 124 269 125 
rect 268 125 269 126 
rect 268 126 269 127 
rect 268 127 269 128 
rect 268 138 269 139 
rect 268 139 269 140 
rect 268 140 269 141 
rect 268 141 269 142 
rect 268 142 269 143 
rect 268 143 269 144 
rect 268 154 269 155 
rect 268 155 269 156 
rect 268 156 269 157 
rect 268 157 269 158 
rect 268 158 269 159 
rect 268 159 269 160 
rect 268 170 269 171 
rect 268 171 269 172 
rect 268 172 269 173 
rect 268 173 269 174 
rect 268 174 269 175 
rect 268 175 269 176 
rect 268 186 269 187 
rect 268 187 269 188 
rect 268 188 269 189 
rect 268 189 269 190 
rect 268 190 269 191 
rect 268 191 269 192 
rect 268 202 269 203 
rect 268 203 269 204 
rect 268 204 269 205 
rect 268 205 269 206 
rect 268 206 269 207 
rect 268 207 269 208 
rect 268 218 269 219 
rect 268 219 269 220 
rect 268 220 269 221 
rect 268 221 269 222 
rect 268 222 269 223 
rect 268 223 269 224 
rect 268 234 269 235 
rect 268 235 269 236 
rect 268 236 269 237 
rect 268 237 269 238 
rect 268 238 269 239 
rect 268 239 269 240 
rect 268 250 269 251 
rect 268 251 269 252 
rect 268 252 269 253 
rect 268 253 269 254 
rect 268 254 269 255 
rect 268 255 269 256 
rect 268 266 269 267 
rect 268 267 269 268 
rect 268 268 269 269 
rect 268 269 269 270 
rect 268 270 269 271 
rect 268 271 269 272 
rect 268 282 269 283 
rect 268 283 269 284 
rect 268 284 269 285 
rect 268 285 269 286 
rect 268 286 269 287 
rect 268 287 269 288 
rect 268 298 269 299 
rect 268 299 269 300 
rect 268 300 269 301 
rect 268 301 269 302 
rect 268 302 269 303 
rect 268 303 269 304 
rect 269 10 270 11 
rect 269 11 270 12 
rect 269 12 270 13 
rect 269 13 270 14 
rect 269 14 270 15 
rect 269 15 270 16 
rect 269 26 270 27 
rect 269 27 270 28 
rect 269 28 270 29 
rect 269 29 270 30 
rect 269 30 270 31 
rect 269 31 270 32 
rect 269 42 270 43 
rect 269 43 270 44 
rect 269 44 270 45 
rect 269 45 270 46 
rect 269 46 270 47 
rect 269 47 270 48 
rect 269 58 270 59 
rect 269 59 270 60 
rect 269 60 270 61 
rect 269 61 270 62 
rect 269 62 270 63 
rect 269 63 270 64 
rect 269 74 270 75 
rect 269 75 270 76 
rect 269 76 270 77 
rect 269 77 270 78 
rect 269 78 270 79 
rect 269 79 270 80 
rect 269 90 270 91 
rect 269 91 270 92 
rect 269 92 270 93 
rect 269 93 270 94 
rect 269 94 270 95 
rect 269 95 270 96 
rect 269 106 270 107 
rect 269 107 270 108 
rect 269 108 270 109 
rect 269 109 270 110 
rect 269 110 270 111 
rect 269 111 270 112 
rect 269 122 270 123 
rect 269 123 270 124 
rect 269 124 270 125 
rect 269 125 270 126 
rect 269 126 270 127 
rect 269 127 270 128 
rect 269 138 270 139 
rect 269 139 270 140 
rect 269 140 270 141 
rect 269 141 270 142 
rect 269 142 270 143 
rect 269 143 270 144 
rect 269 154 270 155 
rect 269 155 270 156 
rect 269 156 270 157 
rect 269 157 270 158 
rect 269 158 270 159 
rect 269 159 270 160 
rect 269 170 270 171 
rect 269 171 270 172 
rect 269 172 270 173 
rect 269 173 270 174 
rect 269 174 270 175 
rect 269 175 270 176 
rect 269 186 270 187 
rect 269 187 270 188 
rect 269 188 270 189 
rect 269 189 270 190 
rect 269 190 270 191 
rect 269 191 270 192 
rect 269 202 270 203 
rect 269 203 270 204 
rect 269 204 270 205 
rect 269 205 270 206 
rect 269 206 270 207 
rect 269 207 270 208 
rect 269 218 270 219 
rect 269 219 270 220 
rect 269 220 270 221 
rect 269 221 270 222 
rect 269 222 270 223 
rect 269 223 270 224 
rect 269 234 270 235 
rect 269 235 270 236 
rect 269 236 270 237 
rect 269 237 270 238 
rect 269 238 270 239 
rect 269 239 270 240 
rect 269 250 270 251 
rect 269 251 270 252 
rect 269 252 270 253 
rect 269 253 270 254 
rect 269 254 270 255 
rect 269 255 270 256 
rect 269 266 270 267 
rect 269 267 270 268 
rect 269 268 270 269 
rect 269 269 270 270 
rect 269 270 270 271 
rect 269 271 270 272 
rect 269 282 270 283 
rect 269 283 270 284 
rect 269 284 270 285 
rect 269 285 270 286 
rect 269 286 270 287 
rect 269 287 270 288 
rect 269 298 270 299 
rect 269 299 270 300 
rect 269 300 270 301 
rect 269 301 270 302 
rect 269 302 270 303 
rect 269 303 270 304 
rect 270 10 271 11 
rect 270 11 271 12 
rect 270 12 271 13 
rect 270 13 271 14 
rect 270 14 271 15 
rect 270 15 271 16 
rect 270 26 271 27 
rect 270 27 271 28 
rect 270 28 271 29 
rect 270 29 271 30 
rect 270 30 271 31 
rect 270 31 271 32 
rect 270 42 271 43 
rect 270 43 271 44 
rect 270 44 271 45 
rect 270 45 271 46 
rect 270 46 271 47 
rect 270 47 271 48 
rect 270 58 271 59 
rect 270 59 271 60 
rect 270 60 271 61 
rect 270 61 271 62 
rect 270 62 271 63 
rect 270 63 271 64 
rect 270 74 271 75 
rect 270 75 271 76 
rect 270 76 271 77 
rect 270 77 271 78 
rect 270 78 271 79 
rect 270 79 271 80 
rect 270 90 271 91 
rect 270 91 271 92 
rect 270 92 271 93 
rect 270 93 271 94 
rect 270 94 271 95 
rect 270 95 271 96 
rect 270 106 271 107 
rect 270 107 271 108 
rect 270 108 271 109 
rect 270 109 271 110 
rect 270 110 271 111 
rect 270 111 271 112 
rect 270 122 271 123 
rect 270 123 271 124 
rect 270 124 271 125 
rect 270 125 271 126 
rect 270 126 271 127 
rect 270 127 271 128 
rect 270 138 271 139 
rect 270 139 271 140 
rect 270 140 271 141 
rect 270 141 271 142 
rect 270 142 271 143 
rect 270 143 271 144 
rect 270 154 271 155 
rect 270 155 271 156 
rect 270 156 271 157 
rect 270 157 271 158 
rect 270 158 271 159 
rect 270 159 271 160 
rect 270 170 271 171 
rect 270 171 271 172 
rect 270 172 271 173 
rect 270 173 271 174 
rect 270 174 271 175 
rect 270 175 271 176 
rect 270 186 271 187 
rect 270 187 271 188 
rect 270 188 271 189 
rect 270 189 271 190 
rect 270 190 271 191 
rect 270 191 271 192 
rect 270 202 271 203 
rect 270 203 271 204 
rect 270 204 271 205 
rect 270 205 271 206 
rect 270 206 271 207 
rect 270 207 271 208 
rect 270 218 271 219 
rect 270 219 271 220 
rect 270 220 271 221 
rect 270 221 271 222 
rect 270 222 271 223 
rect 270 223 271 224 
rect 270 234 271 235 
rect 270 235 271 236 
rect 270 236 271 237 
rect 270 237 271 238 
rect 270 238 271 239 
rect 270 239 271 240 
rect 270 250 271 251 
rect 270 251 271 252 
rect 270 252 271 253 
rect 270 253 271 254 
rect 270 254 271 255 
rect 270 255 271 256 
rect 270 266 271 267 
rect 270 267 271 268 
rect 270 268 271 269 
rect 270 269 271 270 
rect 270 270 271 271 
rect 270 271 271 272 
rect 270 282 271 283 
rect 270 283 271 284 
rect 270 284 271 285 
rect 270 285 271 286 
rect 270 286 271 287 
rect 270 287 271 288 
rect 270 298 271 299 
rect 270 299 271 300 
rect 270 300 271 301 
rect 270 301 271 302 
rect 270 302 271 303 
rect 270 303 271 304 
rect 271 10 272 11 
rect 271 11 272 12 
rect 271 12 272 13 
rect 271 13 272 14 
rect 271 14 272 15 
rect 271 15 272 16 
rect 271 26 272 27 
rect 271 27 272 28 
rect 271 28 272 29 
rect 271 29 272 30 
rect 271 31 272 32 
rect 271 42 272 43 
rect 271 43 272 44 
rect 271 44 272 45 
rect 271 45 272 46 
rect 271 46 272 47 
rect 271 47 272 48 
rect 271 58 272 59 
rect 271 59 272 60 
rect 271 60 272 61 
rect 271 61 272 62 
rect 271 62 272 63 
rect 271 63 272 64 
rect 271 74 272 75 
rect 271 76 272 77 
rect 271 77 272 78 
rect 271 78 272 79 
rect 271 79 272 80 
rect 271 90 272 91 
rect 271 91 272 92 
rect 271 92 272 93 
rect 271 93 272 94 
rect 271 94 272 95 
rect 271 95 272 96 
rect 271 106 272 107 
rect 271 108 272 109 
rect 271 109 272 110 
rect 271 111 272 112 
rect 271 122 272 123 
rect 271 123 272 124 
rect 271 124 272 125 
rect 271 125 272 126 
rect 271 127 272 128 
rect 271 138 272 139 
rect 271 139 272 140 
rect 271 140 272 141 
rect 271 141 272 142 
rect 271 143 272 144 
rect 271 154 272 155 
rect 271 155 272 156 
rect 271 156 272 157 
rect 271 157 272 158 
rect 271 159 272 160 
rect 271 170 272 171 
rect 271 172 272 173 
rect 271 173 272 174 
rect 271 175 272 176 
rect 271 186 272 187 
rect 271 188 272 189 
rect 271 189 272 190 
rect 271 190 272 191 
rect 271 191 272 192 
rect 271 202 272 203 
rect 271 203 272 204 
rect 271 204 272 205 
rect 271 205 272 206 
rect 271 207 272 208 
rect 271 218 272 219 
rect 271 220 272 221 
rect 271 221 272 222 
rect 271 223 272 224 
rect 271 234 272 235 
rect 271 236 272 237 
rect 271 237 272 238 
rect 271 238 272 239 
rect 271 239 272 240 
rect 271 250 272 251 
rect 271 251 272 252 
rect 271 252 272 253 
rect 271 253 272 254 
rect 271 255 272 256 
rect 271 266 272 267 
rect 271 267 272 268 
rect 271 268 272 269 
rect 271 269 272 270 
rect 271 270 272 271 
rect 271 271 272 272 
rect 271 282 272 283 
rect 271 284 272 285 
rect 271 285 272 286 
rect 271 286 272 287 
rect 271 287 272 288 
rect 271 298 272 299 
rect 271 299 272 300 
rect 271 300 272 301 
rect 271 301 272 302 
rect 271 302 272 303 
rect 271 303 272 304 
rect 282 10 283 11 
rect 282 11 283 12 
rect 282 12 283 13 
rect 282 13 283 14 
rect 282 15 283 16 
rect 282 26 283 27 
rect 282 27 283 28 
rect 282 28 283 29 
rect 282 29 283 30 
rect 282 30 283 31 
rect 282 31 283 32 
rect 282 42 283 43 
rect 282 43 283 44 
rect 282 44 283 45 
rect 282 45 283 46 
rect 282 46 283 47 
rect 282 47 283 48 
rect 282 58 283 59 
rect 282 59 283 60 
rect 282 60 283 61 
rect 282 61 283 62 
rect 282 63 283 64 
rect 282 74 283 75 
rect 282 76 283 77 
rect 282 77 283 78 
rect 282 78 283 79 
rect 282 79 283 80 
rect 282 90 283 91 
rect 282 91 283 92 
rect 282 92 283 93 
rect 282 93 283 94 
rect 282 95 283 96 
rect 282 106 283 107 
rect 282 108 283 109 
rect 282 109 283 110 
rect 282 110 283 111 
rect 282 111 283 112 
rect 282 122 283 123 
rect 282 124 283 125 
rect 282 125 283 126 
rect 282 126 283 127 
rect 282 127 283 128 
rect 282 138 283 139 
rect 282 140 283 141 
rect 282 141 283 142 
rect 282 143 283 144 
rect 282 154 283 155 
rect 282 155 283 156 
rect 282 156 283 157 
rect 282 157 283 158 
rect 282 159 283 160 
rect 282 170 283 171 
rect 282 172 283 173 
rect 282 173 283 174 
rect 282 175 283 176 
rect 282 186 283 187 
rect 282 187 283 188 
rect 282 188 283 189 
rect 282 189 283 190 
rect 282 190 283 191 
rect 282 191 283 192 
rect 282 202 283 203 
rect 282 204 283 205 
rect 282 205 283 206 
rect 282 207 283 208 
rect 282 218 283 219 
rect 282 220 283 221 
rect 282 221 283 222 
rect 282 222 283 223 
rect 282 223 283 224 
rect 282 234 283 235 
rect 282 236 283 237 
rect 282 237 283 238 
rect 282 238 283 239 
rect 282 239 283 240 
rect 282 250 283 251 
rect 282 251 283 252 
rect 282 252 283 253 
rect 282 253 283 254 
rect 282 255 283 256 
rect 282 266 283 267 
rect 282 267 283 268 
rect 282 268 283 269 
rect 282 269 283 270 
rect 282 271 283 272 
rect 282 282 283 283 
rect 282 283 283 284 
rect 282 284 283 285 
rect 282 285 283 286 
rect 282 287 283 288 
rect 282 298 283 299 
rect 282 299 283 300 
rect 282 300 283 301 
rect 282 301 283 302 
rect 282 303 283 304 
rect 283 10 284 11 
rect 283 11 284 12 
rect 283 12 284 13 
rect 283 13 284 14 
rect 283 14 284 15 
rect 283 15 284 16 
rect 283 26 284 27 
rect 283 27 284 28 
rect 283 28 284 29 
rect 283 29 284 30 
rect 283 30 284 31 
rect 283 31 284 32 
rect 283 42 284 43 
rect 283 43 284 44 
rect 283 44 284 45 
rect 283 45 284 46 
rect 283 46 284 47 
rect 283 47 284 48 
rect 283 58 284 59 
rect 283 59 284 60 
rect 283 60 284 61 
rect 283 61 284 62 
rect 283 62 284 63 
rect 283 63 284 64 
rect 283 74 284 75 
rect 283 75 284 76 
rect 283 76 284 77 
rect 283 77 284 78 
rect 283 78 284 79 
rect 283 79 284 80 
rect 283 90 284 91 
rect 283 91 284 92 
rect 283 92 284 93 
rect 283 93 284 94 
rect 283 94 284 95 
rect 283 95 284 96 
rect 283 106 284 107 
rect 283 107 284 108 
rect 283 108 284 109 
rect 283 109 284 110 
rect 283 110 284 111 
rect 283 111 284 112 
rect 283 122 284 123 
rect 283 123 284 124 
rect 283 124 284 125 
rect 283 125 284 126 
rect 283 126 284 127 
rect 283 127 284 128 
rect 283 138 284 139 
rect 283 139 284 140 
rect 283 140 284 141 
rect 283 141 284 142 
rect 283 142 284 143 
rect 283 143 284 144 
rect 283 154 284 155 
rect 283 155 284 156 
rect 283 156 284 157 
rect 283 157 284 158 
rect 283 158 284 159 
rect 283 159 284 160 
rect 283 170 284 171 
rect 283 171 284 172 
rect 283 172 284 173 
rect 283 173 284 174 
rect 283 174 284 175 
rect 283 175 284 176 
rect 283 186 284 187 
rect 283 187 284 188 
rect 283 188 284 189 
rect 283 189 284 190 
rect 283 190 284 191 
rect 283 191 284 192 
rect 283 202 284 203 
rect 283 203 284 204 
rect 283 204 284 205 
rect 283 205 284 206 
rect 283 206 284 207 
rect 283 207 284 208 
rect 283 218 284 219 
rect 283 219 284 220 
rect 283 220 284 221 
rect 283 221 284 222 
rect 283 222 284 223 
rect 283 223 284 224 
rect 283 234 284 235 
rect 283 235 284 236 
rect 283 236 284 237 
rect 283 237 284 238 
rect 283 238 284 239 
rect 283 239 284 240 
rect 283 250 284 251 
rect 283 251 284 252 
rect 283 252 284 253 
rect 283 253 284 254 
rect 283 254 284 255 
rect 283 255 284 256 
rect 283 266 284 267 
rect 283 267 284 268 
rect 283 268 284 269 
rect 283 269 284 270 
rect 283 270 284 271 
rect 283 271 284 272 
rect 283 282 284 283 
rect 283 283 284 284 
rect 283 284 284 285 
rect 283 285 284 286 
rect 283 286 284 287 
rect 283 287 284 288 
rect 283 298 284 299 
rect 283 299 284 300 
rect 283 300 284 301 
rect 283 301 284 302 
rect 283 302 284 303 
rect 283 303 284 304 
rect 284 10 285 11 
rect 284 11 285 12 
rect 284 12 285 13 
rect 284 13 285 14 
rect 284 14 285 15 
rect 284 15 285 16 
rect 284 26 285 27 
rect 284 27 285 28 
rect 284 28 285 29 
rect 284 29 285 30 
rect 284 30 285 31 
rect 284 31 285 32 
rect 284 42 285 43 
rect 284 43 285 44 
rect 284 44 285 45 
rect 284 45 285 46 
rect 284 46 285 47 
rect 284 47 285 48 
rect 284 58 285 59 
rect 284 59 285 60 
rect 284 60 285 61 
rect 284 61 285 62 
rect 284 62 285 63 
rect 284 63 285 64 
rect 284 74 285 75 
rect 284 75 285 76 
rect 284 76 285 77 
rect 284 77 285 78 
rect 284 78 285 79 
rect 284 79 285 80 
rect 284 90 285 91 
rect 284 91 285 92 
rect 284 92 285 93 
rect 284 93 285 94 
rect 284 94 285 95 
rect 284 95 285 96 
rect 284 106 285 107 
rect 284 107 285 108 
rect 284 108 285 109 
rect 284 109 285 110 
rect 284 110 285 111 
rect 284 111 285 112 
rect 284 122 285 123 
rect 284 123 285 124 
rect 284 124 285 125 
rect 284 125 285 126 
rect 284 126 285 127 
rect 284 127 285 128 
rect 284 138 285 139 
rect 284 139 285 140 
rect 284 140 285 141 
rect 284 141 285 142 
rect 284 142 285 143 
rect 284 143 285 144 
rect 284 154 285 155 
rect 284 155 285 156 
rect 284 156 285 157 
rect 284 157 285 158 
rect 284 158 285 159 
rect 284 159 285 160 
rect 284 170 285 171 
rect 284 171 285 172 
rect 284 172 285 173 
rect 284 173 285 174 
rect 284 174 285 175 
rect 284 175 285 176 
rect 284 186 285 187 
rect 284 187 285 188 
rect 284 188 285 189 
rect 284 189 285 190 
rect 284 190 285 191 
rect 284 191 285 192 
rect 284 202 285 203 
rect 284 203 285 204 
rect 284 204 285 205 
rect 284 205 285 206 
rect 284 206 285 207 
rect 284 207 285 208 
rect 284 218 285 219 
rect 284 219 285 220 
rect 284 220 285 221 
rect 284 221 285 222 
rect 284 222 285 223 
rect 284 223 285 224 
rect 284 234 285 235 
rect 284 235 285 236 
rect 284 236 285 237 
rect 284 237 285 238 
rect 284 238 285 239 
rect 284 239 285 240 
rect 284 250 285 251 
rect 284 251 285 252 
rect 284 252 285 253 
rect 284 253 285 254 
rect 284 254 285 255 
rect 284 255 285 256 
rect 284 266 285 267 
rect 284 267 285 268 
rect 284 268 285 269 
rect 284 269 285 270 
rect 284 270 285 271 
rect 284 271 285 272 
rect 284 282 285 283 
rect 284 283 285 284 
rect 284 284 285 285 
rect 284 285 285 286 
rect 284 286 285 287 
rect 284 287 285 288 
rect 284 298 285 299 
rect 284 299 285 300 
rect 284 300 285 301 
rect 284 301 285 302 
rect 284 302 285 303 
rect 284 303 285 304 
rect 285 10 286 11 
rect 285 11 286 12 
rect 285 12 286 13 
rect 285 13 286 14 
rect 285 14 286 15 
rect 285 15 286 16 
rect 285 26 286 27 
rect 285 27 286 28 
rect 285 28 286 29 
rect 285 29 286 30 
rect 285 30 286 31 
rect 285 31 286 32 
rect 285 42 286 43 
rect 285 43 286 44 
rect 285 44 286 45 
rect 285 45 286 46 
rect 285 46 286 47 
rect 285 47 286 48 
rect 285 58 286 59 
rect 285 59 286 60 
rect 285 60 286 61 
rect 285 61 286 62 
rect 285 62 286 63 
rect 285 63 286 64 
rect 285 74 286 75 
rect 285 75 286 76 
rect 285 76 286 77 
rect 285 77 286 78 
rect 285 78 286 79 
rect 285 79 286 80 
rect 285 90 286 91 
rect 285 91 286 92 
rect 285 92 286 93 
rect 285 93 286 94 
rect 285 94 286 95 
rect 285 95 286 96 
rect 285 106 286 107 
rect 285 107 286 108 
rect 285 108 286 109 
rect 285 109 286 110 
rect 285 110 286 111 
rect 285 111 286 112 
rect 285 122 286 123 
rect 285 123 286 124 
rect 285 124 286 125 
rect 285 125 286 126 
rect 285 126 286 127 
rect 285 127 286 128 
rect 285 138 286 139 
rect 285 139 286 140 
rect 285 140 286 141 
rect 285 141 286 142 
rect 285 142 286 143 
rect 285 143 286 144 
rect 285 154 286 155 
rect 285 155 286 156 
rect 285 156 286 157 
rect 285 157 286 158 
rect 285 158 286 159 
rect 285 159 286 160 
rect 285 170 286 171 
rect 285 171 286 172 
rect 285 172 286 173 
rect 285 173 286 174 
rect 285 174 286 175 
rect 285 175 286 176 
rect 285 186 286 187 
rect 285 187 286 188 
rect 285 188 286 189 
rect 285 189 286 190 
rect 285 190 286 191 
rect 285 191 286 192 
rect 285 202 286 203 
rect 285 203 286 204 
rect 285 204 286 205 
rect 285 205 286 206 
rect 285 206 286 207 
rect 285 207 286 208 
rect 285 218 286 219 
rect 285 219 286 220 
rect 285 220 286 221 
rect 285 221 286 222 
rect 285 222 286 223 
rect 285 223 286 224 
rect 285 234 286 235 
rect 285 235 286 236 
rect 285 236 286 237 
rect 285 237 286 238 
rect 285 238 286 239 
rect 285 239 286 240 
rect 285 250 286 251 
rect 285 251 286 252 
rect 285 252 286 253 
rect 285 253 286 254 
rect 285 254 286 255 
rect 285 255 286 256 
rect 285 266 286 267 
rect 285 267 286 268 
rect 285 268 286 269 
rect 285 269 286 270 
rect 285 270 286 271 
rect 285 271 286 272 
rect 285 282 286 283 
rect 285 283 286 284 
rect 285 284 286 285 
rect 285 285 286 286 
rect 285 286 286 287 
rect 285 287 286 288 
rect 285 298 286 299 
rect 285 299 286 300 
rect 285 300 286 301 
rect 285 301 286 302 
rect 285 302 286 303 
rect 285 303 286 304 
rect 286 10 287 11 
rect 286 11 287 12 
rect 286 12 287 13 
rect 286 13 287 14 
rect 286 14 287 15 
rect 286 15 287 16 
rect 286 26 287 27 
rect 286 27 287 28 
rect 286 28 287 29 
rect 286 29 287 30 
rect 286 30 287 31 
rect 286 31 287 32 
rect 286 42 287 43 
rect 286 43 287 44 
rect 286 44 287 45 
rect 286 45 287 46 
rect 286 46 287 47 
rect 286 47 287 48 
rect 286 58 287 59 
rect 286 59 287 60 
rect 286 60 287 61 
rect 286 61 287 62 
rect 286 62 287 63 
rect 286 63 287 64 
rect 286 74 287 75 
rect 286 75 287 76 
rect 286 76 287 77 
rect 286 77 287 78 
rect 286 78 287 79 
rect 286 79 287 80 
rect 286 90 287 91 
rect 286 91 287 92 
rect 286 92 287 93 
rect 286 93 287 94 
rect 286 94 287 95 
rect 286 95 287 96 
rect 286 106 287 107 
rect 286 107 287 108 
rect 286 108 287 109 
rect 286 109 287 110 
rect 286 110 287 111 
rect 286 111 287 112 
rect 286 122 287 123 
rect 286 123 287 124 
rect 286 124 287 125 
rect 286 125 287 126 
rect 286 126 287 127 
rect 286 127 287 128 
rect 286 138 287 139 
rect 286 139 287 140 
rect 286 140 287 141 
rect 286 141 287 142 
rect 286 142 287 143 
rect 286 143 287 144 
rect 286 154 287 155 
rect 286 155 287 156 
rect 286 156 287 157 
rect 286 157 287 158 
rect 286 158 287 159 
rect 286 159 287 160 
rect 286 170 287 171 
rect 286 171 287 172 
rect 286 172 287 173 
rect 286 173 287 174 
rect 286 174 287 175 
rect 286 175 287 176 
rect 286 186 287 187 
rect 286 187 287 188 
rect 286 188 287 189 
rect 286 189 287 190 
rect 286 190 287 191 
rect 286 191 287 192 
rect 286 202 287 203 
rect 286 203 287 204 
rect 286 204 287 205 
rect 286 205 287 206 
rect 286 206 287 207 
rect 286 207 287 208 
rect 286 218 287 219 
rect 286 219 287 220 
rect 286 220 287 221 
rect 286 221 287 222 
rect 286 222 287 223 
rect 286 223 287 224 
rect 286 234 287 235 
rect 286 235 287 236 
rect 286 236 287 237 
rect 286 237 287 238 
rect 286 238 287 239 
rect 286 239 287 240 
rect 286 250 287 251 
rect 286 251 287 252 
rect 286 252 287 253 
rect 286 253 287 254 
rect 286 254 287 255 
rect 286 255 287 256 
rect 286 266 287 267 
rect 286 267 287 268 
rect 286 268 287 269 
rect 286 269 287 270 
rect 286 270 287 271 
rect 286 271 287 272 
rect 286 282 287 283 
rect 286 283 287 284 
rect 286 284 287 285 
rect 286 285 287 286 
rect 286 286 287 287 
rect 286 287 287 288 
rect 286 298 287 299 
rect 286 299 287 300 
rect 286 300 287 301 
rect 286 301 287 302 
rect 286 302 287 303 
rect 286 303 287 304 
rect 287 10 288 11 
rect 287 11 288 12 
rect 287 12 288 13 
rect 287 13 288 14 
rect 287 15 288 16 
rect 287 26 288 27 
rect 287 27 288 28 
rect 287 28 288 29 
rect 287 29 288 30 
rect 287 31 288 32 
rect 287 42 288 43 
rect 287 44 288 45 
rect 287 45 288 46 
rect 287 47 288 48 
rect 287 58 288 59 
rect 287 59 288 60 
rect 287 60 288 61 
rect 287 61 288 62 
rect 287 63 288 64 
rect 287 74 288 75 
rect 287 75 288 76 
rect 287 76 288 77 
rect 287 77 288 78 
rect 287 78 288 79 
rect 287 79 288 80 
rect 287 90 288 91 
rect 287 92 288 93 
rect 287 93 288 94 
rect 287 94 288 95 
rect 287 95 288 96 
rect 287 106 288 107 
rect 287 107 288 108 
rect 287 108 288 109 
rect 287 109 288 110 
rect 287 111 288 112 
rect 287 122 288 123 
rect 287 123 288 124 
rect 287 124 288 125 
rect 287 125 288 126 
rect 287 127 288 128 
rect 287 138 288 139 
rect 287 140 288 141 
rect 287 141 288 142 
rect 287 143 288 144 
rect 287 154 288 155 
rect 287 156 288 157 
rect 287 157 288 158 
rect 287 159 288 160 
rect 287 170 288 171 
rect 287 172 288 173 
rect 287 173 288 174 
rect 287 174 288 175 
rect 287 175 288 176 
rect 287 186 288 187 
rect 287 187 288 188 
rect 287 188 288 189 
rect 287 189 288 190 
rect 287 190 288 191 
rect 287 191 288 192 
rect 287 202 288 203 
rect 287 204 288 205 
rect 287 205 288 206 
rect 287 206 288 207 
rect 287 207 288 208 
rect 287 218 288 219 
rect 287 219 288 220 
rect 287 220 288 221 
rect 287 221 288 222 
rect 287 222 288 223 
rect 287 223 288 224 
rect 287 234 288 235 
rect 287 235 288 236 
rect 287 236 288 237 
rect 287 237 288 238 
rect 287 239 288 240 
rect 287 250 288 251 
rect 287 252 288 253 
rect 287 253 288 254 
rect 287 254 288 255 
rect 287 255 288 256 
rect 287 266 288 267 
rect 287 268 288 269 
rect 287 269 288 270 
rect 287 270 288 271 
rect 287 271 288 272 
rect 287 282 288 283 
rect 287 284 288 285 
rect 287 285 288 286 
rect 287 286 288 287 
rect 287 287 288 288 
rect 287 298 288 299 
rect 287 300 288 301 
rect 287 301 288 302 
rect 287 302 288 303 
rect 287 303 288 304 
rect 298 10 299 11 
rect 298 12 299 13 
rect 298 13 299 14 
rect 298 15 299 16 
rect 298 26 299 27 
rect 298 28 299 29 
rect 298 29 299 30 
rect 298 31 299 32 
rect 298 42 299 43 
rect 298 44 299 45 
rect 298 45 299 46 
rect 298 46 299 47 
rect 298 47 299 48 
rect 298 58 299 59 
rect 298 60 299 61 
rect 298 61 299 62 
rect 298 63 299 64 
rect 298 74 299 75 
rect 298 75 299 76 
rect 298 76 299 77 
rect 298 77 299 78 
rect 298 79 299 80 
rect 298 90 299 91 
rect 298 92 299 93 
rect 298 93 299 94 
rect 298 94 299 95 
rect 298 95 299 96 
rect 298 106 299 107 
rect 298 108 299 109 
rect 298 109 299 110 
rect 298 111 299 112 
rect 298 122 299 123 
rect 298 124 299 125 
rect 298 125 299 126 
rect 298 126 299 127 
rect 298 127 299 128 
rect 298 138 299 139 
rect 298 139 299 140 
rect 298 140 299 141 
rect 298 141 299 142 
rect 298 143 299 144 
rect 298 154 299 155 
rect 298 156 299 157 
rect 298 157 299 158 
rect 298 159 299 160 
rect 298 170 299 171 
rect 298 172 299 173 
rect 298 173 299 174 
rect 298 174 299 175 
rect 298 175 299 176 
rect 298 186 299 187 
rect 298 187 299 188 
rect 298 188 299 189 
rect 298 189 299 190 
rect 298 190 299 191 
rect 298 191 299 192 
rect 298 202 299 203 
rect 298 204 299 205 
rect 298 205 299 206 
rect 298 206 299 207 
rect 298 207 299 208 
rect 298 218 299 219 
rect 298 219 299 220 
rect 298 220 299 221 
rect 298 221 299 222 
rect 298 222 299 223 
rect 298 223 299 224 
rect 298 234 299 235 
rect 298 236 299 237 
rect 298 237 299 238 
rect 298 239 299 240 
rect 298 250 299 251 
rect 298 251 299 252 
rect 298 252 299 253 
rect 298 253 299 254 
rect 298 255 299 256 
rect 298 266 299 267 
rect 298 268 299 269 
rect 298 269 299 270 
rect 298 271 299 272 
rect 298 282 299 283 
rect 298 284 299 285 
rect 298 285 299 286 
rect 298 286 299 287 
rect 298 287 299 288 
rect 298 298 299 299 
rect 298 299 299 300 
rect 298 300 299 301 
rect 298 301 299 302 
rect 298 303 299 304 
rect 299 10 300 11 
rect 299 11 300 12 
rect 299 12 300 13 
rect 299 13 300 14 
rect 299 14 300 15 
rect 299 15 300 16 
rect 299 26 300 27 
rect 299 27 300 28 
rect 299 28 300 29 
rect 299 29 300 30 
rect 299 30 300 31 
rect 299 31 300 32 
rect 299 42 300 43 
rect 299 43 300 44 
rect 299 44 300 45 
rect 299 45 300 46 
rect 299 46 300 47 
rect 299 47 300 48 
rect 299 58 300 59 
rect 299 59 300 60 
rect 299 60 300 61 
rect 299 61 300 62 
rect 299 62 300 63 
rect 299 63 300 64 
rect 299 74 300 75 
rect 299 75 300 76 
rect 299 76 300 77 
rect 299 77 300 78 
rect 299 78 300 79 
rect 299 79 300 80 
rect 299 90 300 91 
rect 299 91 300 92 
rect 299 92 300 93 
rect 299 93 300 94 
rect 299 94 300 95 
rect 299 95 300 96 
rect 299 106 300 107 
rect 299 107 300 108 
rect 299 108 300 109 
rect 299 109 300 110 
rect 299 110 300 111 
rect 299 111 300 112 
rect 299 122 300 123 
rect 299 123 300 124 
rect 299 124 300 125 
rect 299 125 300 126 
rect 299 126 300 127 
rect 299 127 300 128 
rect 299 138 300 139 
rect 299 139 300 140 
rect 299 140 300 141 
rect 299 141 300 142 
rect 299 142 300 143 
rect 299 143 300 144 
rect 299 154 300 155 
rect 299 155 300 156 
rect 299 156 300 157 
rect 299 157 300 158 
rect 299 158 300 159 
rect 299 159 300 160 
rect 299 170 300 171 
rect 299 171 300 172 
rect 299 172 300 173 
rect 299 173 300 174 
rect 299 174 300 175 
rect 299 175 300 176 
rect 299 186 300 187 
rect 299 187 300 188 
rect 299 188 300 189 
rect 299 189 300 190 
rect 299 190 300 191 
rect 299 191 300 192 
rect 299 202 300 203 
rect 299 203 300 204 
rect 299 204 300 205 
rect 299 205 300 206 
rect 299 206 300 207 
rect 299 207 300 208 
rect 299 218 300 219 
rect 299 219 300 220 
rect 299 220 300 221 
rect 299 221 300 222 
rect 299 222 300 223 
rect 299 223 300 224 
rect 299 234 300 235 
rect 299 235 300 236 
rect 299 236 300 237 
rect 299 237 300 238 
rect 299 238 300 239 
rect 299 239 300 240 
rect 299 250 300 251 
rect 299 251 300 252 
rect 299 252 300 253 
rect 299 253 300 254 
rect 299 254 300 255 
rect 299 255 300 256 
rect 299 266 300 267 
rect 299 267 300 268 
rect 299 268 300 269 
rect 299 269 300 270 
rect 299 270 300 271 
rect 299 271 300 272 
rect 299 282 300 283 
rect 299 283 300 284 
rect 299 284 300 285 
rect 299 285 300 286 
rect 299 286 300 287 
rect 299 287 300 288 
rect 299 298 300 299 
rect 299 299 300 300 
rect 299 300 300 301 
rect 299 301 300 302 
rect 299 302 300 303 
rect 299 303 300 304 
rect 300 10 301 11 
rect 300 11 301 12 
rect 300 12 301 13 
rect 300 13 301 14 
rect 300 14 301 15 
rect 300 15 301 16 
rect 300 26 301 27 
rect 300 27 301 28 
rect 300 28 301 29 
rect 300 29 301 30 
rect 300 30 301 31 
rect 300 31 301 32 
rect 300 42 301 43 
rect 300 43 301 44 
rect 300 44 301 45 
rect 300 45 301 46 
rect 300 46 301 47 
rect 300 47 301 48 
rect 300 58 301 59 
rect 300 59 301 60 
rect 300 60 301 61 
rect 300 61 301 62 
rect 300 62 301 63 
rect 300 63 301 64 
rect 300 74 301 75 
rect 300 75 301 76 
rect 300 76 301 77 
rect 300 77 301 78 
rect 300 78 301 79 
rect 300 79 301 80 
rect 300 90 301 91 
rect 300 91 301 92 
rect 300 92 301 93 
rect 300 93 301 94 
rect 300 94 301 95 
rect 300 95 301 96 
rect 300 106 301 107 
rect 300 107 301 108 
rect 300 108 301 109 
rect 300 109 301 110 
rect 300 110 301 111 
rect 300 111 301 112 
rect 300 122 301 123 
rect 300 123 301 124 
rect 300 124 301 125 
rect 300 125 301 126 
rect 300 126 301 127 
rect 300 127 301 128 
rect 300 138 301 139 
rect 300 139 301 140 
rect 300 140 301 141 
rect 300 141 301 142 
rect 300 142 301 143 
rect 300 143 301 144 
rect 300 154 301 155 
rect 300 155 301 156 
rect 300 156 301 157 
rect 300 157 301 158 
rect 300 158 301 159 
rect 300 159 301 160 
rect 300 170 301 171 
rect 300 171 301 172 
rect 300 172 301 173 
rect 300 173 301 174 
rect 300 174 301 175 
rect 300 175 301 176 
rect 300 186 301 187 
rect 300 187 301 188 
rect 300 188 301 189 
rect 300 189 301 190 
rect 300 190 301 191 
rect 300 191 301 192 
rect 300 202 301 203 
rect 300 203 301 204 
rect 300 204 301 205 
rect 300 205 301 206 
rect 300 206 301 207 
rect 300 207 301 208 
rect 300 218 301 219 
rect 300 219 301 220 
rect 300 220 301 221 
rect 300 221 301 222 
rect 300 222 301 223 
rect 300 223 301 224 
rect 300 234 301 235 
rect 300 235 301 236 
rect 300 236 301 237 
rect 300 237 301 238 
rect 300 238 301 239 
rect 300 239 301 240 
rect 300 250 301 251 
rect 300 251 301 252 
rect 300 252 301 253 
rect 300 253 301 254 
rect 300 254 301 255 
rect 300 255 301 256 
rect 300 266 301 267 
rect 300 267 301 268 
rect 300 268 301 269 
rect 300 269 301 270 
rect 300 270 301 271 
rect 300 271 301 272 
rect 300 282 301 283 
rect 300 283 301 284 
rect 300 284 301 285 
rect 300 285 301 286 
rect 300 286 301 287 
rect 300 287 301 288 
rect 300 298 301 299 
rect 300 299 301 300 
rect 300 300 301 301 
rect 300 301 301 302 
rect 300 302 301 303 
rect 300 303 301 304 
rect 301 10 302 11 
rect 301 11 302 12 
rect 301 12 302 13 
rect 301 13 302 14 
rect 301 14 302 15 
rect 301 15 302 16 
rect 301 26 302 27 
rect 301 27 302 28 
rect 301 28 302 29 
rect 301 29 302 30 
rect 301 30 302 31 
rect 301 31 302 32 
rect 301 42 302 43 
rect 301 43 302 44 
rect 301 44 302 45 
rect 301 45 302 46 
rect 301 46 302 47 
rect 301 47 302 48 
rect 301 58 302 59 
rect 301 59 302 60 
rect 301 60 302 61 
rect 301 61 302 62 
rect 301 62 302 63 
rect 301 63 302 64 
rect 301 74 302 75 
rect 301 75 302 76 
rect 301 76 302 77 
rect 301 77 302 78 
rect 301 78 302 79 
rect 301 79 302 80 
rect 301 90 302 91 
rect 301 91 302 92 
rect 301 92 302 93 
rect 301 93 302 94 
rect 301 94 302 95 
rect 301 95 302 96 
rect 301 106 302 107 
rect 301 107 302 108 
rect 301 108 302 109 
rect 301 109 302 110 
rect 301 110 302 111 
rect 301 111 302 112 
rect 301 122 302 123 
rect 301 123 302 124 
rect 301 124 302 125 
rect 301 125 302 126 
rect 301 126 302 127 
rect 301 127 302 128 
rect 301 138 302 139 
rect 301 139 302 140 
rect 301 140 302 141 
rect 301 141 302 142 
rect 301 142 302 143 
rect 301 143 302 144 
rect 301 154 302 155 
rect 301 155 302 156 
rect 301 156 302 157 
rect 301 157 302 158 
rect 301 158 302 159 
rect 301 159 302 160 
rect 301 170 302 171 
rect 301 171 302 172 
rect 301 172 302 173 
rect 301 173 302 174 
rect 301 174 302 175 
rect 301 175 302 176 
rect 301 186 302 187 
rect 301 187 302 188 
rect 301 188 302 189 
rect 301 189 302 190 
rect 301 190 302 191 
rect 301 191 302 192 
rect 301 202 302 203 
rect 301 203 302 204 
rect 301 204 302 205 
rect 301 205 302 206 
rect 301 206 302 207 
rect 301 207 302 208 
rect 301 218 302 219 
rect 301 219 302 220 
rect 301 220 302 221 
rect 301 221 302 222 
rect 301 222 302 223 
rect 301 223 302 224 
rect 301 234 302 235 
rect 301 235 302 236 
rect 301 236 302 237 
rect 301 237 302 238 
rect 301 238 302 239 
rect 301 239 302 240 
rect 301 250 302 251 
rect 301 251 302 252 
rect 301 252 302 253 
rect 301 253 302 254 
rect 301 254 302 255 
rect 301 255 302 256 
rect 301 266 302 267 
rect 301 267 302 268 
rect 301 268 302 269 
rect 301 269 302 270 
rect 301 270 302 271 
rect 301 271 302 272 
rect 301 282 302 283 
rect 301 283 302 284 
rect 301 284 302 285 
rect 301 285 302 286 
rect 301 286 302 287 
rect 301 287 302 288 
rect 301 298 302 299 
rect 301 299 302 300 
rect 301 300 302 301 
rect 301 301 302 302 
rect 301 302 302 303 
rect 301 303 302 304 
rect 302 10 303 11 
rect 302 11 303 12 
rect 302 12 303 13 
rect 302 13 303 14 
rect 302 14 303 15 
rect 302 15 303 16 
rect 302 26 303 27 
rect 302 27 303 28 
rect 302 28 303 29 
rect 302 29 303 30 
rect 302 30 303 31 
rect 302 31 303 32 
rect 302 42 303 43 
rect 302 43 303 44 
rect 302 44 303 45 
rect 302 45 303 46 
rect 302 46 303 47 
rect 302 47 303 48 
rect 302 58 303 59 
rect 302 59 303 60 
rect 302 60 303 61 
rect 302 61 303 62 
rect 302 62 303 63 
rect 302 63 303 64 
rect 302 74 303 75 
rect 302 75 303 76 
rect 302 76 303 77 
rect 302 77 303 78 
rect 302 78 303 79 
rect 302 79 303 80 
rect 302 90 303 91 
rect 302 91 303 92 
rect 302 92 303 93 
rect 302 93 303 94 
rect 302 94 303 95 
rect 302 95 303 96 
rect 302 106 303 107 
rect 302 107 303 108 
rect 302 108 303 109 
rect 302 109 303 110 
rect 302 110 303 111 
rect 302 111 303 112 
rect 302 122 303 123 
rect 302 123 303 124 
rect 302 124 303 125 
rect 302 125 303 126 
rect 302 126 303 127 
rect 302 127 303 128 
rect 302 138 303 139 
rect 302 139 303 140 
rect 302 140 303 141 
rect 302 141 303 142 
rect 302 142 303 143 
rect 302 143 303 144 
rect 302 154 303 155 
rect 302 155 303 156 
rect 302 156 303 157 
rect 302 157 303 158 
rect 302 158 303 159 
rect 302 159 303 160 
rect 302 170 303 171 
rect 302 171 303 172 
rect 302 172 303 173 
rect 302 173 303 174 
rect 302 174 303 175 
rect 302 175 303 176 
rect 302 186 303 187 
rect 302 187 303 188 
rect 302 188 303 189 
rect 302 189 303 190 
rect 302 190 303 191 
rect 302 191 303 192 
rect 302 202 303 203 
rect 302 203 303 204 
rect 302 204 303 205 
rect 302 205 303 206 
rect 302 206 303 207 
rect 302 207 303 208 
rect 302 218 303 219 
rect 302 219 303 220 
rect 302 220 303 221 
rect 302 221 303 222 
rect 302 222 303 223 
rect 302 223 303 224 
rect 302 234 303 235 
rect 302 235 303 236 
rect 302 236 303 237 
rect 302 237 303 238 
rect 302 238 303 239 
rect 302 239 303 240 
rect 302 250 303 251 
rect 302 251 303 252 
rect 302 252 303 253 
rect 302 253 303 254 
rect 302 254 303 255 
rect 302 255 303 256 
rect 302 266 303 267 
rect 302 267 303 268 
rect 302 268 303 269 
rect 302 269 303 270 
rect 302 270 303 271 
rect 302 271 303 272 
rect 302 282 303 283 
rect 302 283 303 284 
rect 302 284 303 285 
rect 302 285 303 286 
rect 302 286 303 287 
rect 302 287 303 288 
rect 302 298 303 299 
rect 302 299 303 300 
rect 302 300 303 301 
rect 302 301 303 302 
rect 302 302 303 303 
rect 302 303 303 304 
rect 303 10 304 11 
rect 303 12 304 13 
rect 303 13 304 14 
rect 303 14 304 15 
rect 303 15 304 16 
rect 303 26 304 27 
rect 303 28 304 29 
rect 303 29 304 30 
rect 303 31 304 32 
rect 303 42 304 43 
rect 303 44 304 45 
rect 303 45 304 46 
rect 303 47 304 48 
rect 303 58 304 59 
rect 303 59 304 60 
rect 303 60 304 61 
rect 303 61 304 62 
rect 303 62 304 63 
rect 303 63 304 64 
rect 303 74 304 75 
rect 303 76 304 77 
rect 303 77 304 78 
rect 303 79 304 80 
rect 303 90 304 91 
rect 303 91 304 92 
rect 303 92 304 93 
rect 303 93 304 94 
rect 303 95 304 96 
rect 303 106 304 107 
rect 303 107 304 108 
rect 303 108 304 109 
rect 303 109 304 110 
rect 303 111 304 112 
rect 303 122 304 123 
rect 303 124 304 125 
rect 303 125 304 126 
rect 303 126 304 127 
rect 303 127 304 128 
rect 303 138 304 139 
rect 303 140 304 141 
rect 303 141 304 142 
rect 303 142 304 143 
rect 303 143 304 144 
rect 303 154 304 155 
rect 303 156 304 157 
rect 303 157 304 158 
rect 303 159 304 160 
rect 303 170 304 171 
rect 303 171 304 172 
rect 303 172 304 173 
rect 303 173 304 174 
rect 303 175 304 176 
rect 303 186 304 187 
rect 303 187 304 188 
rect 303 188 304 189 
rect 303 189 304 190 
rect 303 190 304 191 
rect 303 191 304 192 
rect 303 202 304 203 
rect 303 203 304 204 
rect 303 204 304 205 
rect 303 205 304 206 
rect 303 206 304 207 
rect 303 207 304 208 
rect 303 218 304 219 
rect 303 220 304 221 
rect 303 221 304 222 
rect 303 222 304 223 
rect 303 223 304 224 
rect 303 234 304 235 
rect 303 235 304 236 
rect 303 236 304 237 
rect 303 237 304 238 
rect 303 238 304 239 
rect 303 239 304 240 
rect 303 250 304 251 
rect 303 251 304 252 
rect 303 252 304 253 
rect 303 253 304 254 
rect 303 254 304 255 
rect 303 255 304 256 
rect 303 266 304 267 
rect 303 268 304 269 
rect 303 269 304 270 
rect 303 271 304 272 
rect 303 282 304 283 
rect 303 283 304 284 
rect 303 284 304 285 
rect 303 285 304 286 
rect 303 287 304 288 
rect 303 298 304 299 
rect 303 299 304 300 
rect 303 300 304 301 
rect 303 301 304 302 
rect 303 302 304 303 
rect 303 303 304 304 
<< labels >>
<< metal1 >>
rect 1 127 2 128 
rect 1 128 2 129 
rect 1 129 2 130 
rect 1 130 2 131 
rect 1 131 2 132 
rect 1 132 2 133 
rect 1 133 2 134 
rect 2 118 3 119 
rect 2 119 3 120 
rect 2 120 3 121 
rect 2 121 3 122 
rect 2 122 3 123 
rect 2 123 3 124 
rect 2 124 3 125 
rect 2 125 3 126 
rect 2 126 3 127 
rect 2 127 3 128 
rect 2 133 3 134 
rect 3 56 4 57 
rect 3 57 4 58 
rect 3 58 4 59 
rect 3 59 4 60 
rect 3 60 4 61 
rect 3 61 4 62 
rect 3 62 4 63 
rect 3 63 4 64 
rect 3 64 4 65 
rect 3 65 4 66 
rect 3 66 4 67 
rect 3 67 4 68 
rect 3 68 4 69 
rect 3 69 4 70 
rect 3 70 4 71 
rect 3 71 4 72 
rect 3 72 4 73 
rect 3 73 4 74 
rect 3 74 4 75 
rect 3 75 4 76 
rect 3 76 4 77 
rect 3 77 4 78 
rect 3 78 4 79 
rect 3 79 4 80 
rect 3 80 4 81 
rect 3 81 4 82 
rect 3 82 4 83 
rect 3 83 4 84 
rect 3 84 4 85 
rect 3 85 4 86 
rect 3 86 4 87 
rect 3 87 4 88 
rect 3 88 4 89 
rect 3 89 4 90 
rect 3 90 4 91 
rect 3 91 4 92 
rect 3 92 4 93 
rect 3 93 4 94 
rect 3 94 4 95 
rect 3 95 4 96 
rect 3 96 4 97 
rect 3 97 4 98 
rect 3 98 4 99 
rect 3 99 4 100 
rect 3 100 4 101 
rect 3 101 4 102 
rect 3 102 4 103 
rect 3 103 4 104 
rect 3 104 4 105 
rect 3 105 4 106 
rect 3 106 4 107 
rect 3 107 4 108 
rect 3 108 4 109 
rect 3 109 4 110 
rect 3 110 4 111 
rect 3 111 4 112 
rect 3 112 4 113 
rect 3 113 4 114 
rect 3 114 4 115 
rect 3 115 4 116 
rect 3 116 4 117 
rect 3 117 4 118 
rect 3 118 4 119 
rect 3 135 4 136 
rect 3 136 4 137 
rect 3 137 4 138 
rect 3 138 4 139 
rect 3 139 4 140 
rect 3 140 4 141 
rect 3 141 4 142 
rect 3 142 4 143 
rect 3 143 4 144 
rect 3 144 4 145 
rect 3 145 4 146 
rect 3 146 4 147 
rect 3 147 4 148 
rect 3 148 4 149 
rect 3 149 4 150 
rect 3 150 4 151 
rect 3 151 4 152 
rect 3 152 4 153 
rect 3 153 4 154 
rect 3 154 4 155 
rect 3 155 4 156 
rect 3 156 4 157 
rect 3 157 4 158 
rect 3 158 4 159 
rect 3 159 4 160 
rect 3 160 4 161 
rect 3 161 4 162 
rect 3 162 4 163 
rect 3 163 4 164 
rect 3 164 4 165 
rect 3 165 4 166 
rect 3 166 4 167 
rect 3 167 4 168 
rect 3 168 4 169 
rect 3 169 4 170 
rect 3 170 4 171 
rect 3 171 4 172 
rect 3 172 4 173 
rect 3 173 4 174 
rect 3 174 4 175 
rect 3 175 4 176 
rect 3 176 4 177 
rect 3 177 4 178 
rect 3 178 4 179 
rect 3 179 4 180 
rect 3 180 4 181 
rect 3 181 4 182 
rect 3 182 4 183 
rect 3 183 4 184 
rect 3 184 4 185 
rect 3 185 4 186 
rect 3 186 4 187 
rect 3 187 4 188 
rect 3 188 4 189 
rect 3 189 4 190 
rect 3 190 4 191 
rect 3 191 4 192 
rect 3 192 4 193 
rect 3 193 4 194 
rect 3 194 4 195 
rect 3 195 4 196 
rect 3 196 4 197 
rect 3 197 4 198 
rect 3 198 4 199 
rect 3 199 4 200 
rect 3 200 4 201 
rect 3 201 4 202 
rect 3 202 4 203 
rect 3 203 4 204 
rect 3 204 4 205 
rect 3 205 4 206 
rect 3 206 4 207 
rect 3 207 4 208 
rect 3 208 4 209 
rect 3 209 4 210 
rect 3 210 4 211 
rect 3 211 4 212 
rect 3 212 4 213 
rect 3 213 4 214 
rect 3 214 4 215 
rect 3 215 4 216 
rect 3 216 4 217 
rect 3 217 4 218 
rect 3 218 4 219 
rect 3 219 4 220 
rect 3 220 4 221 
rect 3 221 4 222 
rect 3 222 4 223 
rect 3 223 4 224 
rect 3 224 4 225 
rect 3 225 4 226 
rect 3 226 4 227 
rect 3 227 4 228 
rect 3 228 4 229 
rect 3 229 4 230 
rect 3 230 4 231 
rect 3 231 4 232 
rect 3 232 4 233 
rect 3 233 4 234 
rect 3 234 4 235 
rect 3 235 4 236 
rect 3 236 4 237 
rect 3 237 4 238 
rect 3 238 4 239 
rect 3 239 4 240 
rect 3 240 4 241 
rect 4 56 5 57 
rect 4 135 5 136 
rect 4 240 5 241 
rect 5 56 6 57 
rect 5 135 6 136 
rect 5 240 6 241 
rect 6 56 7 57 
rect 6 135 7 136 
rect 6 240 7 241 
rect 6 241 7 242 
rect 6 242 7 243 
rect 6 243 7 244 
rect 6 244 7 245 
rect 6 245 7 246 
rect 6 246 7 247 
rect 6 247 7 248 
rect 6 248 7 249 
rect 6 249 7 250 
rect 6 250 7 251 
rect 6 251 7 252 
rect 6 252 7 253 
rect 7 55 8 56 
rect 7 56 8 57 
rect 7 135 8 136 
rect 7 252 8 253 
rect 7 253 8 254 
rect 8 25 9 26 
rect 8 26 9 27 
rect 8 27 9 28 
rect 8 28 9 29 
rect 8 29 9 30 
rect 8 30 9 31 
rect 8 31 9 32 
rect 8 32 9 33 
rect 8 33 9 34 
rect 8 34 9 35 
rect 8 35 9 36 
rect 8 36 9 37 
rect 8 37 9 38 
rect 8 38 9 39 
rect 8 39 9 40 
rect 8 40 9 41 
rect 8 41 9 42 
rect 8 42 9 43 
rect 8 43 9 44 
rect 8 44 9 45 
rect 8 45 9 46 
rect 8 46 9 47 
rect 8 47 9 48 
rect 8 48 9 49 
rect 8 49 9 50 
rect 8 50 9 51 
rect 8 51 9 52 
rect 8 52 9 53 
rect 8 53 9 54 
rect 8 54 9 55 
rect 8 55 9 56 
rect 8 57 9 58 
rect 8 58 9 59 
rect 8 59 9 60 
rect 8 60 9 61 
rect 8 61 9 62 
rect 8 62 9 63 
rect 8 63 9 64 
rect 8 64 9 65 
rect 8 65 9 66 
rect 8 66 9 67 
rect 8 67 9 68 
rect 8 68 9 69 
rect 8 69 9 70 
rect 8 70 9 71 
rect 8 71 9 72 
rect 8 72 9 73 
rect 8 73 9 74 
rect 8 74 9 75 
rect 8 75 9 76 
rect 8 76 9 77 
rect 8 77 9 78 
rect 8 78 9 79 
rect 8 79 9 80 
rect 8 80 9 81 
rect 8 81 9 82 
rect 8 82 9 83 
rect 8 83 9 84 
rect 8 84 9 85 
rect 8 85 9 86 
rect 8 86 9 87 
rect 8 87 9 88 
rect 8 88 9 89 
rect 8 89 9 90 
rect 8 90 9 91 
rect 8 91 9 92 
rect 8 92 9 93 
rect 8 93 9 94 
rect 8 94 9 95 
rect 8 95 9 96 
rect 8 96 9 97 
rect 8 97 9 98 
rect 8 98 9 99 
rect 8 99 9 100 
rect 8 100 9 101 
rect 8 101 9 102 
rect 8 102 9 103 
rect 8 103 9 104 
rect 8 104 9 105 
rect 8 105 9 106 
rect 8 106 9 107 
rect 8 107 9 108 
rect 8 108 9 109 
rect 8 109 9 110 
rect 8 110 9 111 
rect 8 111 9 112 
rect 8 112 9 113 
rect 8 113 9 114 
rect 8 114 9 115 
rect 8 115 9 116 
rect 8 116 9 117 
rect 8 117 9 118 
rect 8 118 9 119 
rect 8 119 9 120 
rect 8 120 9 121 
rect 8 121 9 122 
rect 8 122 9 123 
rect 8 123 9 124 
rect 8 124 9 125 
rect 8 125 9 126 
rect 8 126 9 127 
rect 8 127 9 128 
rect 8 128 9 129 
rect 8 129 9 130 
rect 8 130 9 131 
rect 8 131 9 132 
rect 8 132 9 133 
rect 8 133 9 134 
rect 8 134 9 135 
rect 8 135 9 136 
rect 8 137 9 138 
rect 8 138 9 139 
rect 8 139 9 140 
rect 8 142 9 143 
rect 8 143 9 144 
rect 8 144 9 145 
rect 8 145 9 146 
rect 8 146 9 147 
rect 8 147 9 148 
rect 8 148 9 149 
rect 8 149 9 150 
rect 8 150 9 151 
rect 8 151 9 152 
rect 8 152 9 153 
rect 8 153 9 154 
rect 8 154 9 155 
rect 8 155 9 156 
rect 8 156 9 157 
rect 8 157 9 158 
rect 8 158 9 159 
rect 8 159 9 160 
rect 8 160 9 161 
rect 8 161 9 162 
rect 8 162 9 163 
rect 8 163 9 164 
rect 8 164 9 165 
rect 8 165 9 166 
rect 8 166 9 167 
rect 8 167 9 168 
rect 8 168 9 169 
rect 8 169 9 170 
rect 8 170 9 171 
rect 8 171 9 172 
rect 8 172 9 173 
rect 8 173 9 174 
rect 8 174 9 175 
rect 8 175 9 176 
rect 8 176 9 177 
rect 8 177 9 178 
rect 8 178 9 179 
rect 8 179 9 180 
rect 8 180 9 181 
rect 8 181 9 182 
rect 8 182 9 183 
rect 8 183 9 184 
rect 8 184 9 185 
rect 8 185 9 186 
rect 8 186 9 187 
rect 8 187 9 188 
rect 8 188 9 189 
rect 8 189 9 190 
rect 8 190 9 191 
rect 8 191 9 192 
rect 8 192 9 193 
rect 8 193 9 194 
rect 8 194 9 195 
rect 8 195 9 196 
rect 8 196 9 197 
rect 8 197 9 198 
rect 8 198 9 199 
rect 8 199 9 200 
rect 8 200 9 201 
rect 8 201 9 202 
rect 8 202 9 203 
rect 8 203 9 204 
rect 8 205 9 206 
rect 8 206 9 207 
rect 8 217 9 218 
rect 8 218 9 219 
rect 8 219 9 220 
rect 8 235 9 236 
rect 8 236 9 237 
rect 8 237 9 238 
rect 8 238 9 239 
rect 8 239 9 240 
rect 8 240 9 241 
rect 8 241 9 242 
rect 8 242 9 243 
rect 8 243 9 244 
rect 8 244 9 245 
rect 8 245 9 246 
rect 8 246 9 247 
rect 8 247 9 248 
rect 8 248 9 249 
rect 8 249 9 250 
rect 8 250 9 251 
rect 8 251 9 252 
rect 8 253 9 254 
rect 8 254 9 255 
rect 8 255 9 256 
rect 8 256 9 257 
rect 8 257 9 258 
rect 8 258 9 259 
rect 8 259 9 260 
rect 8 260 9 261 
rect 8 261 9 262 
rect 8 262 9 263 
rect 8 263 9 264 
rect 8 264 9 265 
rect 8 265 9 266 
rect 8 266 9 267 
rect 8 267 9 268 
rect 8 268 9 269 
rect 8 269 9 270 
rect 8 270 9 271 
rect 8 271 9 272 
rect 8 272 9 273 
rect 8 273 9 274 
rect 8 274 9 275 
rect 8 275 9 276 
rect 8 276 9 277 
rect 8 277 9 278 
rect 8 278 9 279 
rect 8 279 9 280 
rect 8 280 9 281 
rect 8 281 9 282 
rect 8 282 9 283 
rect 8 283 9 284 
rect 8 284 9 285 
rect 8 285 9 286 
rect 8 286 9 287 
rect 8 287 9 288 
rect 8 288 9 289 
rect 8 289 9 290 
rect 8 290 9 291 
rect 8 291 9 292 
rect 8 292 9 293 
rect 8 293 9 294 
rect 8 294 9 295 
rect 8 295 9 296 
rect 8 296 9 297 
rect 8 297 9 298 
rect 8 298 9 299 
rect 8 299 9 300 
rect 9 24 10 25 
rect 9 25 10 26 
rect 9 56 10 57 
rect 9 57 10 58 
rect 9 136 10 137 
rect 9 137 10 138 
rect 9 139 10 140 
rect 9 142 10 143 
rect 9 203 10 204 
rect 9 206 10 207 
rect 9 216 10 217 
rect 9 217 10 218 
rect 9 219 10 220 
rect 9 235 10 236 
rect 9 251 10 252 
rect 9 299 10 300 
rect 10 17 11 18 
rect 10 18 11 19 
rect 10 19 11 20 
rect 10 20 11 21 
rect 10 21 11 22 
rect 10 22 11 23 
rect 10 23 11 24 
rect 10 24 11 25 
rect 10 54 11 55 
rect 10 55 11 56 
rect 10 56 11 57 
rect 10 136 11 137 
rect 10 139 11 140 
rect 10 142 11 143 
rect 10 203 11 204 
rect 10 206 11 207 
rect 10 216 11 217 
rect 10 219 11 220 
rect 10 235 11 236 
rect 10 251 11 252 
rect 10 299 11 300 
rect 11 17 12 18 
rect 11 54 12 55 
rect 11 136 12 137 
rect 11 216 12 217 
rect 12 17 13 18 
rect 12 54 13 55 
rect 12 136 13 137 
rect 12 216 13 217 
rect 13 17 14 18 
rect 13 54 14 55 
rect 13 136 14 137 
rect 13 216 14 217 
rect 14 17 15 18 
rect 14 54 15 55 
rect 14 136 15 137 
rect 14 216 15 217 
rect 15 17 16 18 
rect 15 54 16 55 
rect 15 78 16 79 
rect 15 107 16 108 
rect 15 136 16 137 
rect 15 139 16 140 
rect 15 174 16 175 
rect 15 190 16 191 
rect 15 216 16 217 
rect 15 286 16 287 
rect 16 16 17 17 
rect 16 17 17 18 
rect 16 54 17 55 
rect 16 78 17 79 
rect 16 107 17 108 
rect 16 136 17 137 
rect 16 139 17 140 
rect 16 174 17 175 
rect 16 190 17 191 
rect 16 216 17 217 
rect 16 225 17 226 
rect 16 226 17 227 
rect 16 227 17 228 
rect 16 228 17 229 
rect 16 229 17 230 
rect 16 230 17 231 
rect 16 231 17 232 
rect 16 232 17 233 
rect 16 233 17 234 
rect 16 286 17 287 
rect 16 289 17 290 
rect 16 290 17 291 
rect 16 291 17 292 
rect 16 292 17 293 
rect 16 293 17 294 
rect 16 294 17 295 
rect 16 295 17 296 
rect 16 296 17 297 
rect 16 297 17 298 
rect 17 14 18 15 
rect 17 15 18 16 
rect 17 16 18 17 
rect 17 54 18 55 
rect 17 78 18 79 
rect 17 79 18 80 
rect 17 80 18 81 
rect 17 81 18 82 
rect 17 82 18 83 
rect 17 83 18 84 
rect 17 84 18 85 
rect 17 85 18 86 
rect 17 86 18 87 
rect 17 87 18 88 
rect 17 88 18 89 
rect 17 89 18 90 
rect 17 90 18 91 
rect 17 91 18 92 
rect 17 92 18 93 
rect 17 93 18 94 
rect 17 94 18 95 
rect 17 95 18 96 
rect 17 96 18 97 
rect 17 97 18 98 
rect 17 98 18 99 
rect 17 99 18 100 
rect 17 107 18 108 
rect 17 108 18 109 
rect 17 109 18 110 
rect 17 110 18 111 
rect 17 111 18 112 
rect 17 112 18 113 
rect 17 113 18 114 
rect 17 114 18 115 
rect 17 115 18 116 
rect 17 116 18 117 
rect 17 117 18 118 
rect 17 118 18 119 
rect 17 119 18 120 
rect 17 120 18 121 
rect 17 121 18 122 
rect 17 122 18 123 
rect 17 123 18 124 
rect 17 124 18 125 
rect 17 125 18 126 
rect 17 126 18 127 
rect 17 127 18 128 
rect 17 128 18 129 
rect 17 129 18 130 
rect 17 130 18 131 
rect 17 131 18 132 
rect 17 132 18 133 
rect 17 133 18 134 
rect 17 134 18 135 
rect 17 136 18 137 
rect 17 139 18 140 
rect 17 140 18 141 
rect 17 141 18 142 
rect 17 142 18 143 
rect 17 143 18 144 
rect 17 144 18 145 
rect 17 145 18 146 
rect 17 146 18 147 
rect 17 147 18 148 
rect 17 148 18 149 
rect 17 149 18 150 
rect 17 150 18 151 
rect 17 151 18 152 
rect 17 152 18 153 
rect 17 153 18 154 
rect 17 154 18 155 
rect 17 155 18 156 
rect 17 156 18 157 
rect 17 157 18 158 
rect 17 158 18 159 
rect 17 159 18 160 
rect 17 160 18 161 
rect 17 161 18 162 
rect 17 162 18 163 
rect 17 163 18 164 
rect 17 174 18 175 
rect 17 190 18 191 
rect 17 191 18 192 
rect 17 192 18 193 
rect 17 193 18 194 
rect 17 194 18 195 
rect 17 195 18 196 
rect 17 196 18 197 
rect 17 197 18 198 
rect 17 198 18 199 
rect 17 199 18 200 
rect 17 200 18 201 
rect 17 201 18 202 
rect 17 202 18 203 
rect 17 203 18 204 
rect 17 204 18 205 
rect 17 205 18 206 
rect 17 206 18 207 
rect 17 207 18 208 
rect 17 208 18 209 
rect 17 209 18 210 
rect 17 210 18 211 
rect 17 211 18 212 
rect 17 212 18 213 
rect 17 213 18 214 
rect 17 214 18 215 
rect 17 216 18 217 
rect 17 219 18 220 
rect 17 220 18 221 
rect 17 221 18 222 
rect 17 222 18 223 
rect 17 223 18 224 
rect 17 224 18 225 
rect 17 225 18 226 
rect 17 233 18 234 
rect 17 234 18 235 
rect 17 235 18 236 
rect 17 236 18 237 
rect 17 237 18 238 
rect 17 238 18 239 
rect 17 239 18 240 
rect 17 240 18 241 
rect 17 241 18 242 
rect 17 242 18 243 
rect 17 243 18 244 
rect 17 244 18 245 
rect 17 245 18 246 
rect 17 246 18 247 
rect 17 247 18 248 
rect 17 248 18 249 
rect 17 249 18 250 
rect 17 250 18 251 
rect 17 251 18 252 
rect 17 252 18 253 
rect 17 253 18 254 
rect 17 254 18 255 
rect 17 255 18 256 
rect 17 256 18 257 
rect 17 257 18 258 
rect 17 258 18 259 
rect 17 259 18 260 
rect 17 260 18 261 
rect 17 261 18 262 
rect 17 262 18 263 
rect 17 263 18 264 
rect 17 264 18 265 
rect 17 265 18 266 
rect 17 266 18 267 
rect 17 267 18 268 
rect 17 268 18 269 
rect 17 269 18 270 
rect 17 270 18 271 
rect 17 271 18 272 
rect 17 272 18 273 
rect 17 273 18 274 
rect 17 274 18 275 
rect 17 275 18 276 
rect 17 276 18 277 
rect 17 277 18 278 
rect 17 278 18 279 
rect 17 279 18 280 
rect 17 280 18 281 
rect 17 281 18 282 
rect 17 282 18 283 
rect 17 283 18 284 
rect 17 284 18 285 
rect 17 286 18 287 
rect 17 289 18 290 
rect 17 297 18 298 
rect 17 298 18 299 
rect 17 299 18 300 
rect 17 300 18 301 
rect 17 301 18 302 
rect 17 302 18 303 
rect 18 14 19 15 
rect 18 54 19 55 
rect 18 99 19 100 
rect 18 134 19 135 
rect 18 136 19 137 
rect 18 163 19 164 
rect 18 167 19 168 
rect 18 168 19 169 
rect 18 169 19 170 
rect 18 170 19 171 
rect 18 171 19 172 
rect 18 172 19 173 
rect 18 174 19 175 
rect 18 216 19 217 
rect 18 286 19 287 
rect 18 302 19 303 
rect 19 14 20 15 
rect 19 54 20 55 
rect 19 99 20 100 
rect 19 134 20 135 
rect 19 136 20 137 
rect 19 148 20 149 
rect 19 149 20 150 
rect 19 150 20 151 
rect 19 151 20 152 
rect 19 152 20 153 
rect 19 153 20 154 
rect 19 154 20 155 
rect 19 155 20 156 
rect 19 156 20 157 
rect 19 157 20 158 
rect 19 158 20 159 
rect 19 159 20 160 
rect 19 160 20 161 
rect 19 161 20 162 
rect 19 163 20 164 
rect 19 166 20 167 
rect 19 167 20 168 
rect 19 174 20 175 
rect 19 216 20 217 
rect 19 286 20 287 
rect 19 302 20 303 
rect 20 14 21 15 
rect 20 54 21 55 
rect 20 99 21 100 
rect 20 134 21 135 
rect 20 136 21 137 
rect 20 148 21 149 
rect 20 163 21 164 
rect 20 169 21 170 
rect 20 170 21 171 
rect 20 171 21 172 
rect 20 172 21 173 
rect 20 173 21 174 
rect 20 174 21 175 
rect 20 216 21 217 
rect 20 217 21 218 
rect 20 218 21 219 
rect 20 286 21 287 
rect 20 302 21 303 
rect 21 14 22 15 
rect 21 54 22 55 
rect 21 99 22 100 
rect 21 134 22 135 
rect 21 136 22 137 
rect 21 148 22 149 
rect 21 153 22 154 
rect 21 154 22 155 
rect 21 155 22 156 
rect 21 156 22 157 
rect 21 157 22 158 
rect 21 158 22 159 
rect 21 159 22 160 
rect 21 163 22 164 
rect 21 286 22 287 
rect 21 302 22 303 
rect 22 14 23 15 
rect 22 54 23 55 
rect 22 74 23 75 
rect 22 75 23 76 
rect 22 76 23 77 
rect 22 77 23 78 
rect 22 78 23 79 
rect 22 79 23 80 
rect 22 80 23 81 
rect 22 81 23 82 
rect 22 82 23 83 
rect 22 83 23 84 
rect 22 84 23 85 
rect 22 85 23 86 
rect 22 86 23 87 
rect 22 87 23 88 
rect 22 88 23 89 
rect 22 89 23 90 
rect 22 90 23 91 
rect 22 91 23 92 
rect 22 92 23 93 
rect 22 93 23 94 
rect 22 94 23 95 
rect 22 95 23 96 
rect 22 96 23 97 
rect 22 97 23 98 
rect 22 99 23 100 
rect 22 134 23 135 
rect 22 136 23 137 
rect 22 148 23 149 
rect 22 153 23 154 
rect 22 159 23 160 
rect 22 160 23 161 
rect 22 163 23 164 
rect 22 165 23 166 
rect 22 166 23 167 
rect 22 167 23 168 
rect 22 168 23 169 
rect 22 169 23 170 
rect 22 170 23 171 
rect 22 171 23 172 
rect 22 172 23 173 
rect 22 173 23 174 
rect 22 174 23 175 
rect 22 175 23 176 
rect 22 176 23 177 
rect 22 177 23 178 
rect 22 178 23 179 
rect 22 179 23 180 
rect 22 180 23 181 
rect 22 181 23 182 
rect 22 182 23 183 
rect 22 183 23 184 
rect 22 184 23 185 
rect 22 185 23 186 
rect 22 186 23 187 
rect 22 187 23 188 
rect 22 188 23 189 
rect 22 189 23 190 
rect 22 190 23 191 
rect 22 191 23 192 
rect 22 192 23 193 
rect 22 193 23 194 
rect 22 194 23 195 
rect 22 195 23 196 
rect 22 196 23 197 
rect 22 197 23 198 
rect 22 198 23 199 
rect 22 199 23 200 
rect 22 200 23 201 
rect 22 201 23 202 
rect 22 202 23 203 
rect 22 203 23 204 
rect 22 204 23 205 
rect 22 205 23 206 
rect 22 206 23 207 
rect 22 207 23 208 
rect 22 208 23 209 
rect 22 209 23 210 
rect 22 210 23 211 
rect 22 211 23 212 
rect 22 212 23 213 
rect 22 213 23 214 
rect 22 214 23 215 
rect 22 215 23 216 
rect 22 216 23 217 
rect 22 217 23 218 
rect 22 218 23 219 
rect 22 219 23 220 
rect 22 220 23 221 
rect 22 221 23 222 
rect 22 222 23 223 
rect 22 223 23 224 
rect 22 224 23 225 
rect 22 225 23 226 
rect 22 226 23 227 
rect 22 227 23 228 
rect 22 228 23 229 
rect 22 229 23 230 
rect 22 230 23 231 
rect 22 231 23 232 
rect 22 232 23 233 
rect 22 233 23 234 
rect 22 234 23 235 
rect 22 235 23 236 
rect 22 236 23 237 
rect 22 237 23 238 
rect 22 238 23 239 
rect 22 239 23 240 
rect 22 240 23 241 
rect 22 241 23 242 
rect 22 242 23 243 
rect 22 243 23 244 
rect 22 244 23 245 
rect 22 245 23 246 
rect 22 246 23 247 
rect 22 247 23 248 
rect 22 248 23 249 
rect 22 249 23 250 
rect 22 250 23 251 
rect 22 251 23 252 
rect 22 252 23 253 
rect 22 286 23 287 
rect 22 302 23 303 
rect 22 303 23 304 
rect 22 304 23 305 
rect 22 305 23 306 
rect 23 14 24 15 
rect 23 54 24 55 
rect 23 73 24 74 
rect 23 74 24 75 
rect 23 99 24 100 
rect 23 134 24 135 
rect 23 136 24 137 
rect 23 140 24 141 
rect 23 141 24 142 
rect 23 142 24 143 
rect 23 143 24 144 
rect 23 144 24 145 
rect 23 145 24 146 
rect 23 146 24 147 
rect 23 147 24 148 
rect 23 148 24 149 
rect 23 153 24 154 
rect 23 163 24 164 
rect 23 252 24 253 
rect 23 253 24 254 
rect 23 286 24 287 
rect 23 305 24 306 
rect 23 306 24 307 
rect 24 9 25 10 
rect 24 10 25 11 
rect 24 11 25 12 
rect 24 12 25 13 
rect 24 13 25 14 
rect 24 14 25 15 
rect 24 54 25 55 
rect 24 57 25 58 
rect 24 58 25 59 
rect 24 59 25 60 
rect 24 60 25 61 
rect 24 61 25 62 
rect 24 62 25 63 
rect 24 63 25 64 
rect 24 64 25 65 
rect 24 65 25 66 
rect 24 66 25 67 
rect 24 67 25 68 
rect 24 68 25 69 
rect 24 69 25 70 
rect 24 70 25 71 
rect 24 71 25 72 
rect 24 72 25 73 
rect 24 73 25 74 
rect 24 75 25 76 
rect 24 76 25 77 
rect 24 77 25 78 
rect 24 78 25 79 
rect 24 79 25 80 
rect 24 80 25 81 
rect 24 81 25 82 
rect 24 82 25 83 
rect 24 83 25 84 
rect 24 84 25 85 
rect 24 85 25 86 
rect 24 86 25 87 
rect 24 87 25 88 
rect 24 88 25 89 
rect 24 89 25 90 
rect 24 90 25 91 
rect 24 91 25 92 
rect 24 92 25 93 
rect 24 93 25 94 
rect 24 94 25 95 
rect 24 95 25 96 
rect 24 96 25 97 
rect 24 99 25 100 
rect 24 134 25 135 
rect 24 136 25 137 
rect 24 139 25 140 
rect 24 140 25 141 
rect 24 153 25 154 
rect 24 163 25 164 
rect 24 168 25 169 
rect 24 171 25 172 
rect 24 172 25 173 
rect 24 173 25 174 
rect 24 174 25 175 
rect 24 175 25 176 
rect 24 176 25 177 
rect 24 177 25 178 
rect 24 178 25 179 
rect 24 179 25 180 
rect 24 180 25 181 
rect 24 181 25 182 
rect 24 182 25 183 
rect 24 183 25 184 
rect 24 184 25 185 
rect 24 185 25 186 
rect 24 186 25 187 
rect 24 187 25 188 
rect 24 188 25 189 
rect 24 189 25 190 
rect 24 190 25 191 
rect 24 191 25 192 
rect 24 192 25 193 
rect 24 193 25 194 
rect 24 194 25 195 
rect 24 195 25 196 
rect 24 196 25 197 
rect 24 197 25 198 
rect 24 198 25 199 
rect 24 199 25 200 
rect 24 201 25 202 
rect 24 202 25 203 
rect 24 203 25 204 
rect 24 206 25 207 
rect 24 207 25 208 
rect 24 208 25 209 
rect 24 209 25 210 
rect 24 210 25 211 
rect 24 219 25 220 
rect 24 249 25 250 
rect 24 250 25 251 
rect 24 251 25 252 
rect 24 253 25 254 
rect 24 254 25 255 
rect 24 255 25 256 
rect 24 256 25 257 
rect 24 257 25 258 
rect 24 258 25 259 
rect 24 259 25 260 
rect 24 260 25 261 
rect 24 261 25 262 
rect 24 262 25 263 
rect 24 263 25 264 
rect 24 264 25 265 
rect 24 265 25 266 
rect 24 266 25 267 
rect 24 267 25 268 
rect 24 268 25 269 
rect 24 269 25 270 
rect 24 270 25 271 
rect 24 271 25 272 
rect 24 272 25 273 
rect 24 286 25 287 
rect 24 287 25 288 
rect 24 288 25 289 
rect 24 299 25 300 
rect 24 300 25 301 
rect 24 301 25 302 
rect 24 302 25 303 
rect 24 303 25 304 
rect 24 304 25 305 
rect 24 306 25 307 
rect 24 307 25 308 
rect 25 8 26 9 
rect 25 9 26 10 
rect 25 54 26 55 
rect 25 56 26 57 
rect 25 57 26 58 
rect 25 75 26 76 
rect 25 96 26 97 
rect 25 97 26 98 
rect 25 99 26 100 
rect 25 132 26 133 
rect 25 134 26 135 
rect 25 136 26 137 
rect 25 152 26 153 
rect 25 153 26 154 
rect 25 163 26 164 
rect 25 168 26 169 
rect 25 200 26 201 
rect 25 201 26 202 
rect 25 203 26 204 
rect 25 210 26 211 
rect 25 219 26 220 
rect 25 248 26 249 
rect 25 249 26 250 
rect 25 251 26 252 
rect 25 272 26 273 
rect 25 273 26 274 
rect 25 288 26 289 
rect 25 289 26 290 
rect 25 299 26 300 
rect 25 304 26 305 
rect 25 305 26 306 
rect 25 307 26 308 
rect 26 8 27 9 
rect 26 54 27 55 
rect 26 56 27 57 
rect 26 75 27 76 
rect 26 97 27 98 
rect 26 99 27 100 
rect 26 132 27 133 
rect 26 134 27 135 
rect 26 136 27 137 
rect 26 152 27 153 
rect 26 163 27 164 
rect 26 168 27 169 
rect 26 200 27 201 
rect 26 203 27 204 
rect 26 210 27 211 
rect 26 219 27 220 
rect 26 244 27 245 
rect 26 245 27 246 
rect 26 246 27 247 
rect 26 247 27 248 
rect 26 248 27 249 
rect 26 251 27 252 
rect 26 273 27 274 
rect 26 289 27 290 
rect 26 299 27 300 
rect 26 305 27 306 
rect 26 307 27 308 
rect 27 8 28 9 
rect 27 54 28 55 
rect 27 56 28 57 
rect 27 99 28 100 
rect 27 101 28 102 
rect 27 132 28 133 
rect 27 134 28 135 
rect 27 136 28 137 
rect 27 152 28 153 
rect 27 163 28 164 
rect 27 168 28 169 
rect 27 200 28 201 
rect 27 210 28 211 
rect 27 244 28 245 
rect 27 273 28 274 
rect 27 289 28 290 
rect 27 305 28 306 
rect 27 307 28 308 
rect 28 8 29 9 
rect 28 54 29 55 
rect 28 56 29 57 
rect 28 99 29 100 
rect 28 101 29 102 
rect 28 132 29 133 
rect 28 134 29 135 
rect 28 136 29 137 
rect 28 152 29 153 
rect 28 163 29 164 
rect 28 168 29 169 
rect 28 200 29 201 
rect 28 210 29 211 
rect 28 244 29 245 
rect 28 273 29 274 
rect 28 289 29 290 
rect 28 305 29 306 
rect 28 307 29 308 
rect 29 8 30 9 
rect 29 54 30 55 
rect 29 56 30 57 
rect 29 99 30 100 
rect 29 101 30 102 
rect 29 126 30 127 
rect 29 127 30 128 
rect 29 128 30 129 
rect 29 129 30 130 
rect 29 130 30 131 
rect 29 131 30 132 
rect 29 132 30 133 
rect 29 134 30 135 
rect 29 136 30 137 
rect 29 152 30 153 
rect 29 163 30 164 
rect 29 168 30 169 
rect 29 200 30 201 
rect 29 210 30 211 
rect 29 244 30 245 
rect 29 273 30 274 
rect 29 289 30 290 
rect 29 305 30 306 
rect 29 307 30 308 
rect 30 8 31 9 
rect 30 54 31 55 
rect 30 56 31 57 
rect 30 99 31 100 
rect 30 101 31 102 
rect 30 124 31 125 
rect 30 125 31 126 
rect 30 126 31 127 
rect 30 134 31 135 
rect 30 136 31 137 
rect 30 152 31 153 
rect 30 163 31 164 
rect 30 168 31 169 
rect 30 200 31 201 
rect 30 210 31 211 
rect 30 244 31 245 
rect 30 273 31 274 
rect 30 289 31 290 
rect 30 305 31 306 
rect 30 307 31 308 
rect 31 8 32 9 
rect 31 14 32 15 
rect 31 54 32 55 
rect 31 56 32 57 
rect 31 59 32 60 
rect 31 62 32 63 
rect 31 99 32 100 
rect 31 101 32 102 
rect 31 134 32 135 
rect 31 136 32 137 
rect 31 145 32 146 
rect 31 146 32 147 
rect 31 147 32 148 
rect 31 148 32 149 
rect 31 149 32 150 
rect 31 150 32 151 
rect 31 151 32 152 
rect 31 152 32 153 
rect 31 155 32 156 
rect 31 161 32 162 
rect 31 163 32 164 
rect 31 168 32 169 
rect 31 200 32 201 
rect 31 210 32 211 
rect 31 222 32 223 
rect 31 235 32 236 
rect 31 244 32 245 
rect 31 251 32 252 
rect 31 273 32 274 
rect 31 283 32 284 
rect 31 289 32 290 
rect 31 299 32 300 
rect 31 305 32 306 
rect 31 307 32 308 
rect 32 8 33 9 
rect 32 14 33 15 
rect 32 54 33 55 
rect 32 56 33 57 
rect 32 59 33 60 
rect 32 62 33 63 
rect 32 99 33 100 
rect 32 101 33 102 
rect 32 102 33 103 
rect 32 103 33 104 
rect 32 104 33 105 
rect 32 105 33 106 
rect 32 112 33 113 
rect 32 113 33 114 
rect 32 114 33 115 
rect 32 115 33 116 
rect 32 116 33 117 
rect 32 117 33 118 
rect 32 118 33 119 
rect 32 119 33 120 
rect 32 120 33 121 
rect 32 121 33 122 
rect 32 122 33 123 
rect 32 123 33 124 
rect 32 124 33 125 
rect 32 125 33 126 
rect 32 126 33 127 
rect 32 127 33 128 
rect 32 128 33 129 
rect 32 129 33 130 
rect 32 130 33 131 
rect 32 134 33 135 
rect 32 136 33 137 
rect 32 145 33 146 
rect 32 155 33 156 
rect 32 161 33 162 
rect 32 163 33 164 
rect 32 165 33 166 
rect 32 166 33 167 
rect 32 167 33 168 
rect 32 168 33 169 
rect 32 200 33 201 
rect 32 210 33 211 
rect 32 222 33 223 
rect 32 235 33 236 
rect 32 244 33 245 
rect 32 251 33 252 
rect 32 273 33 274 
rect 32 274 33 275 
rect 32 275 33 276 
rect 32 276 33 277 
rect 32 277 33 278 
rect 32 278 33 279 
rect 32 279 33 280 
rect 32 280 33 281 
rect 32 281 33 282 
rect 32 283 33 284 
rect 32 289 33 290 
rect 32 299 33 300 
rect 32 305 33 306 
rect 32 307 33 308 
rect 33 8 34 9 
rect 33 14 34 15 
rect 33 54 34 55 
rect 33 56 34 57 
rect 33 59 34 60 
rect 33 62 34 63 
rect 33 63 34 64 
rect 33 64 34 65 
rect 33 65 34 66 
rect 33 66 34 67 
rect 33 67 34 68 
rect 33 99 34 100 
rect 33 105 34 106 
rect 33 106 34 107 
rect 33 107 34 108 
rect 33 108 34 109 
rect 33 109 34 110 
rect 33 110 34 111 
rect 33 111 34 112 
rect 33 112 34 113 
rect 33 130 34 131 
rect 33 134 34 135 
rect 33 136 34 137 
rect 33 145 34 146 
rect 33 155 34 156 
rect 33 161 34 162 
rect 33 163 34 164 
rect 33 165 34 166 
rect 33 200 34 201 
rect 33 210 34 211 
rect 33 222 34 223 
rect 33 235 34 236 
rect 33 244 34 245 
rect 33 251 34 252 
rect 33 281 34 282 
rect 33 282 34 283 
rect 33 283 34 284 
rect 33 289 34 290 
rect 33 299 34 300 
rect 33 305 34 306 
rect 33 307 34 308 
rect 34 8 35 9 
rect 34 14 35 15 
rect 34 54 35 55 
rect 34 56 35 57 
rect 34 59 35 60 
rect 34 67 35 68 
rect 34 99 35 100 
rect 34 130 35 131 
rect 34 134 35 135 
rect 34 136 35 137 
rect 34 145 35 146 
rect 34 155 35 156 
rect 34 161 35 162 
rect 34 163 35 164 
rect 34 165 35 166 
rect 34 200 35 201 
rect 34 210 35 211 
rect 34 222 35 223 
rect 34 235 35 236 
rect 34 244 35 245 
rect 34 251 35 252 
rect 34 289 35 290 
rect 34 299 35 300 
rect 34 305 35 306 
rect 34 307 35 308 
rect 35 8 36 9 
rect 35 14 36 15 
rect 35 54 36 55 
rect 35 56 36 57 
rect 35 59 36 60 
rect 35 155 36 156 
rect 35 161 36 162 
rect 35 163 36 164 
rect 35 165 36 166 
rect 35 200 36 201 
rect 35 210 36 211 
rect 35 222 36 223 
rect 35 235 36 236 
rect 35 244 36 245 
rect 35 251 36 252 
rect 35 289 36 290 
rect 35 299 36 300 
rect 35 305 36 306 
rect 35 307 36 308 
rect 36 8 37 9 
rect 36 11 37 12 
rect 36 12 37 13 
rect 36 13 37 14 
rect 36 14 37 15 
rect 36 54 37 55 
rect 36 56 37 57 
rect 36 59 37 60 
rect 36 60 37 61 
rect 36 61 37 62 
rect 36 62 37 63 
rect 36 63 37 64 
rect 36 64 37 65 
rect 36 65 37 66 
rect 36 66 37 67 
rect 36 67 37 68 
rect 36 68 37 69 
rect 36 69 37 70 
rect 36 70 37 71 
rect 36 71 37 72 
rect 36 72 37 73 
rect 36 73 37 74 
rect 36 74 37 75 
rect 36 75 37 76 
rect 36 76 37 77 
rect 36 77 37 78 
rect 36 78 37 79 
rect 36 79 37 80 
rect 36 80 37 81 
rect 36 82 37 83 
rect 36 83 37 84 
rect 36 84 37 85 
rect 36 85 37 86 
rect 36 86 37 87 
rect 36 87 37 88 
rect 36 88 37 89 
rect 36 89 37 90 
rect 36 90 37 91 
rect 36 91 37 92 
rect 36 92 37 93 
rect 36 93 37 94 
rect 36 94 37 95 
rect 36 95 37 96 
rect 36 96 37 97 
rect 36 97 37 98 
rect 36 98 37 99 
rect 36 99 37 100 
rect 36 100 37 101 
rect 36 101 37 102 
rect 36 102 37 103 
rect 36 103 37 104 
rect 36 104 37 105 
rect 36 105 37 106 
rect 36 106 37 107 
rect 36 107 37 108 
rect 36 108 37 109 
rect 36 109 37 110 
rect 36 110 37 111 
rect 36 111 37 112 
rect 36 112 37 113 
rect 36 113 37 114 
rect 36 114 37 115 
rect 36 115 37 116 
rect 36 116 37 117 
rect 36 117 37 118 
rect 36 118 37 119 
rect 36 119 37 120 
rect 36 120 37 121 
rect 36 121 37 122 
rect 36 122 37 123 
rect 36 123 37 124 
rect 36 124 37 125 
rect 36 125 37 126 
rect 36 126 37 127 
rect 36 127 37 128 
rect 36 128 37 129 
rect 36 129 37 130 
rect 36 130 37 131 
rect 36 131 37 132 
rect 36 132 37 133 
rect 36 133 37 134 
rect 36 134 37 135 
rect 36 135 37 136 
rect 36 136 37 137 
rect 36 137 37 138 
rect 36 138 37 139 
rect 36 139 37 140 
rect 36 140 37 141 
rect 36 141 37 142 
rect 36 142 37 143 
rect 36 143 37 144 
rect 36 144 37 145 
rect 36 145 37 146 
rect 36 146 37 147 
rect 36 147 37 148 
rect 36 148 37 149 
rect 36 149 37 150 
rect 36 150 37 151 
rect 36 151 37 152 
rect 36 152 37 153 
rect 36 153 37 154 
rect 36 154 37 155 
rect 36 155 37 156 
rect 36 158 37 159 
rect 36 159 37 160 
rect 36 160 37 161 
rect 36 161 37 162 
rect 36 163 37 164 
rect 36 210 37 211 
rect 36 215 37 216 
rect 36 216 37 217 
rect 36 217 37 218 
rect 36 218 37 219 
rect 36 219 37 220 
rect 36 220 37 221 
rect 36 221 37 222 
rect 36 222 37 223 
rect 36 235 37 236 
rect 36 244 37 245 
rect 36 246 37 247 
rect 36 247 37 248 
rect 36 248 37 249 
rect 36 249 37 250 
rect 36 250 37 251 
rect 36 251 37 252 
rect 36 289 37 290 
rect 36 292 37 293 
rect 36 293 37 294 
rect 36 294 37 295 
rect 36 295 37 296 
rect 36 296 37 297 
rect 36 297 37 298 
rect 36 298 37 299 
rect 36 299 37 300 
rect 36 305 37 306 
rect 36 307 37 308 
rect 37 8 38 9 
rect 37 11 38 12 
rect 37 54 38 55 
rect 37 56 38 57 
rect 37 80 38 81 
rect 37 82 38 83 
rect 37 163 38 164 
rect 37 166 38 167 
rect 37 167 38 168 
rect 37 168 38 169 
rect 37 169 38 170 
rect 37 170 38 171 
rect 37 171 38 172 
rect 37 172 38 173 
rect 37 173 38 174 
rect 37 174 38 175 
rect 37 175 38 176 
rect 37 176 38 177 
rect 37 177 38 178 
rect 37 178 38 179 
rect 37 179 38 180 
rect 37 180 38 181 
rect 37 181 38 182 
rect 37 182 38 183 
rect 37 183 38 184 
rect 37 184 38 185 
rect 37 185 38 186 
rect 37 186 38 187 
rect 37 187 38 188 
rect 37 188 38 189 
rect 37 189 38 190 
rect 37 190 38 191 
rect 37 191 38 192 
rect 37 192 38 193 
rect 37 193 38 194 
rect 37 194 38 195 
rect 37 195 38 196 
rect 37 196 38 197 
rect 37 197 38 198 
rect 37 198 38 199 
rect 37 199 38 200 
rect 37 200 38 201 
rect 37 201 38 202 
rect 37 202 38 203 
rect 37 203 38 204 
rect 37 204 38 205 
rect 37 205 38 206 
rect 37 206 38 207 
rect 37 210 38 211 
rect 37 215 38 216 
rect 37 235 38 236 
rect 37 244 38 245 
rect 37 246 38 247 
rect 37 289 38 290 
rect 37 292 38 293 
rect 37 305 38 306 
rect 37 307 38 308 
rect 38 8 39 9 
rect 38 11 39 12 
rect 38 54 39 55 
rect 38 56 39 57 
rect 38 80 39 81 
rect 38 82 39 83 
rect 38 85 39 86 
rect 38 86 39 87 
rect 38 87 39 88 
rect 38 88 39 89 
rect 38 89 39 90 
rect 38 90 39 91 
rect 38 91 39 92 
rect 38 92 39 93 
rect 38 93 39 94 
rect 38 94 39 95 
rect 38 95 39 96 
rect 38 96 39 97 
rect 38 97 39 98 
rect 38 98 39 99 
rect 38 99 39 100 
rect 38 100 39 101 
rect 38 101 39 102 
rect 38 102 39 103 
rect 38 103 39 104 
rect 38 104 39 105 
rect 38 105 39 106 
rect 38 106 39 107 
rect 38 107 39 108 
rect 38 108 39 109 
rect 38 109 39 110 
rect 38 110 39 111 
rect 38 111 39 112 
rect 38 112 39 113 
rect 38 113 39 114 
rect 38 114 39 115 
rect 38 115 39 116 
rect 38 116 39 117 
rect 38 117 39 118 
rect 38 118 39 119 
rect 38 119 39 120 
rect 38 120 39 121 
rect 38 121 39 122 
rect 38 122 39 123 
rect 38 123 39 124 
rect 38 124 39 125 
rect 38 125 39 126 
rect 38 126 39 127 
rect 38 127 39 128 
rect 38 128 39 129 
rect 38 129 39 130 
rect 38 130 39 131 
rect 38 131 39 132 
rect 38 132 39 133 
rect 38 135 39 136 
rect 38 136 39 137 
rect 38 137 39 138 
rect 38 138 39 139 
rect 38 139 39 140 
rect 38 140 39 141 
rect 38 141 39 142 
rect 38 142 39 143 
rect 38 143 39 144 
rect 38 144 39 145 
rect 38 145 39 146 
rect 38 146 39 147 
rect 38 147 39 148 
rect 38 148 39 149 
rect 38 149 39 150 
rect 38 150 39 151 
rect 38 151 39 152 
rect 38 152 39 153 
rect 38 153 39 154 
rect 38 154 39 155 
rect 38 155 39 156 
rect 38 156 39 157 
rect 38 157 39 158 
rect 38 158 39 159 
rect 38 159 39 160 
rect 38 160 39 161 
rect 38 161 39 162 
rect 38 163 39 164 
rect 38 166 39 167 
rect 38 206 39 207 
rect 38 210 39 211 
rect 38 215 39 216 
rect 38 235 39 236 
rect 38 244 39 245 
rect 38 246 39 247 
rect 38 289 39 290 
rect 38 292 39 293 
rect 38 305 39 306 
rect 38 307 39 308 
rect 39 7 40 8 
rect 39 8 40 9 
rect 39 11 40 12 
rect 39 54 40 55 
rect 39 56 40 57 
rect 39 82 40 83 
rect 39 163 40 164 
rect 39 194 40 195 
rect 39 206 40 207 
rect 39 210 40 211 
rect 39 215 40 216 
rect 39 235 40 236 
rect 39 244 40 245 
rect 39 246 40 247 
rect 39 289 40 290 
rect 39 292 40 293 
rect 39 305 40 306 
rect 39 307 40 308 
rect 40 3 41 4 
rect 40 4 41 5 
rect 40 5 41 6 
rect 40 6 41 7 
rect 40 7 41 8 
rect 40 9 41 10 
rect 40 10 41 11 
rect 40 11 41 12 
rect 40 43 41 44 
rect 40 44 41 45 
rect 40 45 41 46 
rect 40 46 41 47 
rect 40 47 41 48 
rect 40 48 41 49 
rect 40 54 41 55 
rect 40 56 41 57 
rect 40 82 41 83 
rect 40 91 41 92 
rect 40 92 41 93 
rect 40 93 41 94 
rect 40 94 41 95 
rect 40 95 41 96 
rect 40 96 41 97 
rect 40 97 41 98 
rect 40 98 41 99 
rect 40 99 41 100 
rect 40 100 41 101 
rect 40 101 41 102 
rect 40 102 41 103 
rect 40 103 41 104 
rect 40 104 41 105 
rect 40 105 41 106 
rect 40 106 41 107 
rect 40 107 41 108 
rect 40 108 41 109 
rect 40 109 41 110 
rect 40 110 41 111 
rect 40 111 41 112 
rect 40 112 41 113 
rect 40 113 41 114 
rect 40 114 41 115 
rect 40 115 41 116 
rect 40 116 41 117 
rect 40 117 41 118 
rect 40 118 41 119 
rect 40 119 41 120 
rect 40 120 41 121 
rect 40 121 41 122 
rect 40 122 41 123 
rect 40 123 41 124 
rect 40 124 41 125 
rect 40 125 41 126 
rect 40 126 41 127 
rect 40 127 41 128 
rect 40 128 41 129 
rect 40 129 41 130 
rect 40 130 41 131 
rect 40 131 41 132 
rect 40 132 41 133 
rect 40 133 41 134 
rect 40 134 41 135 
rect 40 135 41 136 
rect 40 136 41 137 
rect 40 137 41 138 
rect 40 138 41 139 
rect 40 139 41 140 
rect 40 140 41 141 
rect 40 141 41 142 
rect 40 142 41 143 
rect 40 143 41 144 
rect 40 144 41 145 
rect 40 153 41 154 
rect 40 154 41 155 
rect 40 155 41 156 
rect 40 156 41 157 
rect 40 157 41 158 
rect 40 158 41 159 
rect 40 159 41 160 
rect 40 160 41 161 
rect 40 163 41 164 
rect 40 165 41 166 
rect 40 166 41 167 
rect 40 167 41 168 
rect 40 168 41 169 
rect 40 169 41 170 
rect 40 170 41 171 
rect 40 171 41 172 
rect 40 187 41 188 
rect 40 188 41 189 
rect 40 189 41 190 
rect 40 190 41 191 
rect 40 191 41 192 
rect 40 192 41 193 
rect 40 194 41 195 
rect 40 195 41 196 
rect 40 206 41 207 
rect 40 210 41 211 
rect 40 215 41 216 
rect 40 219 41 220 
rect 40 220 41 221 
rect 40 221 41 222 
rect 40 222 41 223 
rect 40 223 41 224 
rect 40 224 41 225 
rect 40 233 41 234 
rect 40 234 41 235 
rect 40 235 41 236 
rect 40 244 41 245 
rect 40 246 41 247 
rect 40 254 41 255 
rect 40 255 41 256 
rect 40 256 41 257 
rect 40 267 41 268 
rect 40 268 41 269 
rect 40 269 41 270 
rect 40 270 41 271 
rect 40 271 41 272 
rect 40 272 41 273 
rect 40 289 41 290 
rect 40 292 41 293 
rect 40 305 41 306 
rect 40 307 41 308 
rect 41 3 42 4 
rect 41 8 42 9 
rect 41 9 42 10 
rect 41 43 42 44 
rect 41 48 42 49 
rect 41 49 42 50 
rect 41 54 42 55 
rect 41 56 42 57 
rect 41 82 42 83 
rect 41 91 42 92 
rect 41 152 42 153 
rect 41 153 42 154 
rect 41 163 42 164 
rect 41 171 42 172 
rect 41 187 42 188 
rect 41 192 42 193 
rect 41 193 42 194 
rect 41 195 42 196 
rect 41 206 42 207 
rect 41 210 42 211 
rect 41 215 42 216 
rect 41 219 42 220 
rect 41 224 42 225 
rect 41 225 42 226 
rect 41 232 42 233 
rect 41 233 42 234 
rect 41 244 42 245 
rect 41 246 42 247 
rect 41 254 42 255 
rect 41 256 42 257 
rect 41 257 42 258 
rect 41 267 42 268 
rect 41 272 42 273 
rect 41 273 42 274 
rect 41 289 42 290 
rect 41 292 42 293 
rect 41 305 42 306 
rect 41 307 42 308 
rect 42 3 43 4 
rect 42 8 43 9 
rect 42 43 43 44 
rect 42 49 43 50 
rect 42 54 43 55 
rect 42 56 43 57 
rect 42 82 43 83 
rect 42 91 43 92 
rect 42 97 43 98 
rect 42 98 43 99 
rect 42 99 43 100 
rect 42 100 43 101 
rect 42 101 43 102 
rect 42 102 43 103 
rect 42 103 43 104 
rect 42 113 43 114 
rect 42 145 43 146 
rect 42 146 43 147 
rect 42 147 43 148 
rect 42 148 43 149 
rect 42 149 43 150 
rect 42 150 43 151 
rect 42 151 43 152 
rect 42 152 43 153 
rect 42 163 43 164 
rect 42 171 43 172 
rect 42 187 43 188 
rect 42 193 43 194 
rect 42 195 43 196 
rect 42 206 43 207 
rect 42 210 43 211 
rect 42 215 43 216 
rect 42 219 43 220 
rect 42 225 43 226 
rect 42 226 43 227 
rect 42 227 43 228 
rect 42 228 43 229 
rect 42 232 43 233 
rect 42 244 43 245 
rect 42 246 43 247 
rect 42 254 43 255 
rect 42 257 43 258 
rect 42 267 43 268 
rect 42 273 43 274 
rect 42 289 43 290 
rect 42 292 43 293 
rect 42 305 43 306 
rect 42 307 43 308 
rect 43 3 44 4 
rect 43 8 44 9 
rect 43 49 44 50 
rect 43 54 44 55 
rect 43 56 44 57 
rect 43 82 44 83 
rect 43 113 44 114 
rect 43 145 44 146 
rect 43 163 44 164 
rect 43 193 44 194 
rect 43 195 44 196 
rect 43 210 44 211 
rect 43 215 44 216 
rect 43 228 44 229 
rect 43 232 44 233 
rect 43 244 44 245 
rect 43 246 44 247 
rect 43 257 44 258 
rect 43 273 44 274 
rect 43 289 44 290 
rect 43 292 44 293 
rect 43 305 44 306 
rect 43 307 44 308 
rect 44 3 45 4 
rect 44 8 45 9 
rect 44 49 45 50 
rect 44 54 45 55 
rect 44 56 45 57 
rect 44 82 45 83 
rect 44 113 45 114 
rect 44 145 45 146 
rect 44 163 45 164 
rect 44 193 45 194 
rect 44 195 45 196 
rect 44 210 45 211 
rect 44 215 45 216 
rect 44 228 45 229 
rect 44 232 45 233 
rect 44 244 45 245 
rect 44 246 45 247 
rect 44 257 45 258 
rect 44 273 45 274 
rect 44 289 45 290 
rect 44 292 45 293 
rect 44 305 45 306 
rect 44 307 45 308 
rect 45 3 46 4 
rect 45 8 46 9 
rect 45 49 46 50 
rect 45 54 46 55 
rect 45 82 46 83 
rect 45 113 46 114 
rect 45 145 46 146 
rect 45 163 46 164 
rect 45 193 46 194 
rect 45 195 46 196 
rect 45 210 46 211 
rect 45 215 46 216 
rect 45 228 46 229 
rect 45 232 46 233 
rect 45 244 46 245 
rect 45 246 46 247 
rect 45 257 46 258 
rect 45 273 46 274 
rect 45 289 46 290 
rect 45 292 46 293 
rect 45 305 46 306 
rect 45 307 46 308 
rect 46 3 47 4 
rect 46 8 47 9 
rect 46 49 47 50 
rect 46 54 47 55 
rect 46 82 47 83 
rect 46 113 47 114 
rect 46 114 47 115 
rect 46 145 47 146 
rect 46 163 47 164 
rect 46 193 47 194 
rect 46 195 47 196 
rect 46 210 47 211 
rect 46 211 47 212 
rect 46 212 47 213 
rect 46 215 47 216 
rect 46 228 47 229 
rect 46 232 47 233 
rect 46 244 47 245 
rect 46 246 47 247 
rect 46 257 47 258 
rect 46 273 47 274 
rect 46 289 47 290 
rect 46 292 47 293 
rect 46 305 47 306 
rect 46 307 47 308 
rect 47 3 48 4 
rect 47 8 48 9 
rect 47 49 48 50 
rect 47 54 48 55 
rect 47 82 48 83 
rect 47 114 48 115 
rect 47 115 48 116 
rect 47 163 48 164 
rect 47 193 48 194 
rect 47 195 48 196 
rect 47 196 48 197 
rect 47 197 48 198 
rect 47 232 48 233 
rect 47 244 48 245 
rect 47 246 48 247 
rect 47 257 48 258 
rect 47 270 48 271 
rect 47 273 48 274 
rect 47 289 48 290 
rect 47 292 48 293 
rect 47 305 48 306 
rect 47 307 48 308 
rect 48 3 49 4 
rect 48 8 49 9 
rect 48 82 49 83 
rect 48 97 49 98 
rect 48 98 49 99 
rect 48 99 49 100 
rect 48 100 49 101 
rect 48 101 49 102 
rect 48 144 49 145 
rect 48 145 49 146 
rect 48 146 49 147 
rect 48 147 49 148 
rect 48 148 49 149 
rect 48 149 49 150 
rect 48 150 49 151 
rect 48 151 49 152 
rect 48 152 49 153 
rect 48 163 49 164 
rect 48 208 49 209 
rect 48 209 49 210 
rect 48 210 49 211 
rect 48 211 49 212 
rect 48 212 49 213 
rect 48 213 49 214 
rect 48 214 49 215 
rect 48 215 49 216 
rect 48 216 49 217 
rect 48 224 49 225 
rect 48 225 49 226 
rect 48 226 49 227 
rect 48 227 49 228 
rect 48 228 49 229 
rect 48 229 49 230 
rect 48 230 49 231 
rect 48 232 49 233 
rect 48 244 49 245 
rect 48 246 49 247 
rect 48 257 49 258 
rect 48 270 49 271 
rect 48 273 49 274 
rect 48 289 49 290 
rect 48 292 49 293 
rect 48 305 49 306 
rect 48 307 49 308 
rect 49 3 50 4 
rect 49 8 50 9 
rect 49 18 50 19 
rect 49 19 50 20 
rect 49 20 50 21 
rect 49 21 50 22 
rect 49 22 50 23 
rect 49 23 50 24 
rect 49 24 50 25 
rect 49 25 50 26 
rect 49 26 50 27 
rect 49 27 50 28 
rect 49 28 50 29 
rect 49 29 50 30 
rect 49 30 50 31 
rect 49 31 50 32 
rect 49 32 50 33 
rect 49 33 50 34 
rect 49 34 50 35 
rect 49 35 50 36 
rect 49 36 50 37 
rect 49 37 50 38 
rect 49 38 50 39 
rect 49 39 50 40 
rect 49 40 50 41 
rect 49 41 50 42 
rect 49 42 50 43 
rect 49 43 50 44 
rect 49 44 50 45 
rect 49 45 50 46 
rect 49 46 50 47 
rect 49 47 50 48 
rect 49 48 50 49 
rect 49 49 50 50 
rect 49 50 50 51 
rect 49 51 50 52 
rect 49 52 50 53 
rect 49 53 50 54 
rect 49 54 50 55 
rect 49 55 50 56 
rect 49 56 50 57 
rect 49 57 50 58 
rect 49 58 50 59 
rect 49 59 50 60 
rect 49 60 50 61 
rect 49 61 50 62 
rect 49 62 50 63 
rect 49 63 50 64 
rect 49 64 50 65 
rect 49 65 50 66 
rect 49 66 50 67 
rect 49 67 50 68 
rect 49 68 50 69 
rect 49 69 50 70 
rect 49 70 50 71 
rect 49 71 50 72 
rect 49 72 50 73 
rect 49 73 50 74 
rect 49 74 50 75 
rect 49 75 50 76 
rect 49 76 50 77 
rect 49 77 50 78 
rect 49 78 50 79 
rect 49 79 50 80 
rect 49 82 50 83 
rect 49 103 50 104 
rect 49 104 50 105 
rect 49 105 50 106 
rect 49 106 50 107 
rect 49 107 50 108 
rect 49 108 50 109 
rect 49 109 50 110 
rect 49 110 50 111 
rect 49 111 50 112 
rect 49 112 50 113 
rect 49 113 50 114 
rect 49 114 50 115 
rect 49 115 50 116 
rect 49 116 50 117 
rect 49 117 50 118 
rect 49 118 50 119 
rect 49 119 50 120 
rect 49 120 50 121 
rect 49 121 50 122 
rect 49 122 50 123 
rect 49 123 50 124 
rect 49 124 50 125 
rect 49 125 50 126 
rect 49 126 50 127 
rect 49 127 50 128 
rect 49 128 50 129 
rect 49 129 50 130 
rect 49 130 50 131 
rect 49 131 50 132 
rect 49 132 50 133 
rect 49 133 50 134 
rect 49 134 50 135 
rect 49 135 50 136 
rect 49 136 50 137 
rect 49 137 50 138 
rect 49 138 50 139 
rect 49 139 50 140 
rect 49 140 50 141 
rect 49 141 50 142 
rect 49 142 50 143 
rect 49 143 50 144 
rect 49 144 50 145 
rect 49 152 50 153 
rect 49 153 50 154 
rect 49 154 50 155 
rect 49 155 50 156 
rect 49 156 50 157 
rect 49 157 50 158 
rect 49 158 50 159 
rect 49 159 50 160 
rect 49 160 50 161 
rect 49 163 50 164 
rect 49 165 50 166 
rect 49 166 50 167 
rect 49 167 50 168 
rect 49 168 50 169 
rect 49 169 50 170 
rect 49 170 50 171 
rect 49 171 50 172 
rect 49 172 50 173 
rect 49 173 50 174 
rect 49 174 50 175 
rect 49 175 50 176 
rect 49 176 50 177 
rect 49 177 50 178 
rect 49 178 50 179 
rect 49 179 50 180 
rect 49 180 50 181 
rect 49 181 50 182 
rect 49 182 50 183 
rect 49 183 50 184 
rect 49 184 50 185 
rect 49 185 50 186 
rect 49 186 50 187 
rect 49 187 50 188 
rect 49 188 50 189 
rect 49 189 50 190 
rect 49 190 50 191 
rect 49 191 50 192 
rect 49 192 50 193 
rect 49 193 50 194 
rect 49 194 50 195 
rect 49 195 50 196 
rect 49 196 50 197 
rect 49 197 50 198 
rect 49 198 50 199 
rect 49 199 50 200 
rect 49 200 50 201 
rect 49 201 50 202 
rect 49 202 50 203 
rect 49 203 50 204 
rect 49 204 50 205 
rect 49 205 50 206 
rect 49 206 50 207 
rect 49 207 50 208 
rect 49 208 50 209 
rect 49 216 50 217 
rect 49 217 50 218 
rect 49 218 50 219 
rect 49 219 50 220 
rect 49 220 50 221 
rect 49 221 50 222 
rect 49 222 50 223 
rect 49 223 50 224 
rect 49 224 50 225 
rect 49 232 50 233 
rect 49 244 50 245 
rect 49 246 50 247 
rect 49 257 50 258 
rect 49 261 50 262 
rect 49 262 50 263 
rect 49 263 50 264 
rect 49 264 50 265 
rect 49 265 50 266 
rect 49 266 50 267 
rect 49 267 50 268 
rect 49 268 50 269 
rect 49 269 50 270 
rect 49 270 50 271 
rect 49 273 50 274 
rect 49 289 50 290 
rect 49 292 50 293 
rect 49 305 50 306 
rect 49 307 50 308 
rect 50 3 51 4 
rect 50 8 51 9 
rect 50 18 51 19 
rect 50 79 51 80 
rect 50 82 51 83 
rect 50 84 51 85 
rect 50 85 51 86 
rect 50 86 51 87 
rect 50 87 51 88 
rect 50 88 51 89 
rect 50 89 51 90 
rect 50 90 51 91 
rect 50 91 51 92 
rect 50 92 51 93 
rect 50 93 51 94 
rect 50 94 51 95 
rect 50 95 51 96 
rect 50 96 51 97 
rect 50 97 51 98 
rect 50 98 51 99 
rect 50 99 51 100 
rect 50 100 51 101 
rect 50 103 51 104 
rect 50 163 51 164 
rect 50 210 51 211 
rect 50 211 51 212 
rect 50 212 51 213 
rect 50 213 51 214 
rect 50 214 51 215 
rect 50 232 51 233 
rect 50 234 51 235 
rect 50 235 51 236 
rect 50 236 51 237 
rect 50 237 51 238 
rect 50 238 51 239 
rect 50 239 51 240 
rect 50 240 51 241 
rect 50 241 51 242 
rect 50 244 51 245 
rect 50 257 51 258 
rect 50 261 51 262 
rect 50 273 51 274 
rect 50 289 51 290 
rect 50 292 51 293 
rect 50 305 51 306 
rect 50 307 51 308 
rect 51 2 52 3 
rect 51 3 52 4 
rect 51 8 52 9 
rect 51 18 52 19 
rect 51 50 52 51 
rect 51 51 52 52 
rect 51 52 52 53 
rect 51 53 52 54 
rect 51 54 52 55 
rect 51 55 52 56 
rect 51 82 52 83 
rect 51 100 52 101 
rect 51 103 52 104 
rect 51 105 52 106 
rect 51 106 52 107 
rect 51 107 52 108 
rect 51 108 52 109 
rect 51 109 52 110 
rect 51 110 52 111 
rect 51 111 52 112 
rect 51 112 52 113 
rect 51 113 52 114 
rect 51 114 52 115 
rect 51 115 52 116 
rect 51 116 52 117 
rect 51 117 52 118 
rect 51 118 52 119 
rect 51 119 52 120 
rect 51 120 52 121 
rect 51 121 52 122 
rect 51 122 52 123 
rect 51 123 52 124 
rect 51 124 52 125 
rect 51 125 52 126 
rect 51 126 52 127 
rect 51 127 52 128 
rect 51 128 52 129 
rect 51 129 52 130 
rect 51 130 52 131 
rect 51 131 52 132 
rect 51 132 52 133 
rect 51 133 52 134 
rect 51 134 52 135 
rect 51 135 52 136 
rect 51 136 52 137 
rect 51 137 52 138 
rect 51 138 52 139 
rect 51 139 52 140 
rect 51 140 52 141 
rect 51 141 52 142 
rect 51 142 52 143 
rect 51 143 52 144 
rect 51 144 52 145 
rect 51 145 52 146 
rect 51 146 52 147 
rect 51 147 52 148 
rect 51 148 52 149 
rect 51 149 52 150 
rect 51 150 52 151 
rect 51 151 52 152 
rect 51 152 52 153 
rect 51 153 52 154 
rect 51 154 52 155 
rect 51 155 52 156 
rect 51 156 52 157 
rect 51 157 52 158 
rect 51 158 52 159 
rect 51 159 52 160 
rect 51 160 52 161 
rect 51 163 52 164 
rect 51 165 52 166 
rect 51 166 52 167 
rect 51 167 52 168 
rect 51 168 52 169 
rect 51 169 52 170 
rect 51 170 52 171 
rect 51 171 52 172 
rect 51 172 52 173 
rect 51 173 52 174 
rect 51 174 52 175 
rect 51 175 52 176 
rect 51 176 52 177 
rect 51 177 52 178 
rect 51 178 52 179 
rect 51 179 52 180 
rect 51 180 52 181 
rect 51 181 52 182 
rect 51 182 52 183 
rect 51 183 52 184 
rect 51 184 52 185 
rect 51 185 52 186 
rect 51 186 52 187 
rect 51 187 52 188 
rect 51 188 52 189 
rect 51 189 52 190 
rect 51 190 52 191 
rect 51 191 52 192 
rect 51 192 52 193 
rect 51 193 52 194 
rect 51 194 52 195 
rect 51 195 52 196 
rect 51 196 52 197 
rect 51 197 52 198 
rect 51 198 52 199 
rect 51 199 52 200 
rect 51 200 52 201 
rect 51 201 52 202 
rect 51 202 52 203 
rect 51 203 52 204 
rect 51 204 52 205 
rect 51 205 52 206 
rect 51 206 52 207 
rect 51 207 52 208 
rect 51 208 52 209 
rect 51 209 52 210 
rect 51 210 52 211 
rect 51 232 52 233 
rect 51 241 52 242 
rect 51 244 52 245 
rect 51 257 52 258 
rect 51 261 52 262 
rect 51 273 52 274 
rect 51 289 52 290 
rect 51 292 52 293 
rect 51 305 52 306 
rect 51 307 52 308 
rect 52 2 53 3 
rect 52 8 53 9 
rect 52 18 53 19 
rect 52 55 53 56 
rect 52 82 53 83 
rect 52 103 53 104 
rect 52 163 53 164 
rect 52 232 53 233 
rect 52 241 53 242 
rect 52 244 53 245 
rect 52 257 53 258 
rect 52 261 53 262 
rect 52 273 53 274 
rect 52 289 53 290 
rect 52 292 53 293 
rect 52 305 53 306 
rect 52 307 53 308 
rect 53 2 54 3 
rect 53 8 54 9 
rect 53 18 54 19 
rect 53 55 54 56 
rect 53 80 54 81 
rect 53 82 54 83 
rect 53 103 54 104 
rect 53 152 54 153 
rect 53 163 54 164 
rect 53 196 54 197 
rect 53 197 54 198 
rect 53 198 54 199 
rect 53 199 54 200 
rect 53 232 54 233 
rect 53 241 54 242 
rect 53 244 54 245 
rect 53 257 54 258 
rect 53 261 54 262 
rect 53 273 54 274 
rect 53 289 54 290 
rect 53 292 54 293 
rect 53 305 54 306 
rect 53 307 54 308 
rect 54 2 55 3 
rect 54 8 55 9 
rect 54 18 55 19 
rect 54 55 55 56 
rect 54 77 55 78 
rect 54 78 55 79 
rect 54 79 55 80 
rect 54 80 55 81 
rect 54 82 55 83 
rect 54 103 55 104 
rect 54 130 55 131 
rect 54 131 55 132 
rect 54 132 55 133 
rect 54 133 55 134 
rect 54 134 55 135 
rect 54 135 55 136 
rect 54 136 55 137 
rect 54 137 55 138 
rect 54 138 55 139 
rect 54 139 55 140 
rect 54 140 55 141 
rect 54 141 55 142 
rect 54 142 55 143 
rect 54 143 55 144 
rect 54 144 55 145 
rect 54 145 55 146 
rect 54 146 55 147 
rect 54 147 55 148 
rect 54 148 55 149 
rect 54 149 55 150 
rect 54 150 55 151 
rect 54 151 55 152 
rect 54 152 55 153 
rect 54 163 55 164 
rect 54 165 55 166 
rect 54 166 55 167 
rect 54 167 55 168 
rect 54 168 55 169 
rect 54 169 55 170 
rect 54 170 55 171 
rect 54 171 55 172 
rect 54 172 55 173 
rect 54 173 55 174 
rect 54 174 55 175 
rect 54 175 55 176 
rect 54 176 55 177 
rect 54 177 55 178 
rect 54 178 55 179 
rect 54 179 55 180 
rect 54 180 55 181 
rect 54 181 55 182 
rect 54 182 55 183 
rect 54 183 55 184 
rect 54 184 55 185 
rect 54 185 55 186 
rect 54 186 55 187 
rect 54 187 55 188 
rect 54 188 55 189 
rect 54 189 55 190 
rect 54 190 55 191 
rect 54 191 55 192 
rect 54 199 55 200 
rect 54 200 55 201 
rect 54 201 55 202 
rect 54 202 55 203 
rect 54 203 55 204 
rect 54 204 55 205 
rect 54 205 55 206 
rect 54 206 55 207 
rect 54 207 55 208 
rect 54 208 55 209 
rect 54 209 55 210 
rect 54 210 55 211 
rect 54 211 55 212 
rect 54 212 55 213 
rect 54 213 55 214 
rect 54 214 55 215 
rect 54 215 55 216 
rect 54 216 55 217 
rect 54 217 55 218 
rect 54 218 55 219 
rect 54 219 55 220 
rect 54 220 55 221 
rect 54 221 55 222 
rect 54 222 55 223 
rect 54 223 55 224 
rect 54 224 55 225 
rect 54 225 55 226 
rect 54 226 55 227 
rect 54 227 55 228 
rect 54 228 55 229 
rect 54 229 55 230 
rect 54 230 55 231 
rect 54 232 55 233 
rect 54 241 55 242 
rect 54 244 55 245 
rect 54 257 55 258 
rect 54 261 55 262 
rect 54 273 55 274 
rect 54 289 55 290 
rect 54 292 55 293 
rect 54 305 55 306 
rect 54 307 55 308 
rect 55 2 56 3 
rect 55 8 56 9 
rect 55 18 56 19 
rect 55 55 56 56 
rect 55 76 56 77 
rect 55 77 56 78 
rect 55 82 56 83 
rect 55 103 56 104 
rect 55 153 56 154 
rect 55 154 56 155 
rect 55 155 56 156 
rect 55 156 56 157 
rect 55 157 56 158 
rect 55 158 56 159 
rect 55 159 56 160 
rect 55 163 56 164 
rect 55 191 56 192 
rect 55 192 56 193 
rect 55 193 56 194 
rect 55 194 56 195 
rect 55 195 56 196 
rect 55 232 56 233 
rect 55 241 56 242 
rect 55 244 56 245 
rect 55 246 56 247 
rect 55 257 56 258 
rect 55 261 56 262 
rect 55 263 56 264 
rect 55 264 56 265 
rect 55 265 56 266 
rect 55 266 56 267 
rect 55 267 56 268 
rect 55 268 56 269 
rect 55 269 56 270 
rect 55 273 56 274 
rect 55 289 56 290 
rect 55 292 56 293 
rect 55 305 56 306 
rect 55 307 56 308 
rect 56 2 57 3 
rect 56 8 57 9 
rect 56 18 57 19 
rect 56 55 57 56 
rect 56 57 57 58 
rect 56 58 57 59 
rect 56 59 57 60 
rect 56 60 57 61 
rect 56 61 57 62 
rect 56 62 57 63 
rect 56 63 57 64 
rect 56 64 57 65 
rect 56 65 57 66 
rect 56 66 57 67 
rect 56 67 57 68 
rect 56 68 57 69 
rect 56 69 57 70 
rect 56 70 57 71 
rect 56 71 57 72 
rect 56 72 57 73 
rect 56 73 57 74 
rect 56 74 57 75 
rect 56 75 57 76 
rect 56 76 57 77 
rect 56 78 57 79 
rect 56 79 57 80 
rect 56 80 57 81 
rect 56 82 57 83 
rect 56 103 57 104 
rect 56 105 57 106 
rect 56 106 57 107 
rect 56 107 57 108 
rect 56 108 57 109 
rect 56 109 57 110 
rect 56 110 57 111 
rect 56 111 57 112 
rect 56 112 57 113 
rect 56 113 57 114 
rect 56 114 57 115 
rect 56 115 57 116 
rect 56 116 57 117 
rect 56 117 57 118 
rect 56 118 57 119 
rect 56 119 57 120 
rect 56 120 57 121 
rect 56 121 57 122 
rect 56 122 57 123 
rect 56 123 57 124 
rect 56 124 57 125 
rect 56 125 57 126 
rect 56 126 57 127 
rect 56 127 57 128 
rect 56 128 57 129 
rect 56 129 57 130 
rect 56 130 57 131 
rect 56 131 57 132 
rect 56 132 57 133 
rect 56 133 57 134 
rect 56 134 57 135 
rect 56 135 57 136 
rect 56 136 57 137 
rect 56 137 57 138 
rect 56 138 57 139 
rect 56 139 57 140 
rect 56 140 57 141 
rect 56 141 57 142 
rect 56 142 57 143 
rect 56 143 57 144 
rect 56 144 57 145 
rect 56 145 57 146 
rect 56 146 57 147 
rect 56 147 57 148 
rect 56 148 57 149 
rect 56 149 57 150 
rect 56 150 57 151 
rect 56 151 57 152 
rect 56 152 57 153 
rect 56 153 57 154 
rect 56 159 57 160 
rect 56 160 57 161 
rect 56 163 57 164 
rect 56 165 57 166 
rect 56 166 57 167 
rect 56 167 57 168 
rect 56 168 57 169 
rect 56 169 57 170 
rect 56 170 57 171 
rect 56 171 57 172 
rect 56 172 57 173 
rect 56 173 57 174 
rect 56 174 57 175 
rect 56 175 57 176 
rect 56 176 57 177 
rect 56 177 57 178 
rect 56 178 57 179 
rect 56 179 57 180 
rect 56 180 57 181 
rect 56 181 57 182 
rect 56 182 57 183 
rect 56 183 57 184 
rect 56 184 57 185 
rect 56 185 57 186 
rect 56 186 57 187 
rect 56 187 57 188 
rect 56 188 57 189 
rect 56 189 57 190 
rect 56 190 57 191 
rect 56 195 57 196 
rect 56 196 57 197 
rect 56 197 57 198 
rect 56 198 57 199 
rect 56 199 57 200 
rect 56 200 57 201 
rect 56 201 57 202 
rect 56 202 57 203 
rect 56 203 57 204 
rect 56 204 57 205 
rect 56 205 57 206 
rect 56 206 57 207 
rect 56 207 57 208 
rect 56 208 57 209 
rect 56 209 57 210 
rect 56 210 57 211 
rect 56 211 57 212 
rect 56 212 57 213 
rect 56 213 57 214 
rect 56 214 57 215 
rect 56 215 57 216 
rect 56 216 57 217 
rect 56 217 57 218 
rect 56 218 57 219 
rect 56 219 57 220 
rect 56 220 57 221 
rect 56 221 57 222 
rect 56 222 57 223 
rect 56 223 57 224 
rect 56 224 57 225 
rect 56 232 57 233 
rect 56 235 57 236 
rect 56 241 57 242 
rect 56 244 57 245 
rect 56 246 57 247 
rect 56 247 57 248 
rect 56 248 57 249 
rect 56 249 57 250 
rect 56 250 57 251 
rect 56 251 57 252 
rect 56 257 57 258 
rect 56 261 57 262 
rect 56 263 57 264 
rect 56 269 57 270 
rect 56 270 57 271 
rect 56 273 57 274 
rect 56 275 57 276 
rect 56 276 57 277 
rect 56 277 57 278 
rect 56 278 57 279 
rect 56 279 57 280 
rect 56 280 57 281 
rect 56 281 57 282 
rect 56 282 57 283 
rect 56 283 57 284 
rect 56 284 57 285 
rect 56 285 57 286 
rect 56 286 57 287 
rect 56 289 57 290 
rect 56 292 57 293 
rect 56 302 57 303 
rect 56 305 57 306 
rect 56 307 57 308 
rect 57 2 58 3 
rect 57 8 58 9 
rect 57 18 58 19 
rect 57 55 58 56 
rect 57 57 58 58 
rect 57 78 58 79 
rect 57 80 58 81 
rect 57 82 58 83 
rect 57 104 58 105 
rect 57 105 58 106 
rect 57 163 58 164 
rect 57 190 58 191 
rect 57 224 58 225 
rect 57 225 58 226 
rect 57 232 58 233 
rect 57 235 58 236 
rect 57 241 58 242 
rect 57 244 58 245 
rect 57 251 58 252 
rect 57 257 58 258 
rect 57 263 58 264 
rect 57 273 58 274 
rect 57 286 58 287 
rect 57 289 58 290 
rect 57 292 58 293 
rect 57 302 58 303 
rect 57 305 58 306 
rect 57 307 58 308 
rect 57 309 58 310 
rect 58 2 59 3 
rect 58 8 59 9 
rect 58 18 59 19 
rect 58 55 59 56 
rect 58 78 59 79 
rect 58 82 59 83 
rect 58 98 59 99 
rect 58 99 59 100 
rect 58 100 59 101 
rect 58 101 59 102 
rect 58 102 59 103 
rect 58 103 59 104 
rect 58 104 59 105 
rect 58 163 59 164 
rect 58 190 59 191 
rect 58 225 59 226 
rect 58 232 59 233 
rect 58 235 59 236 
rect 58 241 59 242 
rect 58 244 59 245 
rect 58 251 59 252 
rect 58 257 59 258 
rect 58 259 59 260 
rect 58 260 59 261 
rect 58 261 59 262 
rect 58 262 59 263 
rect 58 263 59 264 
rect 58 273 59 274 
rect 58 286 59 287 
rect 58 289 59 290 
rect 58 292 59 293 
rect 58 302 59 303 
rect 58 305 59 306 
rect 58 307 59 308 
rect 58 309 59 310 
rect 59 2 60 3 
rect 59 8 60 9 
rect 59 18 60 19 
rect 59 55 60 56 
rect 59 82 60 83 
rect 59 98 60 99 
rect 59 163 60 164 
rect 59 225 60 226 
rect 59 232 60 233 
rect 59 241 60 242 
rect 59 244 60 245 
rect 59 257 60 258 
rect 59 259 60 260 
rect 59 273 60 274 
rect 59 289 60 290 
rect 59 292 60 293 
rect 59 305 60 306 
rect 59 307 60 308 
rect 59 309 60 310 
rect 60 2 61 3 
rect 60 8 61 9 
rect 60 18 61 19 
rect 60 55 61 56 
rect 60 82 61 83 
rect 60 98 61 99 
rect 60 163 61 164 
rect 60 225 61 226 
rect 60 232 61 233 
rect 60 241 61 242 
rect 60 244 61 245 
rect 60 257 61 258 
rect 60 259 61 260 
rect 60 273 61 274 
rect 60 289 61 290 
rect 60 292 61 293 
rect 60 305 61 306 
rect 60 307 61 308 
rect 60 309 61 310 
rect 61 2 62 3 
rect 61 8 62 9 
rect 61 18 62 19 
rect 61 51 62 52 
rect 61 55 62 56 
rect 61 82 62 83 
rect 61 98 62 99 
rect 61 163 62 164 
rect 61 225 62 226 
rect 61 232 62 233 
rect 61 241 62 242 
rect 61 244 62 245 
rect 61 257 62 258 
rect 61 259 62 260 
rect 61 273 62 274 
rect 61 274 62 275 
rect 61 275 62 276 
rect 61 289 62 290 
rect 61 292 62 293 
rect 61 305 62 306 
rect 61 307 62 308 
rect 61 309 62 310 
rect 61 310 62 311 
rect 62 2 63 3 
rect 62 8 63 9 
rect 62 18 63 19 
rect 62 51 63 52 
rect 62 55 63 56 
rect 62 82 63 83 
rect 62 98 63 99 
rect 62 163 63 164 
rect 62 225 63 226 
rect 62 232 63 233 
rect 62 241 63 242 
rect 62 244 63 245 
rect 62 257 63 258 
rect 62 259 63 260 
rect 62 275 63 276 
rect 62 289 63 290 
rect 62 292 63 293 
rect 62 305 63 306 
rect 62 307 63 308 
rect 62 310 63 311 
rect 63 2 64 3 
rect 63 8 64 9 
rect 63 18 64 19 
rect 63 43 64 44 
rect 63 51 64 52 
rect 63 55 64 56 
rect 63 62 64 63 
rect 63 82 64 83 
rect 63 98 64 99 
rect 63 139 64 140 
rect 63 163 64 164 
rect 63 232 64 233 
rect 63 241 64 242 
rect 63 244 64 245 
rect 63 257 64 258 
rect 63 259 64 260 
rect 63 275 64 276 
rect 63 289 64 290 
rect 63 292 64 293 
rect 63 305 64 306 
rect 63 307 64 308 
rect 63 310 64 311 
rect 64 2 65 3 
rect 64 8 65 9 
rect 64 18 65 19 
rect 64 43 65 44 
rect 64 51 65 52 
rect 64 55 65 56 
rect 64 62 65 63 
rect 64 82 65 83 
rect 64 139 65 140 
rect 64 232 65 233 
rect 64 241 65 242 
rect 64 244 65 245 
rect 64 257 65 258 
rect 64 259 65 260 
rect 64 275 65 276 
rect 64 289 65 290 
rect 64 292 65 293 
rect 64 305 65 306 
rect 64 307 65 308 
rect 64 310 65 311 
rect 65 2 66 3 
rect 65 8 66 9 
rect 65 14 66 15 
rect 65 15 66 16 
rect 65 16 66 17 
rect 65 17 66 18 
rect 65 18 66 19 
rect 65 27 66 28 
rect 65 28 66 29 
rect 65 29 66 30 
rect 65 30 66 31 
rect 65 31 66 32 
rect 65 32 66 33 
rect 65 33 66 34 
rect 65 34 66 35 
rect 65 35 66 36 
rect 65 36 66 37 
rect 65 37 66 38 
rect 65 38 66 39 
rect 65 39 66 40 
rect 65 40 66 41 
rect 65 41 66 42 
rect 65 42 66 43 
rect 65 43 66 44 
rect 65 51 66 52 
rect 65 55 66 56 
rect 65 56 66 57 
rect 65 57 66 58 
rect 65 58 66 59 
rect 65 59 66 60 
rect 65 60 66 61 
rect 65 62 66 63 
rect 65 63 66 64 
rect 65 64 66 65 
rect 65 65 66 66 
rect 65 66 66 67 
rect 65 67 66 68 
rect 65 68 66 69 
rect 65 69 66 70 
rect 65 70 66 71 
rect 65 71 66 72 
rect 65 72 66 73 
rect 65 73 66 74 
rect 65 75 66 76 
rect 65 76 66 77 
rect 65 77 66 78 
rect 65 78 66 79 
rect 65 79 66 80 
rect 65 80 66 81 
rect 65 81 66 82 
rect 65 82 66 83 
rect 65 85 66 86 
rect 65 86 66 87 
rect 65 87 66 88 
rect 65 88 66 89 
rect 65 89 66 90 
rect 65 90 66 91 
rect 65 91 66 92 
rect 65 92 66 93 
rect 65 93 66 94 
rect 65 94 66 95 
rect 65 95 66 96 
rect 65 96 66 97 
rect 65 97 66 98 
rect 65 98 66 99 
rect 65 99 66 100 
rect 65 100 66 101 
rect 65 101 66 102 
rect 65 102 66 103 
rect 65 103 66 104 
rect 65 104 66 105 
rect 65 105 66 106 
rect 65 106 66 107 
rect 65 107 66 108 
rect 65 108 66 109 
rect 65 109 66 110 
rect 65 110 66 111 
rect 65 111 66 112 
rect 65 112 66 113 
rect 65 113 66 114 
rect 65 114 66 115 
rect 65 115 66 116 
rect 65 116 66 117 
rect 65 117 66 118 
rect 65 118 66 119 
rect 65 119 66 120 
rect 65 120 66 121 
rect 65 121 66 122 
rect 65 122 66 123 
rect 65 123 66 124 
rect 65 124 66 125 
rect 65 125 66 126 
rect 65 126 66 127 
rect 65 127 66 128 
rect 65 128 66 129 
rect 65 129 66 130 
rect 65 130 66 131 
rect 65 131 66 132 
rect 65 132 66 133 
rect 65 133 66 134 
rect 65 134 66 135 
rect 65 135 66 136 
rect 65 136 66 137 
rect 65 137 66 138 
rect 65 139 66 140 
rect 65 140 66 141 
rect 65 141 66 142 
rect 65 142 66 143 
rect 65 143 66 144 
rect 65 144 66 145 
rect 65 145 66 146 
rect 65 146 66 147 
rect 65 147 66 148 
rect 65 148 66 149 
rect 65 149 66 150 
rect 65 150 66 151 
rect 65 151 66 152 
rect 65 152 66 153 
rect 65 153 66 154 
rect 65 154 66 155 
rect 65 155 66 156 
rect 65 156 66 157 
rect 65 157 66 158 
rect 65 158 66 159 
rect 65 159 66 160 
rect 65 160 66 161 
rect 65 161 66 162 
rect 65 162 66 163 
rect 65 163 66 164 
rect 65 164 66 165 
rect 65 165 66 166 
rect 65 166 66 167 
rect 65 167 66 168 
rect 65 168 66 169 
rect 65 169 66 170 
rect 65 170 66 171 
rect 65 171 66 172 
rect 65 172 66 173 
rect 65 173 66 174 
rect 65 174 66 175 
rect 65 175 66 176 
rect 65 176 66 177 
rect 65 177 66 178 
rect 65 178 66 179 
rect 65 179 66 180 
rect 65 180 66 181 
rect 65 181 66 182 
rect 65 182 66 183 
rect 65 183 66 184 
rect 65 184 66 185 
rect 65 185 66 186 
rect 65 186 66 187 
rect 65 187 66 188 
rect 65 188 66 189 
rect 65 189 66 190 
rect 65 190 66 191 
rect 65 191 66 192 
rect 65 192 66 193 
rect 65 193 66 194 
rect 65 194 66 195 
rect 65 195 66 196 
rect 65 196 66 197 
rect 65 197 66 198 
rect 65 198 66 199 
rect 65 199 66 200 
rect 65 200 66 201 
rect 65 201 66 202 
rect 65 202 66 203 
rect 65 203 66 204 
rect 65 204 66 205 
rect 65 205 66 206 
rect 65 206 66 207 
rect 65 207 66 208 
rect 65 208 66 209 
rect 65 209 66 210 
rect 65 210 66 211 
rect 65 211 66 212 
rect 65 212 66 213 
rect 65 213 66 214 
rect 65 214 66 215 
rect 65 215 66 216 
rect 65 216 66 217 
rect 65 217 66 218 
rect 65 218 66 219 
rect 65 219 66 220 
rect 65 220 66 221 
rect 65 221 66 222 
rect 65 222 66 223 
rect 65 223 66 224 
rect 65 224 66 225 
rect 65 225 66 226 
rect 65 226 66 227 
rect 65 227 66 228 
rect 65 228 66 229 
rect 65 229 66 230 
rect 65 230 66 231 
rect 65 231 66 232 
rect 65 232 66 233 
rect 65 241 66 242 
rect 65 243 66 244 
rect 65 244 66 245 
rect 65 257 66 258 
rect 65 259 66 260 
rect 65 275 66 276 
rect 65 289 66 290 
rect 65 292 66 293 
rect 65 305 66 306 
rect 65 307 66 308 
rect 65 310 66 311 
rect 66 2 67 3 
rect 66 8 67 9 
rect 66 14 67 15 
rect 66 27 67 28 
rect 66 51 67 52 
rect 66 60 67 61 
rect 66 61 67 62 
rect 66 75 67 76 
rect 66 137 67 138 
rect 66 138 67 139 
rect 66 239 67 240 
rect 66 241 67 242 
rect 66 243 67 244 
rect 66 257 67 258 
rect 66 259 67 260 
rect 66 275 67 276 
rect 66 289 67 290 
rect 66 292 67 293 
rect 66 305 67 306 
rect 66 307 67 308 
rect 66 310 67 311 
rect 67 2 68 3 
rect 67 8 68 9 
rect 67 14 68 15 
rect 67 27 68 28 
rect 67 51 68 52 
rect 67 61 68 62 
rect 67 62 68 63 
rect 67 63 68 64 
rect 67 64 68 65 
rect 67 65 68 66 
rect 67 75 68 76 
rect 67 90 68 91 
rect 67 91 68 92 
rect 67 92 68 93 
rect 67 93 68 94 
rect 67 94 68 95 
rect 67 95 68 96 
rect 67 96 68 97 
rect 67 138 68 139 
rect 67 139 68 140 
rect 67 140 68 141 
rect 67 141 68 142 
rect 67 142 68 143 
rect 67 143 68 144 
rect 67 144 68 145 
rect 67 145 68 146 
rect 67 146 68 147 
rect 67 147 68 148 
rect 67 148 68 149 
rect 67 149 68 150 
rect 67 150 68 151 
rect 67 151 68 152 
rect 67 152 68 153 
rect 67 153 68 154 
rect 67 154 68 155 
rect 67 155 68 156 
rect 67 156 68 157 
rect 67 157 68 158 
rect 67 158 68 159 
rect 67 159 68 160 
rect 67 160 68 161 
rect 67 161 68 162 
rect 67 162 68 163 
rect 67 163 68 164 
rect 67 164 68 165 
rect 67 165 68 166 
rect 67 198 68 199 
rect 67 199 68 200 
rect 67 200 68 201 
rect 67 201 68 202 
rect 67 202 68 203 
rect 67 203 68 204 
rect 67 204 68 205 
rect 67 205 68 206 
rect 67 206 68 207 
rect 67 207 68 208 
rect 67 208 68 209 
rect 67 209 68 210 
rect 67 210 68 211 
rect 67 213 68 214 
rect 67 214 68 215 
rect 67 215 68 216 
rect 67 216 68 217 
rect 67 217 68 218 
rect 67 218 68 219 
rect 67 219 68 220 
rect 67 220 68 221 
rect 67 221 68 222 
rect 67 222 68 223 
rect 67 223 68 224 
rect 67 224 68 225 
rect 67 225 68 226 
rect 67 226 68 227 
rect 67 227 68 228 
rect 67 228 68 229 
rect 67 229 68 230 
rect 67 230 68 231 
rect 67 231 68 232 
rect 67 232 68 233 
rect 67 233 68 234 
rect 67 234 68 235 
rect 67 235 68 236 
rect 67 236 68 237 
rect 67 237 68 238 
rect 67 238 68 239 
rect 67 239 68 240 
rect 67 241 68 242 
rect 67 243 68 244 
rect 67 245 68 246 
rect 67 257 68 258 
rect 67 259 68 260 
rect 67 275 68 276 
rect 67 289 68 290 
rect 67 292 68 293 
rect 67 305 68 306 
rect 67 307 68 308 
rect 67 310 68 311 
rect 68 2 69 3 
rect 68 8 69 9 
rect 68 14 69 15 
rect 68 27 69 28 
rect 68 51 69 52 
rect 68 65 69 66 
rect 68 75 69 76 
rect 68 89 69 90 
rect 68 90 69 91 
rect 68 96 69 97 
rect 68 97 69 98 
rect 68 98 69 99 
rect 68 99 69 100 
rect 68 100 69 101 
rect 68 101 69 102 
rect 68 102 69 103 
rect 68 103 69 104 
rect 68 104 69 105 
rect 68 105 69 106 
rect 68 106 69 107 
rect 68 107 69 108 
rect 68 108 69 109 
rect 68 109 69 110 
rect 68 110 69 111 
rect 68 111 69 112 
rect 68 112 69 113 
rect 68 113 69 114 
rect 68 114 69 115 
rect 68 115 69 116 
rect 68 116 69 117 
rect 68 117 69 118 
rect 68 118 69 119 
rect 68 119 69 120 
rect 68 120 69 121 
rect 68 121 69 122 
rect 68 122 69 123 
rect 68 123 69 124 
rect 68 124 69 125 
rect 68 125 69 126 
rect 68 126 69 127 
rect 68 127 69 128 
rect 68 128 69 129 
rect 68 129 69 130 
rect 68 130 69 131 
rect 68 131 69 132 
rect 68 165 69 166 
rect 68 168 69 169 
rect 68 241 69 242 
rect 68 243 69 244 
rect 68 245 69 246 
rect 68 257 69 258 
rect 68 259 69 260 
rect 68 275 69 276 
rect 68 289 69 290 
rect 68 292 69 293 
rect 68 305 69 306 
rect 68 307 69 308 
rect 68 310 69 311 
rect 69 2 70 3 
rect 69 8 70 9 
rect 69 14 70 15 
rect 69 27 70 28 
rect 69 42 70 43 
rect 69 43 70 44 
rect 69 44 70 45 
rect 69 45 70 46 
rect 69 46 70 47 
rect 69 47 70 48 
rect 69 48 70 49 
rect 69 49 70 50 
rect 69 50 70 51 
rect 69 51 70 52 
rect 69 165 70 166 
rect 69 168 70 169 
rect 69 169 70 170 
rect 69 170 70 171 
rect 69 171 70 172 
rect 69 172 70 173 
rect 69 173 70 174 
rect 69 174 70 175 
rect 69 175 70 176 
rect 69 176 70 177 
rect 69 177 70 178 
rect 69 178 70 179 
rect 69 179 70 180 
rect 69 180 70 181 
rect 69 181 70 182 
rect 69 182 70 183 
rect 69 183 70 184 
rect 69 184 70 185 
rect 69 185 70 186 
rect 69 186 70 187 
rect 69 187 70 188 
rect 69 188 70 189 
rect 69 189 70 190 
rect 69 190 70 191 
rect 69 191 70 192 
rect 69 192 70 193 
rect 69 193 70 194 
rect 69 194 70 195 
rect 69 195 70 196 
rect 69 196 70 197 
rect 69 197 70 198 
rect 69 198 70 199 
rect 69 199 70 200 
rect 69 200 70 201 
rect 69 201 70 202 
rect 69 202 70 203 
rect 69 203 70 204 
rect 69 204 70 205 
rect 69 205 70 206 
rect 69 206 70 207 
rect 69 207 70 208 
rect 69 208 70 209 
rect 69 209 70 210 
rect 69 210 70 211 
rect 69 211 70 212 
rect 69 212 70 213 
rect 69 213 70 214 
rect 69 214 70 215 
rect 69 215 70 216 
rect 69 216 70 217 
rect 69 241 70 242 
rect 69 243 70 244 
rect 69 245 70 246 
rect 69 257 70 258 
rect 69 275 70 276 
rect 69 289 70 290 
rect 69 292 70 293 
rect 69 305 70 306 
rect 69 307 70 308 
rect 69 310 70 311 
rect 70 2 71 3 
rect 70 8 71 9 
rect 70 13 71 14 
rect 70 14 71 15 
rect 70 27 71 28 
rect 70 40 71 41 
rect 70 41 71 42 
rect 70 42 71 43 
rect 70 58 71 59 
rect 70 59 71 60 
rect 70 60 71 61 
rect 70 61 71 62 
rect 70 62 71 63 
rect 70 63 71 64 
rect 70 64 71 65 
rect 70 65 71 66 
rect 70 66 71 67 
rect 70 67 71 68 
rect 70 68 71 69 
rect 70 69 71 70 
rect 70 70 71 71 
rect 70 71 71 72 
rect 70 72 71 73 
rect 70 73 71 74 
rect 70 74 71 75 
rect 70 75 71 76 
rect 70 76 71 77 
rect 70 77 71 78 
rect 70 78 71 79 
rect 70 79 71 80 
rect 70 80 71 81 
rect 70 81 71 82 
rect 70 82 71 83 
rect 70 83 71 84 
rect 70 84 71 85 
rect 70 85 71 86 
rect 70 86 71 87 
rect 70 87 71 88 
rect 70 88 71 89 
rect 70 89 71 90 
rect 70 90 71 91 
rect 70 91 71 92 
rect 70 92 71 93 
rect 70 93 71 94 
rect 70 94 71 95 
rect 70 95 71 96 
rect 70 96 71 97 
rect 70 97 71 98 
rect 70 98 71 99 
rect 70 99 71 100 
rect 70 100 71 101 
rect 70 101 71 102 
rect 70 102 71 103 
rect 70 103 71 104 
rect 70 104 71 105 
rect 70 105 71 106 
rect 70 106 71 107 
rect 70 107 71 108 
rect 70 108 71 109 
rect 70 109 71 110 
rect 70 110 71 111 
rect 70 111 71 112 
rect 70 112 71 113 
rect 70 113 71 114 
rect 70 114 71 115 
rect 70 115 71 116 
rect 70 116 71 117 
rect 70 117 71 118 
rect 70 118 71 119 
rect 70 119 71 120 
rect 70 120 71 121 
rect 70 121 71 122 
rect 70 122 71 123 
rect 70 123 71 124 
rect 70 124 71 125 
rect 70 125 71 126 
rect 70 126 71 127 
rect 70 127 71 128 
rect 70 128 71 129 
rect 70 129 71 130 
rect 70 130 71 131 
rect 70 131 71 132 
rect 70 132 71 133 
rect 70 133 71 134 
rect 70 134 71 135 
rect 70 135 71 136 
rect 70 136 71 137 
rect 70 137 71 138 
rect 70 138 71 139 
rect 70 139 71 140 
rect 70 140 71 141 
rect 70 141 71 142 
rect 70 142 71 143 
rect 70 143 71 144 
rect 70 144 71 145 
rect 70 145 71 146 
rect 70 146 71 147 
rect 70 147 71 148 
rect 70 148 71 149 
rect 70 149 71 150 
rect 70 150 71 151 
rect 70 151 71 152 
rect 70 152 71 153 
rect 70 153 71 154 
rect 70 154 71 155 
rect 70 155 71 156 
rect 70 156 71 157 
rect 70 157 71 158 
rect 70 158 71 159 
rect 70 159 71 160 
rect 70 160 71 161 
rect 70 161 71 162 
rect 70 165 71 166 
rect 70 216 71 217 
rect 70 218 71 219 
rect 70 219 71 220 
rect 70 220 71 221 
rect 70 221 71 222 
rect 70 222 71 223 
rect 70 223 71 224 
rect 70 224 71 225 
rect 70 225 71 226 
rect 70 226 71 227 
rect 70 227 71 228 
rect 70 241 71 242 
rect 70 243 71 244 
rect 70 245 71 246 
rect 70 275 71 276 
rect 70 289 71 290 
rect 70 292 71 293 
rect 70 305 71 306 
rect 70 307 71 308 
rect 70 310 71 311 
rect 71 1 72 2 
rect 71 2 72 3 
rect 71 7 72 8 
rect 71 8 72 9 
rect 71 12 72 13 
rect 71 13 72 14 
rect 71 27 72 28 
rect 71 39 72 40 
rect 71 40 72 41 
rect 71 57 72 58 
rect 71 58 72 59 
rect 71 161 72 162 
rect 71 162 72 163 
rect 71 289 72 290 
rect 71 292 72 293 
rect 71 305 72 306 
rect 71 307 72 308 
rect 71 310 72 311 
rect 72 1 73 2 
rect 72 3 73 4 
rect 72 4 73 5 
rect 72 5 73 6 
rect 72 6 73 7 
rect 72 7 73 8 
rect 72 9 73 10 
rect 72 10 73 11 
rect 72 11 73 12 
rect 72 12 73 13 
rect 72 14 73 15 
rect 72 15 73 16 
rect 72 16 73 17 
rect 72 27 73 28 
rect 72 39 73 40 
rect 72 41 73 42 
rect 72 42 73 43 
rect 72 43 73 44 
rect 72 44 73 45 
rect 72 45 73 46 
rect 72 46 73 47 
rect 72 47 73 48 
rect 72 48 73 49 
rect 72 49 73 50 
rect 72 50 73 51 
rect 72 51 73 52 
rect 72 52 73 53 
rect 72 53 73 54 
rect 72 54 73 55 
rect 72 55 73 56 
rect 72 56 73 57 
rect 72 57 73 58 
rect 72 59 73 60 
rect 72 60 73 61 
rect 72 61 73 62 
rect 72 62 73 63 
rect 72 63 73 64 
rect 72 64 73 65 
rect 72 65 73 66 
rect 72 66 73 67 
rect 72 67 73 68 
rect 72 68 73 69 
rect 72 69 73 70 
rect 72 70 73 71 
rect 72 71 73 72 
rect 72 72 73 73 
rect 72 73 73 74 
rect 72 74 73 75 
rect 72 75 73 76 
rect 72 76 73 77 
rect 72 77 73 78 
rect 72 78 73 79 
rect 72 79 73 80 
rect 72 80 73 81 
rect 72 81 73 82 
rect 72 82 73 83 
rect 72 83 73 84 
rect 72 84 73 85 
rect 72 85 73 86 
rect 72 86 73 87 
rect 72 87 73 88 
rect 72 88 73 89 
rect 72 89 73 90 
rect 72 90 73 91 
rect 72 91 73 92 
rect 72 92 73 93 
rect 72 93 73 94 
rect 72 94 73 95 
rect 72 95 73 96 
rect 72 96 73 97 
rect 72 97 73 98 
rect 72 98 73 99 
rect 72 99 73 100 
rect 72 100 73 101 
rect 72 101 73 102 
rect 72 102 73 103 
rect 72 103 73 104 
rect 72 104 73 105 
rect 72 105 73 106 
rect 72 106 73 107 
rect 72 107 73 108 
rect 72 108 73 109 
rect 72 109 73 110 
rect 72 110 73 111 
rect 72 111 73 112 
rect 72 112 73 113 
rect 72 113 73 114 
rect 72 114 73 115 
rect 72 115 73 116 
rect 72 116 73 117 
rect 72 117 73 118 
rect 72 118 73 119 
rect 72 119 73 120 
rect 72 120 73 121 
rect 72 121 73 122 
rect 72 122 73 123 
rect 72 123 73 124 
rect 72 124 73 125 
rect 72 125 73 126 
rect 72 126 73 127 
rect 72 127 73 128 
rect 72 128 73 129 
rect 72 129 73 130 
rect 72 130 73 131 
rect 72 131 73 132 
rect 72 132 73 133 
rect 72 133 73 134 
rect 72 134 73 135 
rect 72 135 73 136 
rect 72 136 73 137 
rect 72 137 73 138 
rect 72 138 73 139 
rect 72 139 73 140 
rect 72 140 73 141 
rect 72 141 73 142 
rect 72 142 73 143 
rect 72 143 73 144 
rect 72 144 73 145 
rect 72 145 73 146 
rect 72 146 73 147 
rect 72 147 73 148 
rect 72 148 73 149 
rect 72 149 73 150 
rect 72 150 73 151 
rect 72 151 73 152 
rect 72 152 73 153 
rect 72 153 73 154 
rect 72 154 73 155 
rect 72 155 73 156 
rect 72 156 73 157 
rect 72 157 73 158 
rect 72 158 73 159 
rect 72 159 73 160 
rect 72 160 73 161 
rect 72 162 73 163 
rect 72 163 73 164 
rect 72 164 73 165 
rect 72 165 73 166 
rect 72 166 73 167 
rect 72 167 73 168 
rect 72 168 73 169 
rect 72 169 73 170 
rect 72 170 73 171 
rect 72 171 73 172 
rect 72 172 73 173 
rect 72 173 73 174 
rect 72 174 73 175 
rect 72 175 73 176 
rect 72 176 73 177 
rect 72 177 73 178 
rect 72 178 73 179 
rect 72 179 73 180 
rect 72 180 73 181 
rect 72 181 73 182 
rect 72 182 73 183 
rect 72 183 73 184 
rect 72 184 73 185 
rect 72 185 73 186 
rect 72 186 73 187 
rect 72 187 73 188 
rect 72 188 73 189 
rect 72 189 73 190 
rect 72 190 73 191 
rect 72 191 73 192 
rect 72 192 73 193 
rect 72 193 73 194 
rect 72 194 73 195 
rect 72 195 73 196 
rect 72 196 73 197 
rect 72 197 73 198 
rect 72 198 73 199 
rect 72 199 73 200 
rect 72 200 73 201 
rect 72 201 73 202 
rect 72 202 73 203 
rect 72 203 73 204 
rect 72 204 73 205 
rect 72 205 73 206 
rect 72 206 73 207 
rect 72 207 73 208 
rect 72 208 73 209 
rect 72 209 73 210 
rect 72 210 73 211 
rect 72 211 73 212 
rect 72 212 73 213 
rect 72 213 73 214 
rect 72 214 73 215 
rect 72 215 73 216 
rect 72 216 73 217 
rect 72 217 73 218 
rect 72 218 73 219 
rect 72 219 73 220 
rect 72 220 73 221 
rect 72 221 73 222 
rect 72 222 73 223 
rect 72 223 73 224 
rect 72 224 73 225 
rect 72 225 73 226 
rect 72 226 73 227 
rect 72 227 73 228 
rect 72 228 73 229 
rect 72 229 73 230 
rect 72 230 73 231 
rect 72 231 73 232 
rect 72 232 73 233 
rect 72 233 73 234 
rect 72 234 73 235 
rect 72 235 73 236 
rect 72 236 73 237 
rect 72 237 73 238 
rect 72 238 73 239 
rect 72 239 73 240 
rect 72 240 73 241 
rect 72 241 73 242 
rect 72 242 73 243 
rect 72 243 73 244 
rect 72 244 73 245 
rect 72 245 73 246 
rect 72 246 73 247 
rect 72 247 73 248 
rect 72 248 73 249 
rect 72 249 73 250 
rect 72 250 73 251 
rect 72 251 73 252 
rect 72 252 73 253 
rect 72 253 73 254 
rect 72 254 73 255 
rect 72 255 73 256 
rect 72 256 73 257 
rect 72 257 73 258 
rect 72 258 73 259 
rect 72 259 73 260 
rect 72 260 73 261 
rect 72 261 73 262 
rect 72 262 73 263 
rect 72 263 73 264 
rect 72 264 73 265 
rect 72 265 73 266 
rect 72 266 73 267 
rect 72 267 73 268 
rect 72 268 73 269 
rect 72 269 73 270 
rect 72 270 73 271 
rect 72 271 73 272 
rect 72 272 73 273 
rect 72 273 73 274 
rect 72 274 73 275 
rect 72 275 73 276 
rect 72 276 73 277 
rect 72 277 73 278 
rect 72 278 73 279 
rect 72 279 73 280 
rect 72 280 73 281 
rect 72 281 73 282 
rect 72 282 73 283 
rect 72 283 73 284 
rect 72 289 73 290 
rect 72 292 73 293 
rect 72 305 73 306 
rect 72 307 73 308 
rect 72 310 73 311 
rect 73 1 74 2 
rect 73 3 74 4 
rect 73 8 74 9 
rect 73 9 74 10 
rect 73 14 74 15 
rect 73 16 74 17 
rect 73 17 74 18 
rect 73 40 74 41 
rect 73 41 74 42 
rect 73 59 74 60 
rect 73 160 74 161 
rect 73 161 74 162 
rect 73 283 74 284 
rect 73 289 74 290 
rect 73 292 74 293 
rect 73 305 74 306 
rect 73 307 74 308 
rect 73 310 74 311 
rect 74 1 75 2 
rect 74 3 75 4 
rect 74 8 75 9 
rect 74 14 75 15 
rect 74 17 75 18 
rect 74 18 75 19 
rect 74 19 75 20 
rect 74 20 75 21 
rect 74 21 75 22 
rect 74 22 75 23 
rect 74 23 75 24 
rect 74 36 75 37 
rect 74 37 75 38 
rect 74 38 75 39 
rect 74 39 75 40 
rect 74 40 75 41 
rect 74 55 75 56 
rect 74 59 75 60 
rect 74 66 75 67 
rect 74 97 75 98 
rect 74 98 75 99 
rect 74 99 75 100 
rect 74 100 75 101 
rect 74 101 75 102 
rect 74 102 75 103 
rect 74 129 75 130 
rect 74 134 75 135 
rect 74 148 75 149 
rect 74 161 75 162 
rect 74 164 75 165 
rect 74 242 75 243 
rect 74 244 75 245 
rect 74 257 75 258 
rect 74 283 75 284 
rect 74 289 75 290 
rect 74 292 75 293 
rect 74 305 75 306 
rect 74 307 75 308 
rect 74 310 75 311 
rect 75 1 76 2 
rect 75 3 76 4 
rect 75 8 76 9 
rect 75 23 76 24 
rect 75 36 76 37 
rect 75 55 76 56 
rect 75 66 76 67 
rect 75 68 76 69 
rect 75 69 76 70 
rect 75 70 76 71 
rect 75 72 76 73 
rect 75 97 76 98 
rect 75 129 76 130 
rect 75 131 76 132 
rect 75 134 76 135 
rect 75 136 76 137 
rect 75 148 76 149 
rect 75 152 76 153 
rect 75 161 76 162 
rect 75 164 76 165 
rect 75 210 76 211 
rect 75 211 76 212 
rect 75 212 76 213 
rect 75 213 76 214 
rect 75 214 76 215 
rect 75 215 76 216 
rect 75 232 76 233 
rect 75 242 76 243 
rect 75 244 76 245 
rect 75 257 76 258 
rect 75 289 76 290 
rect 75 292 76 293 
rect 75 305 76 306 
rect 75 307 76 308 
rect 75 310 76 311 
rect 76 1 77 2 
rect 76 3 77 4 
rect 76 8 77 9 
rect 76 23 77 24 
rect 76 36 77 37 
rect 76 55 77 56 
rect 76 66 77 67 
rect 76 68 77 69 
rect 76 72 77 73 
rect 76 97 77 98 
rect 76 99 77 100 
rect 76 129 77 130 
rect 76 131 77 132 
rect 76 134 77 135 
rect 76 136 77 137 
rect 76 148 77 149 
rect 76 152 77 153 
rect 76 161 77 162 
rect 76 164 77 165 
rect 76 215 77 216 
rect 76 225 77 226 
rect 76 232 77 233 
rect 76 242 77 243 
rect 76 244 77 245 
rect 76 257 77 258 
rect 76 289 77 290 
rect 76 292 77 293 
rect 76 305 77 306 
rect 76 307 77 308 
rect 76 310 77 311 
rect 77 1 78 2 
rect 77 3 78 4 
rect 77 8 78 9 
rect 77 23 78 24 
rect 77 36 78 37 
rect 77 55 78 56 
rect 77 66 78 67 
rect 77 68 78 69 
rect 77 72 78 73 
rect 77 97 78 98 
rect 77 99 78 100 
rect 77 129 78 130 
rect 77 131 78 132 
rect 77 134 78 135 
rect 77 136 78 137 
rect 77 148 78 149 
rect 77 152 78 153 
rect 77 161 78 162 
rect 77 164 78 165 
rect 77 215 78 216 
rect 77 225 78 226 
rect 77 232 78 233 
rect 77 242 78 243 
rect 77 244 78 245 
rect 77 257 78 258 
rect 77 289 78 290 
rect 77 292 78 293 
rect 77 305 78 306 
rect 77 307 78 308 
rect 77 310 78 311 
rect 78 1 79 2 
rect 78 3 79 4 
rect 78 8 79 9 
rect 78 23 79 24 
rect 78 36 79 37 
rect 78 55 79 56 
rect 78 66 79 67 
rect 78 68 79 69 
rect 78 72 79 73 
rect 78 97 79 98 
rect 78 99 79 100 
rect 78 129 79 130 
rect 78 131 79 132 
rect 78 134 79 135 
rect 78 136 79 137 
rect 78 148 79 149 
rect 78 152 79 153 
rect 78 161 79 162 
rect 78 164 79 165 
rect 78 215 79 216 
rect 78 225 79 226 
rect 78 226 79 227 
rect 78 227 79 228 
rect 78 228 79 229 
rect 78 232 79 233 
rect 78 242 79 243 
rect 78 244 79 245 
rect 78 257 79 258 
rect 78 289 79 290 
rect 78 292 79 293 
rect 78 305 79 306 
rect 78 307 79 308 
rect 78 310 79 311 
rect 79 1 80 2 
rect 79 3 80 4 
rect 79 8 80 9 
rect 79 23 80 24 
rect 79 36 80 37 
rect 79 46 80 47 
rect 79 55 80 56 
rect 79 66 80 67 
rect 79 68 80 69 
rect 79 72 80 73 
rect 79 97 80 98 
rect 79 99 80 100 
rect 79 129 80 130 
rect 79 131 80 132 
rect 79 134 80 135 
rect 79 136 80 137 
rect 79 139 80 140 
rect 79 148 80 149 
rect 79 152 80 153 
rect 79 155 80 156 
rect 79 161 80 162 
rect 79 164 80 165 
rect 79 215 80 216 
rect 79 216 80 217 
rect 79 228 80 229 
rect 79 229 80 230 
rect 79 230 80 231 
rect 79 232 80 233 
rect 79 238 80 239 
rect 79 242 80 243 
rect 79 244 80 245 
rect 79 257 80 258 
rect 79 283 80 284 
rect 79 286 80 287 
rect 79 289 80 290 
rect 79 292 80 293 
rect 79 302 80 303 
rect 79 305 80 306 
rect 79 307 80 308 
rect 79 310 80 311 
rect 80 1 81 2 
rect 80 3 81 4 
rect 80 8 81 9 
rect 80 23 81 24 
rect 80 32 81 33 
rect 80 33 81 34 
rect 80 34 81 35 
rect 80 35 81 36 
rect 80 36 81 37 
rect 80 38 81 39 
rect 80 46 81 47 
rect 80 55 81 56 
rect 80 66 81 67 
rect 80 68 81 69 
rect 80 72 81 73 
rect 80 73 81 74 
rect 80 96 81 97 
rect 80 97 81 98 
rect 80 99 81 100 
rect 80 112 81 113 
rect 80 113 81 114 
rect 80 114 81 115 
rect 80 115 81 116 
rect 80 116 81 117 
rect 80 117 81 118 
rect 80 118 81 119 
rect 80 119 81 120 
rect 80 129 81 130 
rect 80 131 81 132 
rect 80 134 81 135 
rect 80 136 81 137 
rect 80 139 81 140 
rect 80 148 81 149 
rect 80 152 81 153 
rect 80 153 81 154 
rect 80 155 81 156 
rect 80 161 81 162 
rect 80 164 81 165 
rect 80 216 81 217 
rect 80 217 81 218 
rect 80 230 81 231 
rect 80 232 81 233 
rect 80 233 81 234 
rect 80 238 81 239 
rect 80 242 81 243 
rect 80 244 81 245 
rect 80 256 81 257 
rect 80 257 81 258 
rect 80 283 81 284 
rect 80 286 81 287 
rect 80 289 81 290 
rect 80 292 81 293 
rect 80 302 81 303 
rect 80 305 81 306 
rect 80 307 81 308 
rect 80 310 81 311 
rect 80 311 81 312 
rect 81 1 82 2 
rect 81 3 82 4 
rect 81 8 82 9 
rect 81 23 82 24 
rect 81 25 82 26 
rect 81 26 82 27 
rect 81 27 82 28 
rect 81 28 82 29 
rect 81 29 82 30 
rect 81 30 82 31 
rect 81 31 82 32 
rect 81 32 82 33 
rect 81 38 82 39 
rect 81 46 82 47 
rect 81 55 82 56 
rect 81 66 82 67 
rect 81 68 82 69 
rect 81 73 82 74 
rect 81 89 82 90 
rect 81 90 82 91 
rect 81 91 82 92 
rect 81 92 82 93 
rect 81 93 82 94 
rect 81 94 82 95 
rect 81 95 82 96 
rect 81 96 82 97 
rect 81 99 82 100 
rect 81 112 82 113 
rect 81 119 82 120 
rect 81 120 82 121 
rect 81 121 82 122 
rect 81 122 82 123 
rect 81 123 82 124 
rect 81 124 82 125 
rect 81 125 82 126 
rect 81 126 82 127 
rect 81 129 82 130 
rect 81 131 82 132 
rect 81 134 82 135 
rect 81 136 82 137 
rect 81 138 82 139 
rect 81 139 82 140 
rect 81 145 82 146 
rect 81 146 82 147 
rect 81 147 82 148 
rect 81 148 82 149 
rect 81 153 82 154 
rect 81 154 82 155 
rect 81 155 82 156 
rect 81 161 82 162 
rect 81 164 82 165 
rect 81 165 82 166 
rect 81 166 82 167 
rect 81 167 82 168 
rect 81 168 82 169 
rect 81 169 82 170 
rect 81 170 82 171 
rect 81 171 82 172 
rect 81 172 82 173 
rect 81 173 82 174 
rect 81 174 82 175 
rect 81 175 82 176 
rect 81 176 82 177 
rect 81 177 82 178 
rect 81 178 82 179 
rect 81 179 82 180 
rect 81 180 82 181 
rect 81 181 82 182 
rect 81 182 82 183 
rect 81 183 82 184 
rect 81 184 82 185 
rect 81 185 82 186 
rect 81 186 82 187 
rect 81 187 82 188 
rect 81 188 82 189 
rect 81 189 82 190 
rect 81 190 82 191 
rect 81 191 82 192 
rect 81 192 82 193 
rect 81 193 82 194 
rect 81 194 82 195 
rect 81 195 82 196 
rect 81 196 82 197 
rect 81 197 82 198 
rect 81 198 82 199 
rect 81 199 82 200 
rect 81 200 82 201 
rect 81 201 82 202 
rect 81 202 82 203 
rect 81 203 82 204 
rect 81 204 82 205 
rect 81 205 82 206 
rect 81 206 82 207 
rect 81 207 82 208 
rect 81 208 82 209 
rect 81 209 82 210 
rect 81 210 82 211 
rect 81 211 82 212 
rect 81 212 82 213 
rect 81 213 82 214 
rect 81 214 82 215 
rect 81 215 82 216 
rect 81 217 82 218 
rect 81 230 82 231 
rect 81 233 82 234 
rect 81 234 82 235 
rect 81 235 82 236 
rect 81 237 82 238 
rect 81 238 82 239 
rect 81 242 82 243 
rect 81 244 82 245 
rect 81 254 82 255 
rect 81 255 82 256 
rect 81 256 82 257 
rect 81 280 82 281 
rect 81 281 82 282 
rect 81 282 82 283 
rect 81 283 82 284 
rect 81 285 82 286 
rect 81 286 82 287 
rect 81 289 82 290 
rect 81 292 82 293 
rect 81 302 82 303 
rect 81 305 82 306 
rect 81 307 82 308 
rect 81 311 82 312 
rect 82 1 83 2 
rect 82 3 83 4 
rect 82 8 83 9 
rect 82 21 83 22 
rect 82 23 83 24 
rect 82 38 83 39 
rect 82 46 83 47 
rect 82 55 83 56 
rect 82 66 83 67 
rect 82 68 83 69 
rect 82 69 83 70 
rect 82 73 83 74 
rect 82 75 83 76 
rect 82 76 83 77 
rect 82 77 83 78 
rect 82 78 83 79 
rect 82 79 83 80 
rect 82 80 83 81 
rect 82 81 83 82 
rect 82 82 83 83 
rect 82 83 83 84 
rect 82 84 83 85 
rect 82 85 83 86 
rect 82 86 83 87 
rect 82 87 83 88 
rect 82 88 83 89 
rect 82 89 83 90 
rect 82 99 83 100 
rect 82 112 83 113 
rect 82 129 83 130 
rect 82 131 83 132 
rect 82 134 83 135 
rect 82 136 83 137 
rect 82 138 83 139 
rect 82 145 83 146 
rect 82 161 83 162 
rect 82 215 83 216 
rect 82 217 83 218 
rect 82 229 83 230 
rect 82 235 83 236 
rect 82 242 83 243 
rect 82 244 83 245 
rect 82 254 83 255 
rect 82 280 83 281 
rect 82 284 83 285 
rect 82 285 83 286 
rect 82 289 83 290 
rect 82 292 83 293 
rect 82 305 83 306 
rect 82 307 83 308 
rect 82 309 83 310 
rect 82 311 83 312 
rect 83 1 84 2 
rect 83 3 84 4 
rect 83 8 84 9 
rect 83 21 84 22 
rect 83 23 84 24 
rect 83 38 84 39 
rect 83 46 84 47 
rect 83 55 84 56 
rect 83 66 84 67 
rect 83 69 84 70 
rect 83 71 84 72 
rect 83 73 84 74 
rect 83 99 84 100 
rect 83 100 84 101 
rect 83 101 84 102 
rect 83 102 84 103 
rect 83 112 84 113 
rect 83 129 84 130 
rect 83 131 84 132 
rect 83 134 84 135 
rect 83 136 84 137 
rect 83 145 84 146 
rect 83 161 84 162 
rect 83 164 84 165 
rect 83 165 84 166 
rect 83 166 84 167 
rect 83 199 84 200 
rect 83 215 84 216 
rect 83 217 84 218 
rect 83 229 84 230 
rect 83 235 84 236 
rect 83 242 84 243 
rect 83 244 84 245 
rect 83 254 84 255 
rect 83 280 84 281 
rect 83 282 84 283 
rect 83 283 84 284 
rect 83 284 84 285 
rect 83 289 84 290 
rect 83 292 84 293 
rect 83 305 84 306 
rect 83 307 84 308 
rect 83 309 84 310 
rect 83 311 84 312 
rect 84 1 85 2 
rect 84 3 85 4 
rect 84 8 85 9 
rect 84 21 85 22 
rect 84 23 85 24 
rect 84 38 85 39 
rect 84 44 85 45 
rect 84 45 85 46 
rect 84 46 85 47 
rect 84 55 85 56 
rect 84 66 85 67 
rect 84 69 85 70 
rect 84 71 85 72 
rect 84 73 85 74 
rect 84 88 85 89 
rect 84 102 85 103 
rect 84 112 85 113 
rect 84 129 85 130 
rect 84 131 85 132 
rect 84 136 85 137 
rect 84 145 85 146 
rect 84 161 85 162 
rect 84 164 85 165 
rect 84 199 85 200 
rect 84 215 85 216 
rect 84 217 85 218 
rect 84 229 85 230 
rect 84 235 85 236 
rect 84 242 85 243 
rect 84 244 85 245 
rect 84 254 85 255 
rect 84 278 85 279 
rect 84 280 85 281 
rect 84 289 85 290 
rect 84 292 85 293 
rect 84 305 85 306 
rect 84 307 85 308 
rect 84 309 85 310 
rect 84 311 85 312 
rect 85 1 86 2 
rect 85 3 86 4 
rect 85 8 86 9 
rect 85 21 86 22 
rect 85 23 86 24 
rect 85 38 86 39 
rect 85 42 86 43 
rect 85 43 86 44 
rect 85 44 86 45 
rect 85 55 86 56 
rect 85 66 86 67 
rect 85 69 86 70 
rect 85 71 86 72 
rect 85 73 86 74 
rect 85 88 86 89 
rect 85 102 86 103 
rect 85 110 86 111 
rect 85 111 86 112 
rect 85 112 86 113 
rect 85 129 86 130 
rect 85 131 86 132 
rect 85 136 86 137 
rect 85 145 86 146 
rect 85 161 86 162 
rect 85 164 86 165 
rect 85 199 86 200 
rect 85 215 86 216 
rect 85 217 86 218 
rect 85 229 86 230 
rect 85 235 86 236 
rect 85 242 86 243 
rect 85 244 86 245 
rect 85 254 86 255 
rect 85 278 86 279 
rect 85 280 86 281 
rect 85 289 86 290 
rect 85 292 86 293 
rect 85 305 86 306 
rect 85 307 86 308 
rect 85 309 86 310 
rect 85 311 86 312 
rect 86 1 87 2 
rect 86 3 87 4 
rect 86 8 87 9 
rect 86 21 87 22 
rect 86 23 87 24 
rect 86 38 87 39 
rect 86 40 87 41 
rect 86 41 87 42 
rect 86 42 87 43 
rect 86 45 87 46 
rect 86 46 87 47 
rect 86 47 87 48 
rect 86 48 87 49 
rect 86 49 87 50 
rect 86 51 87 52 
rect 86 52 87 53 
rect 86 53 87 54 
rect 86 54 87 55 
rect 86 55 87 56 
rect 86 66 87 67 
rect 86 69 87 70 
rect 86 71 87 72 
rect 86 73 87 74 
rect 86 88 87 89 
rect 86 99 87 100 
rect 86 100 87 101 
rect 86 102 87 103 
rect 86 129 87 130 
rect 86 131 87 132 
rect 86 136 87 137 
rect 86 152 87 153 
rect 86 153 87 154 
rect 86 154 87 155 
rect 86 155 87 156 
rect 86 156 87 157 
rect 86 161 87 162 
rect 86 164 87 165 
rect 86 199 87 200 
rect 86 215 87 216 
rect 86 217 87 218 
rect 86 229 87 230 
rect 86 235 87 236 
rect 86 242 87 243 
rect 86 244 87 245 
rect 86 254 87 255 
rect 86 278 87 279 
rect 86 280 87 281 
rect 86 289 87 290 
rect 86 292 87 293 
rect 86 305 87 306 
rect 86 307 87 308 
rect 86 309 87 310 
rect 86 311 87 312 
rect 87 1 88 2 
rect 87 3 88 4 
rect 87 8 88 9 
rect 87 21 88 22 
rect 87 23 88 24 
rect 87 38 88 39 
rect 87 40 88 41 
rect 87 43 88 44 
rect 87 44 88 45 
rect 87 45 88 46 
rect 87 49 88 50 
rect 87 50 88 51 
rect 87 66 88 67 
rect 87 71 88 72 
rect 87 73 88 74 
rect 87 87 88 88 
rect 87 88 88 89 
rect 87 99 88 100 
rect 87 102 88 103 
rect 87 129 88 130 
rect 87 131 88 132 
rect 87 136 88 137 
rect 87 147 88 148 
rect 87 148 88 149 
rect 87 149 88 150 
rect 87 150 88 151 
rect 87 151 88 152 
rect 87 152 88 153 
rect 87 156 88 157 
rect 87 157 88 158 
rect 87 161 88 162 
rect 87 164 88 165 
rect 87 199 88 200 
rect 87 215 88 216 
rect 87 217 88 218 
rect 87 229 88 230 
rect 87 235 88 236 
rect 87 242 88 243 
rect 87 244 88 245 
rect 87 254 88 255 
rect 87 278 88 279 
rect 87 280 88 281 
rect 87 289 88 290 
rect 87 292 88 293 
rect 87 305 88 306 
rect 87 307 88 308 
rect 87 309 88 310 
rect 87 311 88 312 
rect 88 1 89 2 
rect 88 3 89 4 
rect 88 8 89 9 
rect 88 21 89 22 
rect 88 23 89 24 
rect 88 37 89 38 
rect 88 38 89 39 
rect 88 41 89 42 
rect 88 42 89 43 
rect 88 43 89 44 
rect 88 46 89 47 
rect 88 47 89 48 
rect 88 48 89 49 
rect 88 50 89 51 
rect 88 51 89 52 
rect 88 52 89 53 
rect 88 53 89 54 
rect 88 54 89 55 
rect 88 55 89 56 
rect 88 56 89 57 
rect 88 57 89 58 
rect 88 58 89 59 
rect 88 59 89 60 
rect 88 60 89 61 
rect 88 61 89 62 
rect 88 62 89 63 
rect 88 66 89 67 
rect 88 69 89 70 
rect 88 70 89 71 
rect 88 71 89 72 
rect 88 73 89 74 
rect 88 86 89 87 
rect 88 87 89 88 
rect 88 89 89 90 
rect 88 90 89 91 
rect 88 91 89 92 
rect 88 92 89 93 
rect 88 93 89 94 
rect 88 94 89 95 
rect 88 95 89 96 
rect 88 96 89 97 
rect 88 97 89 98 
rect 88 98 89 99 
rect 88 99 89 100 
rect 88 102 89 103 
rect 88 105 89 106 
rect 88 106 89 107 
rect 88 107 89 108 
rect 88 108 89 109 
rect 88 109 89 110 
rect 88 110 89 111 
rect 88 111 89 112 
rect 88 112 89 113 
rect 88 113 89 114 
rect 88 114 89 115 
rect 88 115 89 116 
rect 88 116 89 117 
rect 88 117 89 118 
rect 88 118 89 119 
rect 88 119 89 120 
rect 88 120 89 121 
rect 88 121 89 122 
rect 88 122 89 123 
rect 88 123 89 124 
rect 88 124 89 125 
rect 88 125 89 126 
rect 88 126 89 127 
rect 88 127 89 128 
rect 88 128 89 129 
rect 88 129 89 130 
rect 88 131 89 132 
rect 88 133 89 134 
rect 88 136 89 137 
rect 88 138 89 139 
rect 88 139 89 140 
rect 88 140 89 141 
rect 88 141 89 142 
rect 88 142 89 143 
rect 88 143 89 144 
rect 88 144 89 145 
rect 88 145 89 146 
rect 88 146 89 147 
rect 88 147 89 148 
rect 88 153 89 154 
rect 88 154 89 155 
rect 88 155 89 156 
rect 88 157 89 158 
rect 88 158 89 159 
rect 88 161 89 162 
rect 88 164 89 165 
rect 88 174 89 175 
rect 88 175 89 176 
rect 88 176 89 177 
rect 88 185 89 186 
rect 88 186 89 187 
rect 88 187 89 188 
rect 88 199 89 200 
rect 88 215 89 216 
rect 88 217 89 218 
rect 88 218 89 219 
rect 88 219 89 220 
rect 88 220 89 221 
rect 88 221 89 222 
rect 88 222 89 223 
rect 88 223 89 224 
rect 88 224 89 225 
rect 88 229 89 230 
rect 88 235 89 236 
rect 88 236 89 237 
rect 88 237 89 238 
rect 88 238 89 239 
rect 88 242 89 243 
rect 88 244 89 245 
rect 88 249 89 250 
rect 88 250 89 251 
rect 88 251 89 252 
rect 88 252 89 253 
rect 88 253 89 254 
rect 88 254 89 255 
rect 88 263 89 264 
rect 88 264 89 265 
rect 88 265 89 266 
rect 88 266 89 267 
rect 88 267 89 268 
rect 88 277 89 278 
rect 88 278 89 279 
rect 88 280 89 281 
rect 88 289 89 290 
rect 88 292 89 293 
rect 88 305 89 306 
rect 88 307 89 308 
rect 88 309 89 310 
rect 88 311 89 312 
rect 89 1 90 2 
rect 89 3 90 4 
rect 89 8 90 9 
rect 89 21 90 22 
rect 89 23 90 24 
rect 89 36 90 37 
rect 89 37 90 38 
rect 89 40 90 41 
rect 89 41 90 42 
rect 89 46 90 47 
rect 89 48 90 49 
rect 89 49 90 50 
rect 89 62 90 63 
rect 89 66 90 67 
rect 89 69 90 70 
rect 89 72 90 73 
rect 89 73 90 74 
rect 89 86 90 87 
rect 89 88 90 89 
rect 89 89 90 90 
rect 89 104 90 105 
rect 89 105 90 106 
rect 89 132 90 133 
rect 89 133 90 134 
rect 89 136 90 137 
rect 89 152 90 153 
rect 89 153 90 154 
rect 89 155 90 156 
rect 89 158 90 159 
rect 89 161 90 162 
rect 89 164 90 165 
rect 89 174 90 175 
rect 89 176 90 177 
rect 89 177 90 178 
rect 89 184 90 185 
rect 89 185 90 186 
rect 89 187 90 188 
rect 89 199 90 200 
rect 89 215 90 216 
rect 89 224 90 225 
rect 89 229 90 230 
rect 89 238 90 239 
rect 89 242 90 243 
rect 89 244 90 245 
rect 89 248 90 249 
rect 89 249 90 250 
rect 89 263 90 264 
rect 89 267 90 268 
rect 89 277 90 278 
rect 89 280 90 281 
rect 89 289 90 290 
rect 89 292 90 293 
rect 89 305 90 306 
rect 89 307 90 308 
rect 89 309 90 310 
rect 89 311 90 312 
rect 89 312 90 313 
rect 90 1 91 2 
rect 90 3 91 4 
rect 90 8 91 9 
rect 90 21 91 22 
rect 90 23 91 24 
rect 90 36 91 37 
rect 90 38 91 39 
rect 90 39 91 40 
rect 90 40 91 41 
rect 90 46 91 47 
rect 90 49 91 50 
rect 90 50 91 51 
rect 90 51 91 52 
rect 90 62 91 63 
rect 90 66 91 67 
rect 90 69 91 70 
rect 90 72 91 73 
rect 90 86 91 87 
rect 90 88 91 89 
rect 90 102 91 103 
rect 90 103 91 104 
rect 90 104 91 105 
rect 90 131 91 132 
rect 90 132 91 133 
rect 90 134 91 135 
rect 90 135 91 136 
rect 90 136 91 137 
rect 90 145 91 146 
rect 90 146 91 147 
rect 90 147 91 148 
rect 90 148 91 149 
rect 90 149 91 150 
rect 90 150 91 151 
rect 90 151 91 152 
rect 90 152 91 153 
rect 90 155 91 156 
rect 90 158 91 159 
rect 90 161 91 162 
rect 90 164 91 165 
rect 90 174 91 175 
rect 90 177 91 178 
rect 90 184 91 185 
rect 90 187 91 188 
rect 90 195 91 196 
rect 90 199 91 200 
rect 90 215 91 216 
rect 90 225 91 226 
rect 90 226 91 227 
rect 90 227 91 228 
rect 90 228 91 229 
rect 90 229 91 230 
rect 90 238 91 239 
rect 90 242 91 243 
rect 90 244 91 245 
rect 90 247 91 248 
rect 90 248 91 249 
rect 90 263 91 264 
rect 90 267 91 268 
rect 90 277 91 278 
rect 90 280 91 281 
rect 90 289 91 290 
rect 90 292 91 293 
rect 90 305 91 306 
rect 90 307 91 308 
rect 90 309 91 310 
rect 90 310 91 311 
rect 90 312 91 313 
rect 91 1 92 2 
rect 91 3 92 4 
rect 91 8 92 9 
rect 91 21 92 22 
rect 91 23 92 24 
rect 91 36 92 37 
rect 91 38 92 39 
rect 91 51 92 52 
rect 91 66 92 67 
rect 91 69 92 70 
rect 91 72 92 73 
rect 91 86 92 87 
rect 91 88 92 89 
rect 91 102 92 103 
rect 91 131 92 132 
rect 91 134 92 135 
rect 91 145 92 146 
rect 91 161 92 162 
rect 91 164 92 165 
rect 91 177 92 178 
rect 91 184 92 185 
rect 91 195 92 196 
rect 91 199 92 200 
rect 91 215 92 216 
rect 91 225 92 226 
rect 91 242 92 243 
rect 91 244 92 245 
rect 91 247 92 248 
rect 91 263 92 264 
rect 91 277 92 278 
rect 91 280 92 281 
rect 91 289 92 290 
rect 91 292 92 293 
rect 91 305 92 306 
rect 91 307 92 308 
rect 91 310 92 311 
rect 91 312 92 313 
rect 92 1 93 2 
rect 92 3 93 4 
rect 92 8 93 9 
rect 92 21 93 22 
rect 92 23 93 24 
rect 92 36 93 37 
rect 92 38 93 39 
rect 92 51 93 52 
rect 92 65 93 66 
rect 92 66 93 67 
rect 92 69 93 70 
rect 92 72 93 73 
rect 92 86 93 87 
rect 92 88 93 89 
rect 92 102 93 103 
rect 92 131 93 132 
rect 92 134 93 135 
rect 92 145 93 146 
rect 92 161 93 162 
rect 92 164 93 165 
rect 92 177 93 178 
rect 92 184 93 185 
rect 92 195 93 196 
rect 92 199 93 200 
rect 92 215 93 216 
rect 92 225 93 226 
rect 92 242 93 243 
rect 92 244 93 245 
rect 92 247 93 248 
rect 92 263 93 264 
rect 92 277 93 278 
rect 92 280 93 281 
rect 92 289 93 290 
rect 92 292 93 293 
rect 92 305 93 306 
rect 92 307 93 308 
rect 92 310 93 311 
rect 92 312 93 313 
rect 93 1 94 2 
rect 93 3 94 4 
rect 93 8 94 9 
rect 93 21 94 22 
rect 93 23 94 24 
rect 93 36 94 37 
rect 93 38 94 39 
rect 93 51 94 52 
rect 93 69 94 70 
rect 93 72 94 73 
rect 93 86 94 87 
rect 93 88 94 89 
rect 93 102 94 103 
rect 93 131 94 132 
rect 93 134 94 135 
rect 93 145 94 146 
rect 93 161 94 162 
rect 93 164 94 165 
rect 93 177 94 178 
rect 93 184 94 185 
rect 93 195 94 196 
rect 93 199 94 200 
rect 93 215 94 216 
rect 93 225 94 226 
rect 93 242 94 243 
rect 93 244 94 245 
rect 93 247 94 248 
rect 93 263 94 264 
rect 93 277 94 278 
rect 93 280 94 281 
rect 93 289 94 290 
rect 93 292 94 293 
rect 93 305 94 306 
rect 93 307 94 308 
rect 93 310 94 311 
rect 93 312 94 313 
rect 94 1 95 2 
rect 94 3 95 4 
rect 94 8 95 9 
rect 94 18 95 19 
rect 94 19 95 20 
rect 94 20 95 21 
rect 94 21 95 22 
rect 94 23 95 24 
rect 94 36 95 37 
rect 94 38 95 39 
rect 94 51 95 52 
rect 94 52 95 53 
rect 94 65 95 66 
rect 94 66 95 67 
rect 94 67 95 68 
rect 94 68 95 69 
rect 94 69 95 70 
rect 94 72 95 73 
rect 94 86 95 87 
rect 94 88 95 89 
rect 94 102 95 103 
rect 94 129 95 130 
rect 94 130 95 131 
rect 94 131 95 132 
rect 94 134 95 135 
rect 94 145 95 146 
rect 94 161 95 162 
rect 94 164 95 165 
rect 94 177 95 178 
rect 94 184 95 185 
rect 94 195 95 196 
rect 94 199 95 200 
rect 94 215 95 216 
rect 94 216 95 217 
rect 94 225 95 226 
rect 94 242 95 243 
rect 94 244 95 245 
rect 94 247 95 248 
rect 94 263 95 264 
rect 94 273 95 274 
rect 94 274 95 275 
rect 94 275 95 276 
rect 94 276 95 277 
rect 94 277 95 278 
rect 94 280 95 281 
rect 94 289 95 290 
rect 94 292 95 293 
rect 94 305 95 306 
rect 94 307 95 308 
rect 94 310 95 311 
rect 94 312 95 313 
rect 95 1 96 2 
rect 95 3 96 4 
rect 95 8 96 9 
rect 95 18 96 19 
rect 95 23 96 24 
rect 95 27 96 28 
rect 95 36 96 37 
rect 95 38 96 39 
rect 95 46 96 47 
rect 95 52 96 53 
rect 95 65 96 66 
rect 95 72 96 73 
rect 95 85 96 86 
rect 95 86 96 87 
rect 95 88 96 89 
rect 95 101 96 102 
rect 95 102 96 103 
rect 95 129 96 130 
rect 95 134 96 135 
rect 95 139 96 140 
rect 95 145 96 146 
rect 95 155 96 156 
rect 95 158 96 159 
rect 95 161 96 162 
rect 95 164 96 165 
rect 95 165 96 166 
rect 95 177 96 178 
rect 95 184 96 185 
rect 95 187 96 188 
rect 95 195 96 196 
rect 95 199 96 200 
rect 95 206 96 207 
rect 95 216 96 217 
rect 95 222 96 223 
rect 95 225 96 226 
rect 95 238 96 239 
rect 95 242 96 243 
rect 95 244 96 245 
rect 95 245 96 246 
rect 95 247 96 248 
rect 95 251 96 252 
rect 95 263 96 264 
rect 95 273 96 274 
rect 95 280 96 281 
rect 95 289 96 290 
rect 95 292 96 293 
rect 95 305 96 306 
rect 95 307 96 308 
rect 95 310 96 311 
rect 95 312 96 313 
rect 96 1 97 2 
rect 96 3 97 4 
rect 96 8 97 9 
rect 96 18 97 19 
rect 96 23 97 24 
rect 96 27 97 28 
rect 96 36 97 37 
rect 96 38 97 39 
rect 96 46 97 47 
rect 96 52 97 53 
rect 96 65 97 66 
rect 96 72 97 73 
rect 96 128 97 129 
rect 96 129 97 130 
rect 96 134 97 135 
rect 96 139 97 140 
rect 96 145 97 146 
rect 96 155 97 156 
rect 96 158 97 159 
rect 96 161 97 162 
rect 96 165 97 166 
rect 96 177 97 178 
rect 96 184 97 185 
rect 96 187 97 188 
rect 96 195 97 196 
rect 96 199 97 200 
rect 96 206 97 207 
rect 96 216 97 217 
rect 96 222 97 223 
rect 96 224 97 225 
rect 96 225 97 226 
rect 96 238 97 239 
rect 96 242 97 243 
rect 96 245 97 246 
rect 96 247 97 248 
rect 96 251 97 252 
rect 96 272 97 273 
rect 96 273 97 274 
rect 96 280 97 281 
rect 96 289 97 290 
rect 96 292 97 293 
rect 96 305 97 306 
rect 96 307 97 308 
rect 96 310 97 311 
rect 96 312 97 313 
rect 97 1 98 2 
rect 97 3 98 4 
rect 97 8 98 9 
rect 97 18 98 19 
rect 97 20 98 21 
rect 97 23 98 24 
rect 97 27 98 28 
rect 97 28 98 29 
rect 97 29 98 30 
rect 97 30 98 31 
rect 97 31 98 32 
rect 97 32 98 33 
rect 97 33 98 34 
rect 97 34 98 35 
rect 97 35 98 36 
rect 97 36 98 37 
rect 97 38 98 39 
rect 97 46 98 47 
rect 97 47 98 48 
rect 97 48 98 49 
rect 97 49 98 50 
rect 97 50 98 51 
rect 97 52 98 53 
rect 97 56 98 57 
rect 97 57 98 58 
rect 97 58 98 59 
rect 97 59 98 60 
rect 97 60 98 61 
rect 97 61 98 62 
rect 97 62 98 63 
rect 97 63 98 64 
rect 97 64 98 65 
rect 97 65 98 66 
rect 97 68 98 69 
rect 97 69 98 70 
rect 97 72 98 73 
rect 97 81 98 82 
rect 97 82 98 83 
rect 97 83 98 84 
rect 97 84 98 85 
rect 97 85 98 86 
rect 97 86 98 87 
rect 97 87 98 88 
rect 97 88 98 89 
rect 97 89 98 90 
rect 97 90 98 91 
rect 97 91 98 92 
rect 97 92 98 93 
rect 97 93 98 94 
rect 97 94 98 95 
rect 97 95 98 96 
rect 97 96 98 97 
rect 97 97 98 98 
rect 97 98 98 99 
rect 97 99 98 100 
rect 97 100 98 101 
rect 97 101 98 102 
rect 97 102 98 103 
rect 97 103 98 104 
rect 97 104 98 105 
rect 97 105 98 106 
rect 97 106 98 107 
rect 97 107 98 108 
rect 97 108 98 109 
rect 97 109 98 110 
rect 97 110 98 111 
rect 97 111 98 112 
rect 97 112 98 113 
rect 97 113 98 114 
rect 97 114 98 115 
rect 97 115 98 116 
rect 97 116 98 117 
rect 97 117 98 118 
rect 97 118 98 119 
rect 97 119 98 120 
rect 97 120 98 121 
rect 97 121 98 122 
rect 97 122 98 123 
rect 97 123 98 124 
rect 97 124 98 125 
rect 97 125 98 126 
rect 97 126 98 127 
rect 97 127 98 128 
rect 97 128 98 129 
rect 97 134 98 135 
rect 97 139 98 140 
rect 97 140 98 141 
rect 97 141 98 142 
rect 97 142 98 143 
rect 97 143 98 144 
rect 97 145 98 146 
rect 97 147 98 148 
rect 97 148 98 149 
rect 97 149 98 150 
rect 97 150 98 151 
rect 97 151 98 152 
rect 97 152 98 153 
rect 97 153 98 154 
rect 97 154 98 155 
rect 97 155 98 156 
rect 97 158 98 159 
rect 97 159 98 160 
rect 97 161 98 162 
rect 97 165 98 166 
rect 97 166 98 167 
rect 97 177 98 178 
rect 97 184 98 185 
rect 97 187 98 188 
rect 97 195 98 196 
rect 97 199 98 200 
rect 97 206 98 207 
rect 97 216 98 217 
rect 97 219 98 220 
rect 97 220 98 221 
rect 97 221 98 222 
rect 97 222 98 223 
rect 97 224 98 225 
rect 97 235 98 236 
rect 97 236 98 237 
rect 97 237 98 238 
rect 97 238 98 239 
rect 97 242 98 243 
rect 97 247 98 248 
rect 97 249 98 250 
rect 97 251 98 252 
rect 97 252 98 253 
rect 97 253 98 254 
rect 97 254 98 255 
rect 97 255 98 256 
rect 97 256 98 257 
rect 97 257 98 258 
rect 97 258 98 259 
rect 97 259 98 260 
rect 97 260 98 261 
rect 97 261 98 262 
rect 97 262 98 263 
rect 97 263 98 264 
rect 97 264 98 265 
rect 97 265 98 266 
rect 97 266 98 267 
rect 97 267 98 268 
rect 97 268 98 269 
rect 97 269 98 270 
rect 97 270 98 271 
rect 97 271 98 272 
rect 97 272 98 273 
rect 97 280 98 281 
rect 97 289 98 290 
rect 97 292 98 293 
rect 97 305 98 306 
rect 97 307 98 308 
rect 97 310 98 311 
rect 97 312 98 313 
rect 98 1 99 2 
rect 98 3 99 4 
rect 98 8 99 9 
rect 98 18 99 19 
rect 98 20 99 21 
rect 98 23 99 24 
rect 98 38 99 39 
rect 98 50 99 51 
rect 98 52 99 53 
rect 98 56 99 57 
rect 98 68 99 69 
rect 98 72 99 73 
rect 98 81 99 82 
rect 98 134 99 135 
rect 98 145 99 146 
rect 98 147 99 148 
rect 98 161 99 162 
rect 98 166 99 167 
rect 98 177 99 178 
rect 98 184 99 185 
rect 98 187 99 188 
rect 98 190 99 191 
rect 98 191 99 192 
rect 98 192 99 193 
rect 98 193 99 194 
rect 98 194 99 195 
rect 98 195 99 196 
rect 98 199 99 200 
rect 98 202 99 203 
rect 98 203 99 204 
rect 98 204 99 205 
rect 98 205 99 206 
rect 98 206 99 207 
rect 98 216 99 217 
rect 98 224 99 225 
rect 98 235 99 236 
rect 98 242 99 243 
rect 98 247 99 248 
rect 98 249 99 250 
rect 98 280 99 281 
rect 98 289 99 290 
rect 98 292 99 293 
rect 98 303 99 304 
rect 98 305 99 306 
rect 98 308 99 309 
rect 98 309 99 310 
rect 98 310 99 311 
rect 98 312 99 313 
rect 99 1 100 2 
rect 99 3 100 4 
rect 99 8 100 9 
rect 99 18 100 19 
rect 99 20 100 21 
rect 99 23 100 24 
rect 99 38 100 39 
rect 99 50 100 51 
rect 99 52 100 53 
rect 99 56 100 57 
rect 99 68 100 69 
rect 99 72 100 73 
rect 99 81 100 82 
rect 99 87 100 88 
rect 99 94 100 95 
rect 99 95 100 96 
rect 99 96 100 97 
rect 99 97 100 98 
rect 99 101 100 102 
rect 99 119 100 120 
rect 99 134 100 135 
rect 99 135 100 136 
rect 99 145 100 146 
rect 99 147 100 148 
rect 99 161 100 162 
rect 99 166 100 167 
rect 99 177 100 178 
rect 99 184 100 185 
rect 99 187 100 188 
rect 99 199 100 200 
rect 99 216 100 217 
rect 99 224 100 225 
rect 99 235 100 236 
rect 99 242 100 243 
rect 99 247 100 248 
rect 99 249 100 250 
rect 99 250 100 251 
rect 99 251 100 252 
rect 99 252 100 253 
rect 99 253 100 254 
rect 99 254 100 255 
rect 99 255 100 256 
rect 99 256 100 257 
rect 99 257 100 258 
rect 99 258 100 259 
rect 99 259 100 260 
rect 99 260 100 261 
rect 99 261 100 262 
rect 99 262 100 263 
rect 99 263 100 264 
rect 99 264 100 265 
rect 99 265 100 266 
rect 99 266 100 267 
rect 99 267 100 268 
rect 99 268 100 269 
rect 99 269 100 270 
rect 99 270 100 271 
rect 99 271 100 272 
rect 99 272 100 273 
rect 99 273 100 274 
rect 99 274 100 275 
rect 99 275 100 276 
rect 99 276 100 277 
rect 99 280 100 281 
rect 99 289 100 290 
rect 99 292 100 293 
rect 99 303 100 304 
rect 99 305 100 306 
rect 99 308 100 309 
rect 99 311 100 312 
rect 99 312 100 313 
rect 100 1 101 2 
rect 100 3 101 4 
rect 100 8 101 9 
rect 100 18 101 19 
rect 100 20 101 21 
rect 100 23 101 24 
rect 100 38 101 39 
rect 100 50 101 51 
rect 100 52 101 53 
rect 100 56 101 57 
rect 100 68 101 69 
rect 100 72 101 73 
rect 100 81 101 82 
rect 100 84 101 85 
rect 100 87 101 88 
rect 100 94 101 95 
rect 100 101 101 102 
rect 100 115 101 116 
rect 100 116 101 117 
rect 100 117 101 118 
rect 100 118 101 119 
rect 100 119 101 120 
rect 100 135 101 136 
rect 100 145 101 146 
rect 100 147 101 148 
rect 100 161 101 162 
rect 100 166 101 167 
rect 100 177 101 178 
rect 100 184 101 185 
rect 100 187 101 188 
rect 100 188 101 189 
rect 100 189 101 190 
rect 100 190 101 191 
rect 100 191 101 192 
rect 100 192 101 193 
rect 100 193 101 194 
rect 100 194 101 195 
rect 100 195 101 196 
rect 100 199 101 200 
rect 100 216 101 217 
rect 100 224 101 225 
rect 100 235 101 236 
rect 100 242 101 243 
rect 100 247 101 248 
rect 100 276 101 277 
rect 100 280 101 281 
rect 100 289 101 290 
rect 100 292 101 293 
rect 100 303 101 304 
rect 100 305 101 306 
rect 100 308 101 309 
rect 100 310 101 311 
rect 100 311 101 312 
rect 101 1 102 2 
rect 101 3 102 4 
rect 101 8 102 9 
rect 101 18 102 19 
rect 101 20 102 21 
rect 101 23 102 24 
rect 101 38 102 39 
rect 101 50 102 51 
rect 101 52 102 53 
rect 101 56 102 57 
rect 101 68 102 69 
rect 101 72 102 73 
rect 101 81 102 82 
rect 101 84 102 85 
rect 101 87 102 88 
rect 101 94 102 95 
rect 101 101 102 102 
rect 101 114 102 115 
rect 101 115 102 116 
rect 101 135 102 136 
rect 101 145 102 146 
rect 101 147 102 148 
rect 101 161 102 162 
rect 101 166 102 167 
rect 101 216 102 217 
rect 101 224 102 225 
rect 101 235 102 236 
rect 101 242 102 243 
rect 101 247 102 248 
rect 101 276 102 277 
rect 101 280 102 281 
rect 101 289 102 290 
rect 101 292 102 293 
rect 101 303 102 304 
rect 101 305 102 306 
rect 101 308 102 309 
rect 101 310 102 311 
rect 101 312 102 313 
rect 101 313 102 314 
rect 102 1 103 2 
rect 102 3 103 4 
rect 102 8 103 9 
rect 102 18 103 19 
rect 102 20 103 21 
rect 102 23 103 24 
rect 102 38 103 39 
rect 102 50 103 51 
rect 102 52 103 53 
rect 102 56 103 57 
rect 102 68 103 69 
rect 102 72 103 73 
rect 102 81 103 82 
rect 102 84 103 85 
rect 102 87 103 88 
rect 102 94 103 95 
rect 102 101 103 102 
rect 102 114 103 115 
rect 102 116 103 117 
rect 102 117 103 118 
rect 102 118 103 119 
rect 102 119 103 120 
rect 102 120 103 121 
rect 102 121 103 122 
rect 102 122 103 123 
rect 102 123 103 124 
rect 102 124 103 125 
rect 102 125 103 126 
rect 102 126 103 127 
rect 102 127 103 128 
rect 102 128 103 129 
rect 102 129 103 130 
rect 102 130 103 131 
rect 102 131 103 132 
rect 102 132 103 133 
rect 102 135 103 136 
rect 102 145 103 146 
rect 102 147 103 148 
rect 102 161 103 162 
rect 102 166 103 167 
rect 102 167 103 168 
rect 102 168 103 169 
rect 102 169 103 170 
rect 102 170 103 171 
rect 102 171 103 172 
rect 102 172 103 173 
rect 102 173 103 174 
rect 102 174 103 175 
rect 102 175 103 176 
rect 102 176 103 177 
rect 102 177 103 178 
rect 102 178 103 179 
rect 102 179 103 180 
rect 102 180 103 181 
rect 102 181 103 182 
rect 102 182 103 183 
rect 102 183 103 184 
rect 102 184 103 185 
rect 102 185 103 186 
rect 102 186 103 187 
rect 102 187 103 188 
rect 102 188 103 189 
rect 102 189 103 190 
rect 102 190 103 191 
rect 102 191 103 192 
rect 102 192 103 193 
rect 102 193 103 194 
rect 102 194 103 195 
rect 102 195 103 196 
rect 102 196 103 197 
rect 102 197 103 198 
rect 102 198 103 199 
rect 102 199 103 200 
rect 102 200 103 201 
rect 102 201 103 202 
rect 102 202 103 203 
rect 102 203 103 204 
rect 102 204 103 205 
rect 102 205 103 206 
rect 102 206 103 207 
rect 102 207 103 208 
rect 102 208 103 209 
rect 102 209 103 210 
rect 102 210 103 211 
rect 102 211 103 212 
rect 102 212 103 213 
rect 102 213 103 214 
rect 102 214 103 215 
rect 102 216 103 217 
rect 102 219 103 220 
rect 102 220 103 221 
rect 102 221 103 222 
rect 102 222 103 223 
rect 102 223 103 224 
rect 102 224 103 225 
rect 102 235 103 236 
rect 102 242 103 243 
rect 102 247 103 248 
rect 102 276 103 277 
rect 102 280 103 281 
rect 102 289 103 290 
rect 102 292 103 293 
rect 102 303 103 304 
rect 102 305 103 306 
rect 102 308 103 309 
rect 102 310 103 311 
rect 102 312 103 313 
rect 103 1 104 2 
rect 103 3 104 4 
rect 103 8 104 9 
rect 103 18 104 19 
rect 103 20 104 21 
rect 103 23 104 24 
rect 103 38 104 39 
rect 103 50 104 51 
rect 103 52 104 53 
rect 103 56 104 57 
rect 103 68 104 69 
rect 103 69 104 70 
rect 103 72 104 73 
rect 103 81 104 82 
rect 103 84 104 85 
rect 103 87 104 88 
rect 103 94 104 95 
rect 103 101 104 102 
rect 103 114 104 115 
rect 103 135 104 136 
rect 103 145 104 146 
rect 103 147 104 148 
rect 103 161 104 162 
rect 103 214 104 215 
rect 103 216 104 217 
rect 103 235 104 236 
rect 103 242 104 243 
rect 103 247 104 248 
rect 103 276 104 277 
rect 103 280 104 281 
rect 103 289 104 290 
rect 103 292 104 293 
rect 103 303 104 304 
rect 103 305 104 306 
rect 103 308 104 309 
rect 103 310 104 311 
rect 103 312 104 313 
rect 104 1 105 2 
rect 104 3 105 4 
rect 104 8 105 9 
rect 104 18 105 19 
rect 104 20 105 21 
rect 104 23 105 24 
rect 104 38 105 39 
rect 104 50 105 51 
rect 104 52 105 53 
rect 104 56 105 57 
rect 104 59 105 60 
rect 104 60 105 61 
rect 104 61 105 62 
rect 104 62 105 63 
rect 104 63 105 64 
rect 104 64 105 65 
rect 104 65 105 66 
rect 104 69 105 70 
rect 104 72 105 73 
rect 104 81 105 82 
rect 104 84 105 85 
rect 104 87 105 88 
rect 104 94 105 95 
rect 104 101 105 102 
rect 104 105 105 106 
rect 104 106 105 107 
rect 104 107 105 108 
rect 104 114 105 115 
rect 104 119 105 120 
rect 104 120 105 121 
rect 104 121 105 122 
rect 104 122 105 123 
rect 104 123 105 124 
rect 104 124 105 125 
rect 104 125 105 126 
rect 104 126 105 127 
rect 104 135 105 136 
rect 104 136 105 137 
rect 104 145 105 146 
rect 104 147 105 148 
rect 104 161 105 162 
rect 104 169 105 170 
rect 104 170 105 171 
rect 104 171 105 172 
rect 104 172 105 173 
rect 104 173 105 174 
rect 104 174 105 175 
rect 104 175 105 176 
rect 104 176 105 177 
rect 104 177 105 178 
rect 104 178 105 179 
rect 104 179 105 180 
rect 104 180 105 181 
rect 104 181 105 182 
rect 104 182 105 183 
rect 104 183 105 184 
rect 104 184 105 185 
rect 104 185 105 186 
rect 104 186 105 187 
rect 104 187 105 188 
rect 104 188 105 189 
rect 104 189 105 190 
rect 104 190 105 191 
rect 104 191 105 192 
rect 104 192 105 193 
rect 104 193 105 194 
rect 104 194 105 195 
rect 104 195 105 196 
rect 104 196 105 197 
rect 104 197 105 198 
rect 104 198 105 199 
rect 104 199 105 200 
rect 104 200 105 201 
rect 104 201 105 202 
rect 104 202 105 203 
rect 104 203 105 204 
rect 104 204 105 205 
rect 104 205 105 206 
rect 104 206 105 207 
rect 104 207 105 208 
rect 104 208 105 209 
rect 104 209 105 210 
rect 104 210 105 211 
rect 104 211 105 212 
rect 104 212 105 213 
rect 104 214 105 215 
rect 104 216 105 217 
rect 104 219 105 220 
rect 104 220 105 221 
rect 104 221 105 222 
rect 104 222 105 223 
rect 104 223 105 224 
rect 104 224 105 225 
rect 104 225 105 226 
rect 104 233 105 234 
rect 104 234 105 235 
rect 104 235 105 236 
rect 104 242 105 243 
rect 104 247 105 248 
rect 104 276 105 277 
rect 104 280 105 281 
rect 104 289 105 290 
rect 104 292 105 293 
rect 104 302 105 303 
rect 104 303 105 304 
rect 104 305 105 306 
rect 104 308 105 309 
rect 104 310 105 311 
rect 104 312 105 313 
rect 105 1 106 2 
rect 105 3 106 4 
rect 105 8 106 9 
rect 105 18 106 19 
rect 105 20 106 21 
rect 105 23 106 24 
rect 105 38 106 39 
rect 105 50 106 51 
rect 105 52 106 53 
rect 105 56 106 57 
rect 105 59 106 60 
rect 105 65 106 66 
rect 105 69 106 70 
rect 105 72 106 73 
rect 105 81 106 82 
rect 105 84 106 85 
rect 105 87 106 88 
rect 105 94 106 95 
rect 105 101 106 102 
rect 105 104 106 105 
rect 105 105 106 106 
rect 105 107 106 108 
rect 105 114 106 115 
rect 105 126 106 127 
rect 105 136 106 137 
rect 105 145 106 146 
rect 105 147 106 148 
rect 105 161 106 162 
rect 105 168 106 169 
rect 105 169 106 170 
rect 105 214 106 215 
rect 105 216 106 217 
rect 105 225 106 226 
rect 105 226 106 227 
rect 105 227 106 228 
rect 105 228 106 229 
rect 105 229 106 230 
rect 105 230 106 231 
rect 105 231 106 232 
rect 105 232 106 233 
rect 105 233 106 234 
rect 105 242 106 243 
rect 105 247 106 248 
rect 105 276 106 277 
rect 105 280 106 281 
rect 105 289 106 290 
rect 105 292 106 293 
rect 105 302 106 303 
rect 105 305 106 306 
rect 105 308 106 309 
rect 105 310 106 311 
rect 105 312 106 313 
rect 106 1 107 2 
rect 106 3 107 4 
rect 106 8 107 9 
rect 106 18 107 19 
rect 106 20 107 21 
rect 106 23 107 24 
rect 106 38 107 39 
rect 106 50 107 51 
rect 106 52 107 53 
rect 106 56 107 57 
rect 106 59 107 60 
rect 106 65 107 66 
rect 106 69 107 70 
rect 106 72 107 73 
rect 106 81 107 82 
rect 106 84 107 85 
rect 106 87 107 88 
rect 106 94 107 95 
rect 106 101 107 102 
rect 106 102 107 103 
rect 106 104 107 105 
rect 106 107 107 108 
rect 106 114 107 115 
rect 106 126 107 127 
rect 106 136 107 137 
rect 106 145 107 146 
rect 106 147 107 148 
rect 106 161 107 162 
rect 106 168 107 169 
rect 106 194 107 195 
rect 106 214 107 215 
rect 106 216 107 217 
rect 106 242 107 243 
rect 106 247 107 248 
rect 106 276 107 277 
rect 106 280 107 281 
rect 106 289 107 290 
rect 106 292 107 293 
rect 106 302 107 303 
rect 106 305 107 306 
rect 106 308 107 309 
rect 106 310 107 311 
rect 106 312 107 313 
rect 107 1 108 2 
rect 107 3 108 4 
rect 107 8 108 9 
rect 107 18 108 19 
rect 107 20 108 21 
rect 107 23 108 24 
rect 107 38 108 39 
rect 107 50 108 51 
rect 107 52 108 53 
rect 107 56 108 57 
rect 107 65 108 66 
rect 107 69 108 70 
rect 107 72 108 73 
rect 107 81 108 82 
rect 107 84 108 85 
rect 107 87 108 88 
rect 107 102 108 103 
rect 107 104 108 105 
rect 107 114 108 115 
rect 107 136 108 137 
rect 107 145 108 146 
rect 107 147 108 148 
rect 107 161 108 162 
rect 107 168 108 169 
rect 107 194 108 195 
rect 107 214 108 215 
rect 107 216 108 217 
rect 107 242 108 243 
rect 107 247 108 248 
rect 107 276 108 277 
rect 107 280 108 281 
rect 107 289 108 290 
rect 107 292 108 293 
rect 107 305 108 306 
rect 107 308 108 309 
rect 107 310 108 311 
rect 107 312 108 313 
rect 108 1 109 2 
rect 108 3 109 4 
rect 108 8 109 9 
rect 108 18 109 19 
rect 108 20 109 21 
rect 108 23 109 24 
rect 108 38 109 39 
rect 108 50 109 51 
rect 108 52 109 53 
rect 108 56 109 57 
rect 108 65 109 66 
rect 108 69 109 70 
rect 108 72 109 73 
rect 108 81 109 82 
rect 108 84 109 85 
rect 108 87 109 88 
rect 108 102 109 103 
rect 108 104 109 105 
rect 108 114 109 115 
rect 108 136 109 137 
rect 108 145 109 146 
rect 108 147 109 148 
rect 108 161 109 162 
rect 108 168 109 169 
rect 108 194 109 195 
rect 108 214 109 215 
rect 108 216 109 217 
rect 108 242 109 243 
rect 108 247 109 248 
rect 108 276 109 277 
rect 108 280 109 281 
rect 108 289 109 290 
rect 108 292 109 293 
rect 108 305 109 306 
rect 108 308 109 309 
rect 108 310 109 311 
rect 108 312 109 313 
rect 109 1 110 2 
rect 109 3 110 4 
rect 109 8 110 9 
rect 109 18 110 19 
rect 109 20 110 21 
rect 109 23 110 24 
rect 109 38 110 39 
rect 109 50 110 51 
rect 109 52 110 53 
rect 109 56 110 57 
rect 109 65 110 66 
rect 109 69 110 70 
rect 109 72 110 73 
rect 109 81 110 82 
rect 109 84 110 85 
rect 109 87 110 88 
rect 109 102 110 103 
rect 109 104 110 105 
rect 109 114 110 115 
rect 109 136 110 137 
rect 109 145 110 146 
rect 109 147 110 148 
rect 109 161 110 162 
rect 109 166 110 167 
rect 109 167 110 168 
rect 109 168 110 169 
rect 109 194 110 195 
rect 109 214 110 215 
rect 109 216 110 217 
rect 109 242 110 243 
rect 109 247 110 248 
rect 109 276 110 277 
rect 109 280 110 281 
rect 109 289 110 290 
rect 109 292 110 293 
rect 109 305 110 306 
rect 109 308 110 309 
rect 109 310 110 311 
rect 109 312 110 313 
rect 110 1 111 2 
rect 110 3 111 4 
rect 110 8 111 9 
rect 110 18 111 19 
rect 110 20 111 21 
rect 110 23 111 24 
rect 110 38 111 39 
rect 110 50 111 51 
rect 110 52 111 53 
rect 110 56 111 57 
rect 110 65 111 66 
rect 110 69 111 70 
rect 110 72 111 73 
rect 110 81 111 82 
rect 110 84 111 85 
rect 110 87 111 88 
rect 110 102 111 103 
rect 110 104 111 105 
rect 110 114 111 115 
rect 110 136 111 137 
rect 110 145 111 146 
rect 110 147 111 148 
rect 110 149 111 150 
rect 110 150 111 151 
rect 110 151 111 152 
rect 110 152 111 153 
rect 110 161 111 162 
rect 110 166 111 167 
rect 110 194 111 195 
rect 110 214 111 215 
rect 110 216 111 217 
rect 110 242 111 243 
rect 110 247 111 248 
rect 110 276 111 277 
rect 110 280 111 281 
rect 110 289 111 290 
rect 110 292 111 293 
rect 110 305 111 306 
rect 110 308 111 309 
rect 110 310 111 311 
rect 110 312 111 313 
rect 111 1 112 2 
rect 111 3 112 4 
rect 111 8 112 9 
rect 111 18 112 19 
rect 111 20 112 21 
rect 111 23 112 24 
rect 111 27 112 28 
rect 111 38 112 39 
rect 111 50 112 51 
rect 111 52 112 53 
rect 111 56 112 57 
rect 111 65 112 66 
rect 111 69 112 70 
rect 111 72 112 73 
rect 111 75 112 76 
rect 111 81 112 82 
rect 111 84 112 85 
rect 111 87 112 88 
rect 111 102 112 103 
rect 111 104 112 105 
rect 111 114 112 115 
rect 111 136 112 137 
rect 111 145 112 146 
rect 111 147 112 148 
rect 111 152 112 153 
rect 111 158 112 159 
rect 111 161 112 162 
rect 111 166 112 167 
rect 111 171 112 172 
rect 111 174 112 175 
rect 111 177 112 178 
rect 111 178 112 179 
rect 111 179 112 180 
rect 111 180 112 181 
rect 111 181 112 182 
rect 111 194 112 195 
rect 111 206 112 207 
rect 111 214 112 215 
rect 111 216 112 217 
rect 111 222 112 223 
rect 111 241 112 242 
rect 111 242 112 243 
rect 111 247 112 248 
rect 111 251 112 252 
rect 111 270 112 271 
rect 111 276 112 277 
rect 111 280 112 281 
rect 111 289 112 290 
rect 111 292 112 293 
rect 111 302 112 303 
rect 111 305 112 306 
rect 111 308 112 309 
rect 111 310 112 311 
rect 111 312 112 313 
rect 112 1 113 2 
rect 112 3 113 4 
rect 112 8 113 9 
rect 112 18 113 19 
rect 112 20 113 21 
rect 112 23 113 24 
rect 112 27 113 28 
rect 112 38 113 39 
rect 112 50 113 51 
rect 112 52 113 53 
rect 112 56 113 57 
rect 112 65 113 66 
rect 112 72 113 73 
rect 112 73 113 74 
rect 112 75 113 76 
rect 112 80 113 81 
rect 112 81 113 82 
rect 112 84 113 85 
rect 112 87 113 88 
rect 112 102 113 103 
rect 112 104 113 105 
rect 112 114 113 115 
rect 112 136 113 137 
rect 112 144 113 145 
rect 112 145 113 146 
rect 112 147 113 148 
rect 112 152 113 153 
rect 112 158 113 159 
rect 112 161 113 162 
rect 112 166 113 167 
rect 112 171 113 172 
rect 112 174 113 175 
rect 112 176 113 177 
rect 112 177 113 178 
rect 112 194 113 195 
rect 112 206 113 207 
rect 112 214 113 215 
rect 112 216 113 217 
rect 112 217 113 218 
rect 112 222 113 223 
rect 112 247 113 248 
rect 112 251 113 252 
rect 112 270 113 271 
rect 112 276 113 277 
rect 112 280 113 281 
rect 112 289 113 290 
rect 112 292 113 293 
rect 112 302 113 303 
rect 112 305 113 306 
rect 112 308 113 309 
rect 112 310 113 311 
rect 112 312 113 313 
rect 113 1 114 2 
rect 113 3 114 4 
rect 113 8 114 9 
rect 113 18 114 19 
rect 113 20 114 21 
rect 113 23 114 24 
rect 113 27 114 28 
rect 113 28 114 29 
rect 113 29 114 30 
rect 113 30 114 31 
rect 113 31 114 32 
rect 113 32 114 33 
rect 113 33 114 34 
rect 113 34 114 35 
rect 113 35 114 36 
rect 113 36 114 37 
rect 113 38 114 39 
rect 113 50 114 51 
rect 113 52 114 53 
rect 113 56 114 57 
rect 113 65 114 66 
rect 113 66 114 67 
rect 113 67 114 68 
rect 113 68 114 69 
rect 113 69 114 70 
rect 113 70 114 71 
rect 113 73 114 74 
rect 113 74 114 75 
rect 113 75 114 76 
rect 113 77 114 78 
rect 113 78 114 79 
rect 113 79 114 80 
rect 113 80 114 81 
rect 113 84 114 85 
rect 113 87 114 88 
rect 113 102 114 103 
rect 113 104 114 105 
rect 113 114 114 115 
rect 113 115 114 116 
rect 113 116 114 117 
rect 113 117 114 118 
rect 113 118 114 119 
rect 113 119 114 120 
rect 113 120 114 121 
rect 113 121 114 122 
rect 113 122 114 123 
rect 113 123 114 124 
rect 113 136 114 137 
rect 113 138 114 139 
rect 113 139 114 140 
rect 113 140 114 141 
rect 113 141 114 142 
rect 113 142 114 143 
rect 113 143 114 144 
rect 113 144 114 145 
rect 113 146 114 147 
rect 113 147 114 148 
rect 113 152 114 153 
rect 113 153 114 154 
rect 113 154 114 155 
rect 113 155 114 156 
rect 113 156 114 157 
rect 113 157 114 158 
rect 113 158 114 159 
rect 113 161 114 162 
rect 113 166 114 167 
rect 113 171 114 172 
rect 113 174 114 175 
rect 113 175 114 176 
rect 113 176 114 177 
rect 113 194 114 195 
rect 113 206 114 207 
rect 113 214 114 215 
rect 113 215 114 216 
rect 113 217 114 218 
rect 113 218 114 219 
rect 113 219 114 220 
rect 113 220 114 221 
rect 113 221 114 222 
rect 113 222 114 223 
rect 113 224 114 225 
rect 113 225 114 226 
rect 113 226 114 227 
rect 113 227 114 228 
rect 113 228 114 229 
rect 113 229 114 230 
rect 113 230 114 231 
rect 113 231 114 232 
rect 113 232 114 233 
rect 113 233 114 234 
rect 113 234 114 235 
rect 113 235 114 236 
rect 113 236 114 237 
rect 113 237 114 238 
rect 113 238 114 239 
rect 113 239 114 240 
rect 113 240 114 241 
rect 113 241 114 242 
rect 113 242 114 243 
rect 113 243 114 244 
rect 113 244 114 245 
rect 113 247 114 248 
rect 113 249 114 250 
rect 113 250 114 251 
rect 113 251 114 252 
rect 113 257 114 258 
rect 113 258 114 259 
rect 113 259 114 260 
rect 113 260 114 261 
rect 113 261 114 262 
rect 113 262 114 263 
rect 113 263 114 264 
rect 113 264 114 265 
rect 113 265 114 266 
rect 113 266 114 267 
rect 113 267 114 268 
rect 113 268 114 269 
rect 113 269 114 270 
rect 113 270 114 271 
rect 113 276 114 277 
rect 113 280 114 281 
rect 113 282 114 283 
rect 113 289 114 290 
rect 113 292 114 293 
rect 113 297 114 298 
rect 113 298 114 299 
rect 113 299 114 300 
rect 113 300 114 301 
rect 113 301 114 302 
rect 113 302 114 303 
rect 113 305 114 306 
rect 113 308 114 309 
rect 113 310 114 311 
rect 113 312 114 313 
rect 114 1 115 2 
rect 114 3 115 4 
rect 114 8 115 9 
rect 114 18 115 19 
rect 114 20 115 21 
rect 114 23 115 24 
rect 114 76 115 77 
rect 114 77 115 78 
rect 114 84 115 85 
rect 114 87 115 88 
rect 114 102 115 103 
rect 114 104 115 105 
rect 114 123 115 124 
rect 114 134 115 135 
rect 114 136 115 137 
rect 114 145 115 146 
rect 114 146 115 147 
rect 114 161 115 162 
rect 114 165 115 166 
rect 114 166 115 167 
rect 114 171 115 172 
rect 114 194 115 195 
rect 114 206 115 207 
rect 114 215 115 216 
rect 114 216 115 217 
rect 114 247 115 248 
rect 114 257 115 258 
rect 114 276 115 277 
rect 114 280 115 281 
rect 114 282 115 283 
rect 114 289 115 290 
rect 114 292 115 293 
rect 114 297 115 298 
rect 114 305 115 306 
rect 114 308 115 309 
rect 114 310 115 311 
rect 114 312 115 313 
rect 115 1 116 2 
rect 115 3 116 4 
rect 115 8 116 9 
rect 115 18 116 19 
rect 115 20 116 21 
rect 115 23 116 24 
rect 115 25 116 26 
rect 115 26 116 27 
rect 115 27 116 28 
rect 115 28 116 29 
rect 115 29 116 30 
rect 115 30 116 31 
rect 115 31 116 32 
rect 115 32 116 33 
rect 115 33 116 34 
rect 115 34 116 35 
rect 115 35 116 36 
rect 115 36 116 37 
rect 115 37 116 38 
rect 115 38 116 39 
rect 115 39 116 40 
rect 115 40 116 41 
rect 115 41 116 42 
rect 115 42 116 43 
rect 115 43 116 44 
rect 115 44 116 45 
rect 115 45 116 46 
rect 115 46 116 47 
rect 115 47 116 48 
rect 115 48 116 49 
rect 115 49 116 50 
rect 115 50 116 51 
rect 115 51 116 52 
rect 115 52 116 53 
rect 115 53 116 54 
rect 115 54 116 55 
rect 115 55 116 56 
rect 115 56 116 57 
rect 115 57 116 58 
rect 115 58 116 59 
rect 115 59 116 60 
rect 115 60 116 61 
rect 115 61 116 62 
rect 115 62 116 63 
rect 115 63 116 64 
rect 115 64 116 65 
rect 115 65 116 66 
rect 115 66 116 67 
rect 115 67 116 68 
rect 115 68 116 69 
rect 115 69 116 70 
rect 115 70 116 71 
rect 115 71 116 72 
rect 115 72 116 73 
rect 115 73 116 74 
rect 115 74 116 75 
rect 115 75 116 76 
rect 115 76 116 77 
rect 115 86 116 87 
rect 115 87 116 88 
rect 115 102 116 103 
rect 115 104 116 105 
rect 115 123 116 124 
rect 115 134 116 135 
rect 115 136 116 137 
rect 115 138 116 139 
rect 115 139 116 140 
rect 115 140 116 141 
rect 115 141 116 142 
rect 115 142 116 143 
rect 115 143 116 144 
rect 115 144 116 145 
rect 115 145 116 146 
rect 115 161 116 162 
rect 115 165 116 166 
rect 115 171 116 172 
rect 115 194 116 195 
rect 115 206 116 207 
rect 115 216 116 217 
rect 115 217 116 218 
rect 115 218 116 219 
rect 115 219 116 220 
rect 115 220 116 221 
rect 115 221 116 222 
rect 115 222 116 223 
rect 115 223 116 224 
rect 115 224 116 225 
rect 115 225 116 226 
rect 115 226 116 227 
rect 115 227 116 228 
rect 115 228 116 229 
rect 115 229 116 230 
rect 115 230 116 231 
rect 115 231 116 232 
rect 115 232 116 233 
rect 115 233 116 234 
rect 115 234 116 235 
rect 115 235 116 236 
rect 115 236 116 237 
rect 115 237 116 238 
rect 115 238 116 239 
rect 115 239 116 240 
rect 115 240 116 241 
rect 115 241 116 242 
rect 115 242 116 243 
rect 115 243 116 244 
rect 115 244 116 245 
rect 115 245 116 246 
rect 115 247 116 248 
rect 115 250 116 251 
rect 115 251 116 252 
rect 115 257 116 258 
rect 115 260 116 261 
rect 115 276 116 277 
rect 115 280 116 281 
rect 115 282 116 283 
rect 115 289 116 290 
rect 115 292 116 293 
rect 115 297 116 298 
rect 115 305 116 306 
rect 115 308 116 309 
rect 115 310 116 311 
rect 115 312 116 313 
rect 116 1 117 2 
rect 116 3 117 4 
rect 116 8 117 9 
rect 116 16 117 17 
rect 116 18 117 19 
rect 116 20 117 21 
rect 116 23 117 24 
rect 116 102 117 103 
rect 116 104 117 105 
rect 116 123 117 124 
rect 116 132 117 133 
rect 116 134 117 135 
rect 116 136 117 137 
rect 116 161 117 162 
rect 116 165 117 166 
rect 116 171 117 172 
rect 116 194 117 195 
rect 116 206 117 207 
rect 116 247 117 248 
rect 116 251 117 252 
rect 116 252 117 253 
rect 116 253 117 254 
rect 116 254 117 255 
rect 116 255 117 256 
rect 116 256 117 257 
rect 116 257 117 258 
rect 116 260 117 261 
rect 116 262 117 263 
rect 116 263 117 264 
rect 116 276 117 277 
rect 116 280 117 281 
rect 116 282 117 283 
rect 116 289 117 290 
rect 116 292 117 293 
rect 116 297 117 298 
rect 116 305 117 306 
rect 116 308 117 309 
rect 116 310 117 311 
rect 116 312 117 313 
rect 117 1 118 2 
rect 117 3 118 4 
rect 117 8 118 9 
rect 117 16 118 17 
rect 117 18 118 19 
rect 117 20 118 21 
rect 117 23 118 24 
rect 117 37 118 38 
rect 117 38 118 39 
rect 117 39 118 40 
rect 117 40 118 41 
rect 117 41 118 42 
rect 117 42 118 43 
rect 117 43 118 44 
rect 117 44 118 45 
rect 117 45 118 46 
rect 117 46 118 47 
rect 117 47 118 48 
rect 117 48 118 49 
rect 117 49 118 50 
rect 117 50 118 51 
rect 117 51 118 52 
rect 117 52 118 53 
rect 117 53 118 54 
rect 117 54 118 55 
rect 117 55 118 56 
rect 117 56 118 57 
rect 117 57 118 58 
rect 117 58 118 59 
rect 117 59 118 60 
rect 117 60 118 61 
rect 117 61 118 62 
rect 117 62 118 63 
rect 117 63 118 64 
rect 117 64 118 65 
rect 117 65 118 66 
rect 117 66 118 67 
rect 117 67 118 68 
rect 117 68 118 69 
rect 117 69 118 70 
rect 117 70 118 71 
rect 117 71 118 72 
rect 117 72 118 73 
rect 117 73 118 74 
rect 117 74 118 75 
rect 117 75 118 76 
rect 117 76 118 77 
rect 117 77 118 78 
rect 117 78 118 79 
rect 117 79 118 80 
rect 117 80 118 81 
rect 117 81 118 82 
rect 117 82 118 83 
rect 117 83 118 84 
rect 117 84 118 85 
rect 117 85 118 86 
rect 117 86 118 87 
rect 117 87 118 88 
rect 117 88 118 89 
rect 117 89 118 90 
rect 117 90 118 91 
rect 117 91 118 92 
rect 117 92 118 93 
rect 117 93 118 94 
rect 117 94 118 95 
rect 117 95 118 96 
rect 117 96 118 97 
rect 117 97 118 98 
rect 117 102 118 103 
rect 117 104 118 105 
rect 117 123 118 124 
rect 117 132 118 133 
rect 117 134 118 135 
rect 117 136 118 137 
rect 117 161 118 162 
rect 117 165 118 166 
rect 117 171 118 172 
rect 117 172 118 173 
rect 117 173 118 174 
rect 117 174 118 175 
rect 117 175 118 176 
rect 117 176 118 177 
rect 117 177 118 178 
rect 117 178 118 179 
rect 117 179 118 180 
rect 117 180 118 181 
rect 117 194 118 195 
rect 117 195 118 196 
rect 117 206 118 207 
rect 117 207 118 208 
rect 117 208 118 209 
rect 117 209 118 210 
rect 117 210 118 211 
rect 117 211 118 212 
rect 117 212 118 213 
rect 117 213 118 214 
rect 117 214 118 215 
rect 117 215 118 216 
rect 117 216 118 217 
rect 117 217 118 218 
rect 117 218 118 219 
rect 117 219 118 220 
rect 117 220 118 221 
rect 117 221 118 222 
rect 117 222 118 223 
rect 117 223 118 224 
rect 117 224 118 225 
rect 117 225 118 226 
rect 117 231 118 232 
rect 117 232 118 233 
rect 117 233 118 234 
rect 117 234 118 235 
rect 117 235 118 236 
rect 117 236 118 237 
rect 117 237 118 238 
rect 117 238 118 239 
rect 117 239 118 240 
rect 117 240 118 241 
rect 117 241 118 242 
rect 117 242 118 243 
rect 117 243 118 244 
rect 117 244 118 245 
rect 117 245 118 246 
rect 117 246 118 247 
rect 117 247 118 248 
rect 117 260 118 261 
rect 117 262 118 263 
rect 117 276 118 277 
rect 117 280 118 281 
rect 117 282 118 283 
rect 117 283 118 284 
rect 117 289 118 290 
rect 117 292 118 293 
rect 117 297 118 298 
rect 117 305 118 306 
rect 117 308 118 309 
rect 117 310 118 311 
rect 117 312 118 313 
rect 118 1 119 2 
rect 118 3 119 4 
rect 118 8 119 9 
rect 118 16 119 17 
rect 118 18 119 19 
rect 118 20 119 21 
rect 118 23 119 24 
rect 118 123 119 124 
rect 118 131 119 132 
rect 118 132 119 133 
rect 118 134 119 135 
rect 118 136 119 137 
rect 118 161 119 162 
rect 118 165 119 166 
rect 118 230 119 231 
rect 118 231 119 232 
rect 118 260 119 261 
rect 118 262 119 263 
rect 118 280 119 281 
rect 118 283 119 284 
rect 118 284 119 285 
rect 118 289 119 290 
rect 118 292 119 293 
rect 118 297 119 298 
rect 118 305 119 306 
rect 118 308 119 309 
rect 118 310 119 311 
rect 118 312 119 313 
rect 119 1 120 2 
rect 119 3 120 4 
rect 119 8 120 9 
rect 119 11 120 12 
rect 119 12 120 13 
rect 119 13 120 14 
rect 119 14 120 15 
rect 119 15 120 16 
rect 119 16 120 17 
rect 119 18 120 19 
rect 119 20 120 21 
rect 119 23 120 24 
rect 119 30 120 31 
rect 119 31 120 32 
rect 119 32 120 33 
rect 119 33 120 34 
rect 119 34 120 35 
rect 119 35 120 36 
rect 119 36 120 37 
rect 119 37 120 38 
rect 119 38 120 39 
rect 119 39 120 40 
rect 119 40 120 41 
rect 119 41 120 42 
rect 119 42 120 43 
rect 119 43 120 44 
rect 119 44 120 45 
rect 119 45 120 46 
rect 119 46 120 47 
rect 119 47 120 48 
rect 119 48 120 49 
rect 119 49 120 50 
rect 119 50 120 51 
rect 119 51 120 52 
rect 119 52 120 53 
rect 119 53 120 54 
rect 119 54 120 55 
rect 119 55 120 56 
rect 119 56 120 57 
rect 119 57 120 58 
rect 119 58 120 59 
rect 119 59 120 60 
rect 119 60 120 61 
rect 119 61 120 62 
rect 119 62 120 63 
rect 119 63 120 64 
rect 119 64 120 65 
rect 119 65 120 66 
rect 119 66 120 67 
rect 119 67 120 68 
rect 119 68 120 69 
rect 119 69 120 70 
rect 119 70 120 71 
rect 119 71 120 72 
rect 119 72 120 73 
rect 119 73 120 74 
rect 119 74 120 75 
rect 119 75 120 76 
rect 119 76 120 77 
rect 119 77 120 78 
rect 119 78 120 79 
rect 119 79 120 80 
rect 119 80 120 81 
rect 119 81 120 82 
rect 119 82 120 83 
rect 119 83 120 84 
rect 119 84 120 85 
rect 119 85 120 86 
rect 119 86 120 87 
rect 119 87 120 88 
rect 119 88 120 89 
rect 119 89 120 90 
rect 119 90 120 91 
rect 119 91 120 92 
rect 119 92 120 93 
rect 119 93 120 94 
rect 119 94 120 95 
rect 119 95 120 96 
rect 119 96 120 97 
rect 119 97 120 98 
rect 119 98 120 99 
rect 119 99 120 100 
rect 119 100 120 101 
rect 119 101 120 102 
rect 119 102 120 103 
rect 119 103 120 104 
rect 119 104 120 105 
rect 119 105 120 106 
rect 119 106 120 107 
rect 119 107 120 108 
rect 119 108 120 109 
rect 119 109 120 110 
rect 119 110 120 111 
rect 119 111 120 112 
rect 119 123 120 124 
rect 119 130 120 131 
rect 119 131 120 132 
rect 119 133 120 134 
rect 119 134 120 135 
rect 119 136 120 137 
rect 119 140 120 141 
rect 119 141 120 142 
rect 119 142 120 143 
rect 119 143 120 144 
rect 119 144 120 145 
rect 119 145 120 146 
rect 119 146 120 147 
rect 119 147 120 148 
rect 119 161 120 162 
rect 119 165 120 166 
rect 119 168 120 169 
rect 119 169 120 170 
rect 119 170 120 171 
rect 119 171 120 172 
rect 119 172 120 173 
rect 119 173 120 174 
rect 119 174 120 175 
rect 119 175 120 176 
rect 119 176 120 177 
rect 119 177 120 178 
rect 119 178 120 179 
rect 119 179 120 180 
rect 119 180 120 181 
rect 119 181 120 182 
rect 119 182 120 183 
rect 119 183 120 184 
rect 119 184 120 185 
rect 119 185 120 186 
rect 119 186 120 187 
rect 119 187 120 188 
rect 119 188 120 189 
rect 119 189 120 190 
rect 119 190 120 191 
rect 119 191 120 192 
rect 119 192 120 193 
rect 119 193 120 194 
rect 119 194 120 195 
rect 119 195 120 196 
rect 119 196 120 197 
rect 119 197 120 198 
rect 119 198 120 199 
rect 119 199 120 200 
rect 119 200 120 201 
rect 119 201 120 202 
rect 119 202 120 203 
rect 119 203 120 204 
rect 119 204 120 205 
rect 119 205 120 206 
rect 119 206 120 207 
rect 119 207 120 208 
rect 119 208 120 209 
rect 119 209 120 210 
rect 119 210 120 211 
rect 119 211 120 212 
rect 119 212 120 213 
rect 119 213 120 214 
rect 119 214 120 215 
rect 119 215 120 216 
rect 119 216 120 217 
rect 119 217 120 218 
rect 119 218 120 219 
rect 119 219 120 220 
rect 119 220 120 221 
rect 119 221 120 222 
rect 119 222 120 223 
rect 119 223 120 224 
rect 119 224 120 225 
rect 119 225 120 226 
rect 119 226 120 227 
rect 119 227 120 228 
rect 119 228 120 229 
rect 119 229 120 230 
rect 119 230 120 231 
rect 119 232 120 233 
rect 119 233 120 234 
rect 119 234 120 235 
rect 119 235 120 236 
rect 119 236 120 237 
rect 119 237 120 238 
rect 119 238 120 239 
rect 119 239 120 240 
rect 119 240 120 241 
rect 119 241 120 242 
rect 119 242 120 243 
rect 119 243 120 244 
rect 119 244 120 245 
rect 119 245 120 246 
rect 119 246 120 247 
rect 119 247 120 248 
rect 119 248 120 249 
rect 119 249 120 250 
rect 119 250 120 251 
rect 119 251 120 252 
rect 119 252 120 253 
rect 119 253 120 254 
rect 119 260 120 261 
rect 119 262 120 263 
rect 119 276 120 277 
rect 119 277 120 278 
rect 119 280 120 281 
rect 119 282 120 283 
rect 119 284 120 285 
rect 119 285 120 286 
rect 119 286 120 287 
rect 119 289 120 290 
rect 119 292 120 293 
rect 119 294 120 295 
rect 119 295 120 296 
rect 119 296 120 297 
rect 119 297 120 298 
rect 119 305 120 306 
rect 119 308 120 309 
rect 119 310 120 311 
rect 119 312 120 313 
rect 120 1 121 2 
rect 120 3 121 4 
rect 120 8 121 9 
rect 120 11 121 12 
rect 120 18 121 19 
rect 120 20 121 21 
rect 120 23 121 24 
rect 120 30 121 31 
rect 120 111 121 112 
rect 120 112 121 113 
rect 120 123 121 124 
rect 120 130 121 131 
rect 120 133 121 134 
rect 120 136 121 137 
rect 120 139 121 140 
rect 120 140 121 141 
rect 120 147 121 148 
rect 120 161 121 162 
rect 120 165 121 166 
rect 120 168 121 169 
rect 120 232 121 233 
rect 120 253 121 254 
rect 120 254 121 255 
rect 120 260 121 261 
rect 120 262 121 263 
rect 120 276 121 277 
rect 120 280 121 281 
rect 120 282 121 283 
rect 120 283 121 284 
rect 120 286 121 287 
rect 120 289 121 290 
rect 120 292 121 293 
rect 120 294 121 295 
rect 120 305 121 306 
rect 120 308 121 309 
rect 120 310 121 311 
rect 120 312 121 313 
rect 121 1 122 2 
rect 121 3 122 4 
rect 121 8 122 9 
rect 121 11 122 12 
rect 121 18 122 19 
rect 121 20 122 21 
rect 121 23 122 24 
rect 121 30 122 31 
rect 121 49 122 50 
rect 121 70 122 71 
rect 121 112 122 113 
rect 121 113 122 114 
rect 121 123 122 124 
rect 121 130 122 131 
rect 121 133 122 134 
rect 121 136 122 137 
rect 121 139 122 140 
rect 121 147 122 148 
rect 121 161 122 162 
rect 121 165 122 166 
rect 121 168 122 169 
rect 121 181 122 182 
rect 121 194 122 195 
rect 121 197 122 198 
rect 121 232 122 233 
rect 121 254 122 255 
rect 121 260 122 261 
rect 121 262 122 263 
rect 121 276 122 277 
rect 121 280 122 281 
rect 121 283 122 284 
rect 121 286 122 287 
rect 121 289 122 290 
rect 121 292 122 293 
rect 121 294 122 295 
rect 121 305 122 306 
rect 121 308 122 309 
rect 121 310 122 311 
rect 121 312 122 313 
rect 122 1 123 2 
rect 122 3 123 4 
rect 122 8 123 9 
rect 122 11 123 12 
rect 122 18 123 19 
rect 122 20 123 21 
rect 122 23 123 24 
rect 122 30 123 31 
rect 122 49 123 50 
rect 122 70 123 71 
rect 122 113 123 114 
rect 122 123 123 124 
rect 122 130 123 131 
rect 122 133 123 134 
rect 122 136 123 137 
rect 122 139 123 140 
rect 122 147 123 148 
rect 122 161 123 162 
rect 122 165 123 166 
rect 122 168 123 169 
rect 122 181 123 182 
rect 122 194 123 195 
rect 122 197 123 198 
rect 122 228 123 229 
rect 122 232 123 233 
rect 122 241 123 242 
rect 122 243 123 244 
rect 122 254 123 255 
rect 122 260 123 261 
rect 122 262 123 263 
rect 122 276 123 277 
rect 122 280 123 281 
rect 122 283 123 284 
rect 122 286 123 287 
rect 122 289 123 290 
rect 122 292 123 293 
rect 122 294 123 295 
rect 122 305 123 306 
rect 122 308 123 309 
rect 122 310 123 311 
rect 122 312 123 313 
rect 123 1 124 2 
rect 123 3 124 4 
rect 123 8 124 9 
rect 123 17 124 18 
rect 123 18 124 19 
rect 123 20 124 21 
rect 123 23 124 24 
rect 123 49 124 50 
rect 123 70 124 71 
rect 123 71 124 72 
rect 123 72 124 73 
rect 123 113 124 114 
rect 123 129 124 130 
rect 123 130 124 131 
rect 123 132 124 133 
rect 123 133 124 134 
rect 123 136 124 137 
rect 123 147 124 148 
rect 123 148 124 149 
rect 123 149 124 150 
rect 123 150 124 151 
rect 123 151 124 152 
rect 123 152 124 153 
rect 123 161 124 162 
rect 123 165 124 166 
rect 123 166 124 167 
rect 123 168 124 169 
rect 123 181 124 182 
rect 123 194 124 195 
rect 123 197 124 198 
rect 123 198 124 199 
rect 123 199 124 200 
rect 123 200 124 201 
rect 123 228 124 229 
rect 123 232 124 233 
rect 123 241 124 242 
rect 123 243 124 244 
rect 123 257 124 258 
rect 123 258 124 259 
rect 123 259 124 260 
rect 123 260 124 261 
rect 123 262 124 263 
rect 123 273 124 274 
rect 123 274 124 275 
rect 123 275 124 276 
rect 123 276 124 277 
rect 123 280 124 281 
rect 123 289 124 290 
rect 123 291 124 292 
rect 123 292 124 293 
rect 123 294 124 295 
rect 123 305 124 306 
rect 123 308 124 309 
rect 123 310 124 311 
rect 123 312 124 313 
rect 124 1 125 2 
rect 124 3 125 4 
rect 124 8 125 9 
rect 124 17 125 18 
rect 124 20 125 21 
rect 124 23 125 24 
rect 124 49 125 50 
rect 124 72 125 73 
rect 124 113 125 114 
rect 124 129 125 130 
rect 124 132 125 133 
rect 124 136 125 137 
rect 124 152 125 153 
rect 124 161 125 162 
rect 124 166 125 167 
rect 124 168 125 169 
rect 124 181 125 182 
rect 124 194 125 195 
rect 124 200 125 201 
rect 124 228 125 229 
rect 124 232 125 233 
rect 124 241 125 242 
rect 124 243 125 244 
rect 124 257 125 258 
rect 124 261 125 262 
rect 124 262 125 263 
rect 124 273 125 274 
rect 124 280 125 281 
rect 124 289 125 290 
rect 124 291 125 292 
rect 124 293 125 294 
rect 124 294 125 295 
rect 124 305 125 306 
rect 124 308 125 309 
rect 124 310 125 311 
rect 124 312 125 313 
rect 125 1 126 2 
rect 125 3 126 4 
rect 125 8 126 9 
rect 125 17 126 18 
rect 125 20 126 21 
rect 125 23 126 24 
rect 125 49 126 50 
rect 125 72 126 73 
rect 125 113 126 114 
rect 125 129 126 130 
rect 125 132 126 133 
rect 125 136 126 137 
rect 125 152 126 153 
rect 125 161 126 162 
rect 125 168 126 169 
rect 125 181 126 182 
rect 125 194 126 195 
rect 125 200 126 201 
rect 125 228 126 229 
rect 125 232 126 233 
rect 125 241 126 242 
rect 125 243 126 244 
rect 125 257 126 258 
rect 125 261 126 262 
rect 125 273 126 274 
rect 125 280 126 281 
rect 125 289 126 290 
rect 125 291 126 292 
rect 125 305 126 306 
rect 125 308 126 309 
rect 125 310 126 311 
rect 125 312 126 313 
rect 126 1 127 2 
rect 126 3 127 4 
rect 126 8 127 9 
rect 126 17 127 18 
rect 126 20 127 21 
rect 126 23 127 24 
rect 126 49 127 50 
rect 126 72 127 73 
rect 126 113 127 114 
rect 126 129 127 130 
rect 126 132 127 133 
rect 126 136 127 137 
rect 126 152 127 153 
rect 126 161 127 162 
rect 126 168 127 169 
rect 126 181 127 182 
rect 126 194 127 195 
rect 126 200 127 201 
rect 126 228 127 229 
rect 126 232 127 233 
rect 126 241 127 242 
rect 126 243 127 244 
rect 126 257 127 258 
rect 126 261 127 262 
rect 126 273 127 274 
rect 126 280 127 281 
rect 126 289 127 290 
rect 126 291 127 292 
rect 126 305 127 306 
rect 126 308 127 309 
rect 126 310 127 311 
rect 126 312 127 313 
rect 127 1 128 2 
rect 127 3 128 4 
rect 127 8 128 9 
rect 127 14 128 15 
rect 127 17 128 18 
rect 127 20 128 21 
rect 127 23 128 24 
rect 127 49 128 50 
rect 127 72 128 73 
rect 127 113 128 114 
rect 127 129 128 130 
rect 127 132 128 133 
rect 127 136 128 137 
rect 127 139 128 140 
rect 127 152 128 153 
rect 127 161 128 162 
rect 127 164 128 165 
rect 127 165 128 166 
rect 127 166 128 167 
rect 127 167 128 168 
rect 127 168 128 169 
rect 127 181 128 182 
rect 127 182 128 183 
rect 127 183 128 184 
rect 127 194 128 195 
rect 127 200 128 201 
rect 127 219 128 220 
rect 127 228 128 229 
rect 127 232 128 233 
rect 127 238 128 239 
rect 127 241 128 242 
rect 127 243 128 244 
rect 127 254 128 255 
rect 127 257 128 258 
rect 127 261 128 262 
rect 127 273 128 274 
rect 127 280 128 281 
rect 127 289 128 290 
rect 127 291 128 292 
rect 127 305 128 306 
rect 127 308 128 309 
rect 127 310 128 311 
rect 127 312 128 313 
rect 128 1 129 2 
rect 128 3 129 4 
rect 128 8 129 9 
rect 128 14 129 15 
rect 128 17 129 18 
rect 128 20 129 21 
rect 128 23 129 24 
rect 128 48 129 49 
rect 128 49 129 50 
rect 128 72 129 73 
rect 128 73 129 74 
rect 128 113 129 114 
rect 128 128 129 129 
rect 128 129 129 130 
rect 128 132 129 133 
rect 128 136 129 137 
rect 128 139 129 140 
rect 128 152 129 153 
rect 128 161 129 162 
rect 128 164 129 165 
rect 128 183 129 184 
rect 128 194 129 195 
rect 128 200 129 201 
rect 128 201 129 202 
rect 128 219 129 220 
rect 128 228 129 229 
rect 128 232 129 233 
rect 128 238 129 239 
rect 128 241 129 242 
rect 128 243 129 244 
rect 128 254 129 255 
rect 128 272 129 273 
rect 128 273 129 274 
rect 128 280 129 281 
rect 128 289 129 290 
rect 128 291 129 292 
rect 128 305 129 306 
rect 128 308 129 309 
rect 128 310 129 311 
rect 128 312 129 313 
rect 129 1 130 2 
rect 129 3 130 4 
rect 129 8 130 9 
rect 129 14 130 15 
rect 129 15 130 16 
rect 129 17 130 18 
rect 129 20 130 21 
rect 129 23 130 24 
rect 129 26 130 27 
rect 129 27 130 28 
rect 129 113 130 114 
rect 129 116 130 117 
rect 129 117 130 118 
rect 129 118 130 119 
rect 129 119 130 120 
rect 129 120 130 121 
rect 129 121 130 122 
rect 129 122 130 123 
rect 129 123 130 124 
rect 129 124 130 125 
rect 129 125 130 126 
rect 129 126 130 127 
rect 129 127 130 128 
rect 129 128 130 129 
rect 129 132 130 133 
rect 129 136 130 137 
rect 129 138 130 139 
rect 129 139 130 140 
rect 129 152 130 153 
rect 129 161 130 162 
rect 129 164 130 165 
rect 129 183 130 184 
rect 129 194 130 195 
rect 129 201 130 202 
rect 129 202 130 203 
rect 129 203 130 204 
rect 129 204 130 205 
rect 129 205 130 206 
rect 129 206 130 207 
rect 129 219 130 220 
rect 129 228 130 229 
rect 129 232 130 233 
rect 129 238 130 239 
rect 129 239 130 240 
rect 129 241 130 242 
rect 129 243 130 244 
rect 129 248 130 249 
rect 129 249 130 250 
rect 129 250 130 251 
rect 129 251 130 252 
rect 129 252 130 253 
rect 129 253 130 254 
rect 129 254 130 255 
rect 129 256 130 257 
rect 129 257 130 258 
rect 129 258 130 259 
rect 129 259 130 260 
rect 129 260 130 261 
rect 129 261 130 262 
rect 129 262 130 263 
rect 129 263 130 264 
rect 129 264 130 265 
rect 129 265 130 266 
rect 129 266 130 267 
rect 129 267 130 268 
rect 129 268 130 269 
rect 129 269 130 270 
rect 129 270 130 271 
rect 129 271 130 272 
rect 129 272 130 273 
rect 129 280 130 281 
rect 129 289 130 290 
rect 129 291 130 292 
rect 129 305 130 306 
rect 129 308 130 309 
rect 129 310 130 311 
rect 129 312 130 313 
rect 130 1 131 2 
rect 130 3 131 4 
rect 130 8 131 9 
rect 130 17 131 18 
rect 130 20 131 21 
rect 130 23 131 24 
rect 130 27 131 28 
rect 130 28 131 29 
rect 130 29 131 30 
rect 130 30 131 31 
rect 130 31 131 32 
rect 130 32 131 33 
rect 130 33 131 34 
rect 130 34 131 35 
rect 130 35 131 36 
rect 130 36 131 37 
rect 130 37 131 38 
rect 130 38 131 39 
rect 130 39 131 40 
rect 130 40 131 41 
rect 130 41 131 42 
rect 130 42 131 43 
rect 130 43 131 44 
rect 130 44 131 45 
rect 130 45 131 46 
rect 130 46 131 47 
rect 130 47 131 48 
rect 130 48 131 49 
rect 130 49 131 50 
rect 130 50 131 51 
rect 130 51 131 52 
rect 130 52 131 53 
rect 130 53 131 54 
rect 130 54 131 55 
rect 130 55 131 56 
rect 130 56 131 57 
rect 130 57 131 58 
rect 130 58 131 59 
rect 130 59 131 60 
rect 130 60 131 61 
rect 130 61 131 62 
rect 130 62 131 63 
rect 130 63 131 64 
rect 130 64 131 65 
rect 130 65 131 66 
rect 130 66 131 67 
rect 130 67 131 68 
rect 130 68 131 69 
rect 130 69 131 70 
rect 130 70 131 71 
rect 130 71 131 72 
rect 130 72 131 73 
rect 130 73 131 74 
rect 130 74 131 75 
rect 130 75 131 76 
rect 130 76 131 77 
rect 130 77 131 78 
rect 130 78 131 79 
rect 130 79 131 80 
rect 130 80 131 81 
rect 130 81 131 82 
rect 130 82 131 83 
rect 130 83 131 84 
rect 130 84 131 85 
rect 130 85 131 86 
rect 130 86 131 87 
rect 130 87 131 88 
rect 130 88 131 89 
rect 130 89 131 90 
rect 130 90 131 91 
rect 130 91 131 92 
rect 130 92 131 93 
rect 130 93 131 94 
rect 130 94 131 95 
rect 130 95 131 96 
rect 130 96 131 97 
rect 130 97 131 98 
rect 130 98 131 99 
rect 130 99 131 100 
rect 130 100 131 101 
rect 130 101 131 102 
rect 130 102 131 103 
rect 130 103 131 104 
rect 130 104 131 105 
rect 130 105 131 106 
rect 130 106 131 107 
rect 130 107 131 108 
rect 130 108 131 109 
rect 130 109 131 110 
rect 130 110 131 111 
rect 130 111 131 112 
rect 130 113 131 114 
rect 130 116 131 117 
rect 130 132 131 133 
rect 130 136 131 137 
rect 130 138 131 139 
rect 130 141 131 142 
rect 130 152 131 153 
rect 130 161 131 162 
rect 130 164 131 165 
rect 130 183 131 184 
rect 130 194 131 195 
rect 130 206 131 207 
rect 130 219 131 220 
rect 130 228 131 229 
rect 130 232 131 233 
rect 130 241 131 242 
rect 130 243 131 244 
rect 130 248 131 249 
rect 130 255 131 256 
rect 130 256 131 257 
rect 130 280 131 281 
rect 130 289 131 290 
rect 130 291 131 292 
rect 130 305 131 306 
rect 130 308 131 309 
rect 130 310 131 311 
rect 130 312 131 313 
rect 131 1 132 2 
rect 131 3 132 4 
rect 131 8 132 9 
rect 131 17 132 18 
rect 131 20 132 21 
rect 131 23 132 24 
rect 131 113 132 114 
rect 131 116 132 117 
rect 131 132 132 133 
rect 131 136 132 137 
rect 131 138 132 139 
rect 131 141 132 142 
rect 131 142 132 143 
rect 131 143 132 144 
rect 131 144 132 145 
rect 131 145 132 146 
rect 131 146 132 147 
rect 131 147 132 148 
rect 131 148 132 149 
rect 131 152 132 153 
rect 131 161 132 162 
rect 131 164 132 165 
rect 131 183 132 184 
rect 131 194 132 195 
rect 131 206 132 207 
rect 131 219 132 220 
rect 131 221 132 222 
rect 131 222 132 223 
rect 131 223 132 224 
rect 131 224 132 225 
rect 131 225 132 226 
rect 131 226 132 227 
rect 131 227 132 228 
rect 131 228 132 229 
rect 131 232 132 233 
rect 131 241 132 242 
rect 131 243 132 244 
rect 131 248 132 249 
rect 131 250 132 251 
rect 131 251 132 252 
rect 131 252 132 253 
rect 131 253 132 254 
rect 131 254 132 255 
rect 131 255 132 256 
rect 131 280 132 281 
rect 131 289 132 290 
rect 131 291 132 292 
rect 131 305 132 306 
rect 131 308 132 309 
rect 131 310 132 311 
rect 131 312 132 313 
rect 132 1 133 2 
rect 132 3 133 4 
rect 132 8 133 9 
rect 132 17 133 18 
rect 132 20 133 21 
rect 132 23 133 24 
rect 132 36 133 37 
rect 132 37 133 38 
rect 132 38 133 39 
rect 132 39 133 40 
rect 132 40 133 41 
rect 132 41 133 42 
rect 132 42 133 43 
rect 132 43 133 44 
rect 132 44 133 45 
rect 132 45 133 46 
rect 132 46 133 47 
rect 132 47 133 48 
rect 132 87 133 88 
rect 132 88 133 89 
rect 132 89 133 90 
rect 132 90 133 91 
rect 132 91 133 92 
rect 132 92 133 93 
rect 132 93 133 94 
rect 132 94 133 95 
rect 132 95 133 96 
rect 132 98 133 99 
rect 132 99 133 100 
rect 132 100 133 101 
rect 132 113 133 114 
rect 132 116 133 117 
rect 132 132 133 133 
rect 132 136 133 137 
rect 132 138 133 139 
rect 132 152 133 153 
rect 132 161 133 162 
rect 132 164 133 165 
rect 132 183 133 184 
rect 132 194 133 195 
rect 132 206 133 207 
rect 132 219 133 220 
rect 132 221 133 222 
rect 132 232 133 233 
rect 132 241 133 242 
rect 132 243 133 244 
rect 132 248 133 249 
rect 132 250 133 251 
rect 132 280 133 281 
rect 132 289 133 290 
rect 132 291 133 292 
rect 132 305 133 306 
rect 132 308 133 309 
rect 132 310 133 311 
rect 132 312 133 313 
rect 133 1 134 2 
rect 133 3 134 4 
rect 133 8 134 9 
rect 133 17 134 18 
rect 133 20 134 21 
rect 133 23 134 24 
rect 133 36 134 37 
rect 133 95 134 96 
rect 133 96 134 97 
rect 133 100 134 101 
rect 133 113 134 114 
rect 133 132 134 133 
rect 133 136 134 137 
rect 133 152 134 153 
rect 133 161 134 162 
rect 133 164 134 165 
rect 133 183 134 184 
rect 133 194 134 195 
rect 133 206 134 207 
rect 133 219 134 220 
rect 133 232 134 233 
rect 133 241 134 242 
rect 133 243 134 244 
rect 133 248 134 249 
rect 133 253 134 254 
rect 133 254 134 255 
rect 133 255 134 256 
rect 133 256 134 257 
rect 133 257 134 258 
rect 133 258 134 259 
rect 133 259 134 260 
rect 133 280 134 281 
rect 133 289 134 290 
rect 133 291 134 292 
rect 133 305 134 306 
rect 133 308 134 309 
rect 133 310 134 311 
rect 133 312 134 313 
rect 134 1 135 2 
rect 134 3 135 4 
rect 134 8 135 9 
rect 134 17 135 18 
rect 134 20 135 21 
rect 134 23 135 24 
rect 134 36 135 37 
rect 134 70 135 71 
rect 134 71 135 72 
rect 134 72 135 73 
rect 134 73 135 74 
rect 134 74 135 75 
rect 134 75 135 76 
rect 134 76 135 77 
rect 134 77 135 78 
rect 134 78 135 79 
rect 134 79 135 80 
rect 134 80 135 81 
rect 134 81 135 82 
rect 134 82 135 83 
rect 134 83 135 84 
rect 134 84 135 85 
rect 134 96 135 97 
rect 134 97 135 98 
rect 134 100 135 101 
rect 134 101 135 102 
rect 134 102 135 103 
rect 134 103 135 104 
rect 134 104 135 105 
rect 134 105 135 106 
rect 134 106 135 107 
rect 134 107 135 108 
rect 134 108 135 109 
rect 134 109 135 110 
rect 134 110 135 111 
rect 134 111 135 112 
rect 134 113 135 114 
rect 134 114 135 115 
rect 134 115 135 116 
rect 134 116 135 117 
rect 134 117 135 118 
rect 134 132 135 133 
rect 134 136 135 137 
rect 134 152 135 153 
rect 134 161 135 162 
rect 134 164 135 165 
rect 134 183 135 184 
rect 134 194 135 195 
rect 134 195 135 196 
rect 134 206 135 207 
rect 134 207 135 208 
rect 134 208 135 209 
rect 134 209 135 210 
rect 134 210 135 211 
rect 134 211 135 212 
rect 134 219 135 220 
rect 134 220 135 221 
rect 134 221 135 222 
rect 134 222 135 223 
rect 134 223 135 224 
rect 134 224 135 225 
rect 134 225 135 226 
rect 134 226 135 227 
rect 134 227 135 228 
rect 134 228 135 229 
rect 134 229 135 230 
rect 134 232 135 233 
rect 134 241 135 242 
rect 134 243 135 244 
rect 134 244 135 245 
rect 134 245 135 246 
rect 134 246 135 247 
rect 134 248 135 249 
rect 134 259 135 260 
rect 134 280 135 281 
rect 134 289 135 290 
rect 134 291 135 292 
rect 134 305 135 306 
rect 134 308 135 309 
rect 134 310 135 311 
rect 134 312 135 313 
rect 135 1 136 2 
rect 135 3 136 4 
rect 135 8 136 9 
rect 135 17 136 18 
rect 135 20 136 21 
rect 135 23 136 24 
rect 135 36 136 37 
rect 135 289 136 290 
rect 135 291 136 292 
rect 135 305 136 306 
rect 135 308 136 309 
rect 135 310 136 311 
rect 135 312 136 313 
rect 136 1 137 2 
rect 136 3 137 4 
rect 136 8 137 9 
rect 136 17 137 18 
rect 136 20 137 21 
rect 136 23 137 24 
rect 136 34 137 35 
rect 136 35 137 36 
rect 136 36 137 37 
rect 136 41 137 42 
rect 136 42 137 43 
rect 136 43 137 44 
rect 136 44 137 45 
rect 136 45 137 46 
rect 136 46 137 47 
rect 136 47 137 48 
rect 136 48 137 49 
rect 136 49 137 50 
rect 136 50 137 51 
rect 136 51 137 52 
rect 136 52 137 53 
rect 136 53 137 54 
rect 136 54 137 55 
rect 136 55 137 56 
rect 136 56 137 57 
rect 136 57 137 58 
rect 136 58 137 59 
rect 136 59 137 60 
rect 136 60 137 61 
rect 136 61 137 62 
rect 136 62 137 63 
rect 136 63 137 64 
rect 136 64 137 65 
rect 136 65 137 66 
rect 136 66 137 67 
rect 136 67 137 68 
rect 136 68 137 69 
rect 136 69 137 70 
rect 136 70 137 71 
rect 136 71 137 72 
rect 136 72 137 73 
rect 136 73 137 74 
rect 136 74 137 75 
rect 136 75 137 76 
rect 136 76 137 77 
rect 136 77 137 78 
rect 136 78 137 79 
rect 136 79 137 80 
rect 136 80 137 81 
rect 136 81 137 82 
rect 136 82 137 83 
rect 136 83 137 84 
rect 136 84 137 85 
rect 136 85 137 86 
rect 136 86 137 87 
rect 136 87 137 88 
rect 136 88 137 89 
rect 136 89 137 90 
rect 136 90 137 91 
rect 136 91 137 92 
rect 136 92 137 93 
rect 136 93 137 94 
rect 136 94 137 95 
rect 136 95 137 96 
rect 136 96 137 97 
rect 136 97 137 98 
rect 136 98 137 99 
rect 136 99 137 100 
rect 136 100 137 101 
rect 136 101 137 102 
rect 136 102 137 103 
rect 136 103 137 104 
rect 136 104 137 105 
rect 136 105 137 106 
rect 136 106 137 107 
rect 136 107 137 108 
rect 136 110 137 111 
rect 136 111 137 112 
rect 136 112 137 113 
rect 136 113 137 114 
rect 136 114 137 115 
rect 136 115 137 116 
rect 136 116 137 117 
rect 136 117 137 118 
rect 136 118 137 119 
rect 136 119 137 120 
rect 136 120 137 121 
rect 136 121 137 122 
rect 136 122 137 123 
rect 136 123 137 124 
rect 136 124 137 125 
rect 136 125 137 126 
rect 136 126 137 127 
rect 136 127 137 128 
rect 136 128 137 129 
rect 136 129 137 130 
rect 136 130 137 131 
rect 136 131 137 132 
rect 136 132 137 133 
rect 136 133 137 134 
rect 136 134 137 135 
rect 136 135 137 136 
rect 136 136 137 137 
rect 136 137 137 138 
rect 136 138 137 139 
rect 136 139 137 140 
rect 136 140 137 141 
rect 136 141 137 142 
rect 136 142 137 143 
rect 136 143 137 144 
rect 136 144 137 145 
rect 136 145 137 146 
rect 136 146 137 147 
rect 136 147 137 148 
rect 136 148 137 149 
rect 136 149 137 150 
rect 136 150 137 151 
rect 136 151 137 152 
rect 136 152 137 153 
rect 136 153 137 154 
rect 136 154 137 155 
rect 136 155 137 156 
rect 136 156 137 157 
rect 136 157 137 158 
rect 136 158 137 159 
rect 136 159 137 160 
rect 136 160 137 161 
rect 136 161 137 162 
rect 136 162 137 163 
rect 136 163 137 164 
rect 136 164 137 165 
rect 136 165 137 166 
rect 136 166 137 167 
rect 136 167 137 168 
rect 136 168 137 169 
rect 136 169 137 170 
rect 136 170 137 171 
rect 136 171 137 172 
rect 136 172 137 173 
rect 136 173 137 174 
rect 136 174 137 175 
rect 136 175 137 176 
rect 136 176 137 177 
rect 136 177 137 178 
rect 136 178 137 179 
rect 136 179 137 180 
rect 136 180 137 181 
rect 136 181 137 182 
rect 136 182 137 183 
rect 136 183 137 184 
rect 136 184 137 185 
rect 136 185 137 186 
rect 136 186 137 187 
rect 136 187 137 188 
rect 136 188 137 189 
rect 136 189 137 190 
rect 136 190 137 191 
rect 136 191 137 192 
rect 136 192 137 193 
rect 136 193 137 194 
rect 136 194 137 195 
rect 136 195 137 196 
rect 136 196 137 197 
rect 136 197 137 198 
rect 136 198 137 199 
rect 136 199 137 200 
rect 136 200 137 201 
rect 136 201 137 202 
rect 136 202 137 203 
rect 136 203 137 204 
rect 136 204 137 205 
rect 136 205 137 206 
rect 136 206 137 207 
rect 136 207 137 208 
rect 136 208 137 209 
rect 136 209 137 210 
rect 136 210 137 211 
rect 136 211 137 212 
rect 136 212 137 213 
rect 136 213 137 214 
rect 136 214 137 215 
rect 136 215 137 216 
rect 136 216 137 217 
rect 136 217 137 218 
rect 136 218 137 219 
rect 136 219 137 220 
rect 136 220 137 221 
rect 136 221 137 222 
rect 136 222 137 223 
rect 136 223 137 224 
rect 136 224 137 225 
rect 136 225 137 226 
rect 136 226 137 227 
rect 136 227 137 228 
rect 136 228 137 229 
rect 136 229 137 230 
rect 136 230 137 231 
rect 136 231 137 232 
rect 136 232 137 233 
rect 136 233 137 234 
rect 136 234 137 235 
rect 136 235 137 236 
rect 136 236 137 237 
rect 136 237 137 238 
rect 136 238 137 239 
rect 136 239 137 240 
rect 136 240 137 241 
rect 136 241 137 242 
rect 136 242 137 243 
rect 136 243 137 244 
rect 136 244 137 245 
rect 136 245 137 246 
rect 136 246 137 247 
rect 136 247 137 248 
rect 136 248 137 249 
rect 136 249 137 250 
rect 136 250 137 251 
rect 136 251 137 252 
rect 136 252 137 253 
rect 136 253 137 254 
rect 136 254 137 255 
rect 136 255 137 256 
rect 136 256 137 257 
rect 136 257 137 258 
rect 136 258 137 259 
rect 136 259 137 260 
rect 136 260 137 261 
rect 136 261 137 262 
rect 136 262 137 263 
rect 136 263 137 264 
rect 136 264 137 265 
rect 136 265 137 266 
rect 136 266 137 267 
rect 136 267 137 268 
rect 136 268 137 269 
rect 136 269 137 270 
rect 136 270 137 271 
rect 136 271 137 272 
rect 136 272 137 273 
rect 136 273 137 274 
rect 136 274 137 275 
rect 136 275 137 276 
rect 136 276 137 277 
rect 136 277 137 278 
rect 136 278 137 279 
rect 136 279 137 280 
rect 136 280 137 281 
rect 136 281 137 282 
rect 136 282 137 283 
rect 136 283 137 284 
rect 136 284 137 285 
rect 136 285 137 286 
rect 136 286 137 287 
rect 136 287 137 288 
rect 136 288 137 289 
rect 136 291 137 292 
rect 136 305 137 306 
rect 136 308 137 309 
rect 136 310 137 311 
rect 136 312 137 313 
rect 137 1 138 2 
rect 137 3 138 4 
rect 137 8 138 9 
rect 137 17 138 18 
rect 137 20 138 21 
rect 137 23 138 24 
rect 137 34 138 35 
rect 137 40 138 41 
rect 137 41 138 42 
rect 137 107 138 108 
rect 137 110 138 111 
rect 137 288 138 289 
rect 137 289 138 290 
rect 137 305 138 306 
rect 137 308 138 309 
rect 137 310 138 311 
rect 137 312 138 313 
rect 138 1 139 2 
rect 138 3 139 4 
rect 138 8 139 9 
rect 138 17 139 18 
rect 138 20 139 21 
rect 138 23 139 24 
rect 138 34 139 35 
rect 138 36 139 37 
rect 138 37 139 38 
rect 138 38 139 39 
rect 138 39 139 40 
rect 138 40 139 41 
rect 138 107 139 108 
rect 138 110 139 111 
rect 138 114 139 115 
rect 138 115 139 116 
rect 138 118 139 119 
rect 138 133 139 134 
rect 138 162 139 163 
rect 138 163 139 164 
rect 138 164 139 165 
rect 138 165 139 166 
rect 138 166 139 167 
rect 138 167 139 168 
rect 138 168 139 169 
rect 138 225 139 226 
rect 138 226 139 227 
rect 138 227 139 228 
rect 138 228 139 229 
rect 138 229 139 230 
rect 138 230 139 231 
rect 138 231 139 232 
rect 138 241 139 242 
rect 138 242 139 243 
rect 138 243 139 244 
rect 138 244 139 245 
rect 138 245 139 246 
rect 138 246 139 247 
rect 138 247 139 248 
rect 138 260 139 261 
rect 138 261 139 262 
rect 138 262 139 263 
rect 138 273 139 274 
rect 138 274 139 275 
rect 138 275 139 276 
rect 138 276 139 277 
rect 138 277 139 278 
rect 138 278 139 279 
rect 138 279 139 280 
rect 138 289 139 290 
rect 138 290 139 291 
rect 138 291 139 292 
rect 138 292 139 293 
rect 138 293 139 294 
rect 138 305 139 306 
rect 138 308 139 309 
rect 138 310 139 311 
rect 138 312 139 313 
rect 139 1 140 2 
rect 139 3 140 4 
rect 139 8 140 9 
rect 139 17 140 18 
rect 139 20 140 21 
rect 139 23 140 24 
rect 139 34 140 35 
rect 139 36 140 37 
rect 139 114 140 115 
rect 139 118 140 119 
rect 139 133 140 134 
rect 139 136 140 137 
rect 139 145 140 146 
rect 139 148 140 149 
rect 139 168 140 169 
rect 139 225 140 226 
rect 139 241 140 242 
rect 139 262 140 263 
rect 139 273 140 274 
rect 139 293 140 294 
rect 139 305 140 306 
rect 139 308 140 309 
rect 139 310 140 311 
rect 139 312 140 313 
rect 140 1 141 2 
rect 140 3 141 4 
rect 140 8 141 9 
rect 140 17 141 18 
rect 140 20 141 21 
rect 140 23 141 24 
rect 140 34 141 35 
rect 140 36 141 37 
rect 140 114 141 115 
rect 140 118 141 119 
rect 140 133 141 134 
rect 140 136 141 137 
rect 140 145 141 146 
rect 140 148 141 149 
rect 140 168 141 169 
rect 140 225 141 226 
rect 140 230 141 231 
rect 140 241 141 242 
rect 140 244 141 245 
rect 140 245 141 246 
rect 140 246 141 247 
rect 140 247 141 248 
rect 140 248 141 249 
rect 140 262 141 263 
rect 140 263 141 264 
rect 140 273 141 274 
rect 140 276 141 277 
rect 140 277 141 278 
rect 140 293 141 294 
rect 140 305 141 306 
rect 140 308 141 309 
rect 140 310 141 311 
rect 140 312 141 313 
rect 141 1 142 2 
rect 141 3 142 4 
rect 141 8 142 9 
rect 141 17 142 18 
rect 141 20 142 21 
rect 141 23 142 24 
rect 141 34 142 35 
rect 141 36 142 37 
rect 141 114 142 115 
rect 141 118 142 119 
rect 141 133 142 134 
rect 141 136 142 137 
rect 141 145 142 146 
rect 141 148 142 149 
rect 141 163 142 164 
rect 141 168 142 169 
rect 141 225 142 226 
rect 141 228 142 229 
rect 141 230 142 231 
rect 141 241 142 242 
rect 141 248 142 249 
rect 141 263 142 264 
rect 141 273 142 274 
rect 141 276 142 277 
rect 141 289 142 290 
rect 141 291 142 292 
rect 141 293 142 294 
rect 141 305 142 306 
rect 141 308 142 309 
rect 141 310 142 311 
rect 141 312 142 313 
rect 142 1 143 2 
rect 142 3 143 4 
rect 142 8 143 9 
rect 142 17 143 18 
rect 142 20 143 21 
rect 142 23 143 24 
rect 142 34 143 35 
rect 142 36 143 37 
rect 142 114 143 115 
rect 142 118 143 119 
rect 142 133 143 134 
rect 142 136 143 137 
rect 142 145 143 146 
rect 142 148 143 149 
rect 142 161 143 162 
rect 142 163 143 164 
rect 142 168 143 169 
rect 142 225 143 226 
rect 142 228 143 229 
rect 142 230 143 231 
rect 142 241 143 242 
rect 142 248 143 249 
rect 142 263 143 264 
rect 142 273 143 274 
rect 142 276 143 277 
rect 142 279 143 280 
rect 142 280 143 281 
rect 142 289 143 290 
rect 142 291 143 292 
rect 142 293 143 294 
rect 142 305 143 306 
rect 142 308 143 309 
rect 142 310 143 311 
rect 142 312 143 313 
rect 143 1 144 2 
rect 143 3 144 4 
rect 143 8 144 9 
rect 143 14 144 15 
rect 143 17 144 18 
rect 143 20 144 21 
rect 143 23 144 24 
rect 143 27 144 28 
rect 143 34 144 35 
rect 143 36 144 37 
rect 143 107 144 108 
rect 143 114 144 115 
rect 143 118 144 119 
rect 143 133 144 134 
rect 143 136 144 137 
rect 143 139 144 140 
rect 143 145 144 146 
rect 143 148 144 149 
rect 143 161 144 162 
rect 143 163 144 164 
rect 143 165 144 166 
rect 143 166 144 167 
rect 143 168 144 169 
rect 143 225 144 226 
rect 143 228 144 229 
rect 143 230 144 231 
rect 143 241 144 242 
rect 143 248 144 249 
rect 143 251 144 252 
rect 143 263 144 264 
rect 143 273 144 274 
rect 143 276 144 277 
rect 143 280 144 281 
rect 143 289 144 290 
rect 143 291 144 292 
rect 143 293 144 294 
rect 143 302 144 303 
rect 143 305 144 306 
rect 143 308 144 309 
rect 143 310 144 311 
rect 143 312 144 313 
rect 144 1 145 2 
rect 144 3 145 4 
rect 144 8 145 9 
rect 144 14 145 15 
rect 144 16 145 17 
rect 144 17 145 18 
rect 144 20 145 21 
rect 144 23 145 24 
rect 144 27 145 28 
rect 144 34 145 35 
rect 144 36 145 37 
rect 144 107 145 108 
rect 144 114 145 115 
rect 144 118 145 119 
rect 144 133 145 134 
rect 144 136 145 137 
rect 144 139 145 140 
rect 144 144 145 145 
rect 144 145 145 146 
rect 144 148 145 149 
rect 144 161 145 162 
rect 144 163 145 164 
rect 144 165 145 166 
rect 144 168 145 169 
rect 144 169 145 170 
rect 144 177 145 178 
rect 144 178 145 179 
rect 144 179 145 180 
rect 144 180 145 181 
rect 144 181 145 182 
rect 144 182 145 183 
rect 144 183 145 184 
rect 144 184 145 185 
rect 144 185 145 186 
rect 144 224 145 225 
rect 144 225 145 226 
rect 144 227 145 228 
rect 144 228 145 229 
rect 144 230 145 231 
rect 144 240 145 241 
rect 144 241 145 242 
rect 144 248 145 249 
rect 144 251 145 252 
rect 144 263 145 264 
rect 144 273 145 274 
rect 144 276 145 277 
rect 144 280 145 281 
rect 144 281 145 282 
rect 144 288 145 289 
rect 144 289 145 290 
rect 144 291 145 292 
rect 144 293 145 294 
rect 144 302 145 303 
rect 144 305 145 306 
rect 144 308 145 309 
rect 144 310 145 311 
rect 144 312 145 313 
rect 145 1 146 2 
rect 145 3 146 4 
rect 145 8 146 9 
rect 145 14 146 15 
rect 145 15 146 16 
rect 145 16 146 17 
rect 145 20 146 21 
rect 145 23 146 24 
rect 145 27 146 28 
rect 145 34 146 35 
rect 145 36 146 37 
rect 145 38 146 39 
rect 145 39 146 40 
rect 145 40 146 41 
rect 145 41 146 42 
rect 145 42 146 43 
rect 145 43 146 44 
rect 145 44 146 45 
rect 145 45 146 46 
rect 145 46 146 47 
rect 145 47 146 48 
rect 145 48 146 49 
rect 145 49 146 50 
rect 145 50 146 51 
rect 145 51 146 52 
rect 145 52 146 53 
rect 145 53 146 54 
rect 145 54 146 55 
rect 145 55 146 56 
rect 145 56 146 57 
rect 145 57 146 58 
rect 145 58 146 59 
rect 145 59 146 60 
rect 145 60 146 61 
rect 145 61 146 62 
rect 145 62 146 63 
rect 145 63 146 64 
rect 145 64 146 65 
rect 145 65 146 66 
rect 145 66 146 67 
rect 145 67 146 68 
rect 145 68 146 69 
rect 145 69 146 70 
rect 145 70 146 71 
rect 145 71 146 72 
rect 145 72 146 73 
rect 145 73 146 74 
rect 145 74 146 75 
rect 145 75 146 76 
rect 145 76 146 77 
rect 145 77 146 78 
rect 145 78 146 79 
rect 145 79 146 80 
rect 145 80 146 81 
rect 145 81 146 82 
rect 145 82 146 83 
rect 145 83 146 84 
rect 145 84 146 85 
rect 145 85 146 86 
rect 145 86 146 87 
rect 145 87 146 88 
rect 145 88 146 89 
rect 145 89 146 90 
rect 145 90 146 91 
rect 145 91 146 92 
rect 145 92 146 93 
rect 145 93 146 94 
rect 145 94 146 95 
rect 145 95 146 96 
rect 145 96 146 97 
rect 145 97 146 98 
rect 145 98 146 99 
rect 145 99 146 100 
rect 145 100 146 101 
rect 145 101 146 102 
rect 145 102 146 103 
rect 145 103 146 104 
rect 145 104 146 105 
rect 145 105 146 106 
rect 145 106 146 107 
rect 145 107 146 108 
rect 145 114 146 115 
rect 145 118 146 119 
rect 145 133 146 134 
rect 145 136 146 137 
rect 145 139 146 140 
rect 145 140 146 141 
rect 145 141 146 142 
rect 145 142 146 143 
rect 145 143 146 144 
rect 145 144 146 145 
rect 145 148 146 149 
rect 145 149 146 150 
rect 145 150 146 151 
rect 145 151 146 152 
rect 145 152 146 153 
rect 145 153 146 154 
rect 145 154 146 155 
rect 145 155 146 156 
rect 145 156 146 157 
rect 145 157 146 158 
rect 145 161 146 162 
rect 145 163 146 164 
rect 145 165 146 166 
rect 145 169 146 170 
rect 145 172 146 173 
rect 145 173 146 174 
rect 145 174 146 175 
rect 145 175 146 176 
rect 145 176 146 177 
rect 145 177 146 178 
rect 145 185 146 186 
rect 145 186 146 187 
rect 145 187 146 188 
rect 145 188 146 189 
rect 145 189 146 190 
rect 145 190 146 191 
rect 145 191 146 192 
rect 145 192 146 193 
rect 145 193 146 194 
rect 145 194 146 195 
rect 145 195 146 196 
rect 145 196 146 197 
rect 145 197 146 198 
rect 145 198 146 199 
rect 145 199 146 200 
rect 145 200 146 201 
rect 145 201 146 202 
rect 145 202 146 203 
rect 145 203 146 204 
rect 145 204 146 205 
rect 145 205 146 206 
rect 145 206 146 207 
rect 145 207 146 208 
rect 145 208 146 209 
rect 145 209 146 210 
rect 145 210 146 211 
rect 145 211 146 212 
rect 145 212 146 213 
rect 145 213 146 214 
rect 145 214 146 215 
rect 145 215 146 216 
rect 145 216 146 217 
rect 145 217 146 218 
rect 145 218 146 219 
rect 145 219 146 220 
rect 145 220 146 221 
rect 145 221 146 222 
rect 145 222 146 223 
rect 145 224 146 225 
rect 145 226 146 227 
rect 145 227 146 228 
rect 145 230 146 231 
rect 145 240 146 241 
rect 145 248 146 249 
rect 145 251 146 252 
rect 145 252 146 253 
rect 145 253 146 254 
rect 145 254 146 255 
rect 145 255 146 256 
rect 145 256 146 257 
rect 145 257 146 258 
rect 145 258 146 259 
rect 145 259 146 260 
rect 145 263 146 264 
rect 145 273 146 274 
rect 145 276 146 277 
rect 145 281 146 282 
rect 145 282 146 283 
rect 145 283 146 284 
rect 145 284 146 285 
rect 145 285 146 286 
rect 145 286 146 287 
rect 145 288 146 289 
rect 145 290 146 291 
rect 145 291 146 292 
rect 145 293 146 294 
rect 145 296 146 297 
rect 145 297 146 298 
rect 145 298 146 299 
rect 145 299 146 300 
rect 145 300 146 301 
rect 145 301 146 302 
rect 145 302 146 303 
rect 145 305 146 306 
rect 145 308 146 309 
rect 145 310 146 311 
rect 145 312 146 313 
rect 146 1 147 2 
rect 146 3 147 4 
rect 146 8 147 9 
rect 146 18 147 19 
rect 146 20 147 21 
rect 146 23 147 24 
rect 146 27 147 28 
rect 146 34 147 35 
rect 146 36 147 37 
rect 146 38 147 39 
rect 146 114 147 115 
rect 146 118 147 119 
rect 146 133 147 134 
rect 146 136 147 137 
rect 146 157 147 158 
rect 146 160 147 161 
rect 146 161 147 162 
rect 146 163 147 164 
rect 146 165 147 166 
rect 146 169 147 170 
rect 146 181 147 182 
rect 146 182 147 183 
rect 146 183 147 184 
rect 146 224 147 225 
rect 146 226 147 227 
rect 146 230 147 231 
rect 146 231 147 232 
rect 146 232 147 233 
rect 146 233 147 234 
rect 146 234 147 235 
rect 146 235 147 236 
rect 146 236 147 237 
rect 146 237 147 238 
rect 146 238 147 239 
rect 146 240 147 241 
rect 146 242 147 243 
rect 146 248 147 249 
rect 146 259 147 260 
rect 146 263 147 264 
rect 146 273 147 274 
rect 146 276 147 277 
rect 146 288 147 289 
rect 146 290 147 291 
rect 146 293 147 294 
rect 146 305 147 306 
rect 146 308 147 309 
rect 146 310 147 311 
rect 146 312 147 313 
rect 147 1 148 2 
rect 147 3 148 4 
rect 147 8 148 9 
rect 147 18 148 19 
rect 147 20 148 21 
rect 147 23 148 24 
rect 147 27 148 28 
rect 147 34 148 35 
rect 147 36 148 37 
rect 147 38 148 39 
rect 147 48 148 49 
rect 147 49 148 50 
rect 147 50 148 51 
rect 147 51 148 52 
rect 147 52 148 53 
rect 147 53 148 54 
rect 147 54 148 55 
rect 147 55 148 56 
rect 147 58 148 59 
rect 147 59 148 60 
rect 147 60 148 61 
rect 147 61 148 62 
rect 147 62 148 63 
rect 147 63 148 64 
rect 147 64 148 65 
rect 147 65 148 66 
rect 147 66 148 67 
rect 147 67 148 68 
rect 147 68 148 69 
rect 147 69 148 70 
rect 147 70 148 71 
rect 147 71 148 72 
rect 147 72 148 73 
rect 147 73 148 74 
rect 147 74 148 75 
rect 147 75 148 76 
rect 147 76 148 77 
rect 147 77 148 78 
rect 147 78 148 79 
rect 147 79 148 80 
rect 147 80 148 81 
rect 147 81 148 82 
rect 147 82 148 83 
rect 147 83 148 84 
rect 147 84 148 85 
rect 147 85 148 86 
rect 147 86 148 87 
rect 147 87 148 88 
rect 147 88 148 89 
rect 147 89 148 90 
rect 147 90 148 91 
rect 147 91 148 92 
rect 147 92 148 93 
rect 147 93 148 94 
rect 147 94 148 95 
rect 147 95 148 96 
rect 147 96 148 97 
rect 147 97 148 98 
rect 147 98 148 99 
rect 147 99 148 100 
rect 147 100 148 101 
rect 147 101 148 102 
rect 147 102 148 103 
rect 147 103 148 104 
rect 147 114 148 115 
rect 147 118 148 119 
rect 147 133 148 134 
rect 147 136 148 137 
rect 147 157 148 158 
rect 147 159 148 160 
rect 147 160 148 161 
rect 147 163 148 164 
rect 147 169 148 170 
rect 147 171 148 172 
rect 147 172 148 173 
rect 147 173 148 174 
rect 147 174 148 175 
rect 147 175 148 176 
rect 147 176 148 177 
rect 147 177 148 178 
rect 147 178 148 179 
rect 147 179 148 180 
rect 147 180 148 181 
rect 147 181 148 182 
rect 147 210 148 211 
rect 147 224 148 225 
rect 147 226 148 227 
rect 147 240 148 241 
rect 147 242 148 243 
rect 147 244 148 245 
rect 147 245 148 246 
rect 147 273 148 274 
rect 147 276 148 277 
rect 147 288 148 289 
rect 147 290 148 291 
rect 147 293 148 294 
rect 147 305 148 306 
rect 147 308 148 309 
rect 147 310 148 311 
rect 147 312 148 313 
rect 148 1 149 2 
rect 148 3 149 4 
rect 148 8 149 9 
rect 148 18 149 19 
rect 148 20 149 21 
rect 148 23 149 24 
rect 148 27 149 28 
rect 148 34 149 35 
rect 148 36 149 37 
rect 148 38 149 39 
rect 148 48 149 49 
rect 148 57 149 58 
rect 148 58 149 59 
rect 148 114 149 115 
rect 148 118 149 119 
rect 148 133 149 134 
rect 148 136 149 137 
rect 148 159 149 160 
rect 148 161 149 162 
rect 148 162 149 163 
rect 148 163 149 164 
rect 148 166 149 167 
rect 148 167 149 168 
rect 148 169 149 170 
rect 148 171 149 172 
rect 148 187 149 188 
rect 148 188 149 189 
rect 148 189 149 190 
rect 148 190 149 191 
rect 148 191 149 192 
rect 148 192 149 193 
rect 148 193 149 194 
rect 148 194 149 195 
rect 148 195 149 196 
rect 148 196 149 197 
rect 148 197 149 198 
rect 148 198 149 199 
rect 148 199 149 200 
rect 148 200 149 201 
rect 148 201 149 202 
rect 148 202 149 203 
rect 148 203 149 204 
rect 148 204 149 205 
rect 148 205 149 206 
rect 148 206 149 207 
rect 148 207 149 208 
rect 148 208 149 209 
rect 148 209 149 210 
rect 148 210 149 211 
rect 148 224 149 225 
rect 148 226 149 227 
rect 148 240 149 241 
rect 148 242 149 243 
rect 148 243 149 244 
rect 148 245 149 246 
rect 148 246 149 247 
rect 148 247 149 248 
rect 148 248 149 249 
rect 148 249 149 250 
rect 148 250 149 251 
rect 148 251 149 252 
rect 148 252 149 253 
rect 148 253 149 254 
rect 148 254 149 255 
rect 148 255 149 256 
rect 148 256 149 257 
rect 148 257 149 258 
rect 148 258 149 259 
rect 148 259 149 260 
rect 148 260 149 261 
rect 148 261 149 262 
rect 148 262 149 263 
rect 148 263 149 264 
rect 148 264 149 265 
rect 148 265 149 266 
rect 148 266 149 267 
rect 148 267 149 268 
rect 148 268 149 269 
rect 148 269 149 270 
rect 148 270 149 271 
rect 148 271 149 272 
rect 148 273 149 274 
rect 148 276 149 277 
rect 148 288 149 289 
rect 148 290 149 291 
rect 148 293 149 294 
rect 148 305 149 306 
rect 148 308 149 309 
rect 148 310 149 311 
rect 148 312 149 313 
rect 149 1 150 2 
rect 149 3 150 4 
rect 149 8 150 9 
rect 149 18 150 19 
rect 149 20 150 21 
rect 149 23 150 24 
rect 149 27 150 28 
rect 149 34 150 35 
rect 149 36 150 37 
rect 149 38 150 39 
rect 149 48 150 49 
rect 149 114 150 115 
rect 149 118 150 119 
rect 149 133 150 134 
rect 149 136 150 137 
rect 149 159 150 160 
rect 149 161 150 162 
rect 149 166 150 167 
rect 149 169 150 170 
rect 149 171 150 172 
rect 149 187 150 188 
rect 149 224 150 225 
rect 149 226 150 227 
rect 149 240 150 241 
rect 149 243 150 244 
rect 149 271 150 272 
rect 149 273 150 274 
rect 149 276 150 277 
rect 149 288 150 289 
rect 149 290 150 291 
rect 149 293 150 294 
rect 149 305 150 306 
rect 149 308 150 309 
rect 149 310 150 311 
rect 149 312 150 313 
rect 150 1 151 2 
rect 150 3 151 4 
rect 150 8 151 9 
rect 150 18 151 19 
rect 150 20 151 21 
rect 150 23 151 24 
rect 150 27 151 28 
rect 150 34 151 35 
rect 150 36 151 37 
rect 150 38 151 39 
rect 150 48 151 49 
rect 150 114 151 115 
rect 150 118 151 119 
rect 150 133 151 134 
rect 150 136 151 137 
rect 150 152 151 153 
rect 150 153 151 154 
rect 150 154 151 155 
rect 150 155 151 156 
rect 150 156 151 157 
rect 150 157 151 158 
rect 150 159 151 160 
rect 150 161 151 162 
rect 150 166 151 167 
rect 150 169 151 170 
rect 150 187 151 188 
rect 150 189 151 190 
rect 150 190 151 191 
rect 150 191 151 192 
rect 150 192 151 193 
rect 150 193 151 194 
rect 150 194 151 195 
rect 150 195 151 196 
rect 150 196 151 197 
rect 150 224 151 225 
rect 150 226 151 227 
rect 150 240 151 241 
rect 150 243 151 244 
rect 150 271 151 272 
rect 150 273 151 274 
rect 150 276 151 277 
rect 150 288 151 289 
rect 150 290 151 291 
rect 150 293 151 294 
rect 150 305 151 306 
rect 150 308 151 309 
rect 150 310 151 311 
rect 150 312 151 313 
rect 151 1 152 2 
rect 151 3 152 4 
rect 151 8 152 9 
rect 151 18 152 19 
rect 151 20 152 21 
rect 151 23 152 24 
rect 151 27 152 28 
rect 151 34 152 35 
rect 151 36 152 37 
rect 151 38 152 39 
rect 151 48 152 49 
rect 151 114 152 115 
rect 151 118 152 119 
rect 151 133 152 134 
rect 151 136 152 137 
rect 151 151 152 152 
rect 151 152 152 153 
rect 151 159 152 160 
rect 151 161 152 162 
rect 151 166 152 167 
rect 151 169 152 170 
rect 151 187 152 188 
rect 151 224 152 225 
rect 151 226 152 227 
rect 151 240 152 241 
rect 151 243 152 244 
rect 151 271 152 272 
rect 151 273 152 274 
rect 151 276 152 277 
rect 151 288 152 289 
rect 151 290 152 291 
rect 151 293 152 294 
rect 151 305 152 306 
rect 151 308 152 309 
rect 151 310 152 311 
rect 151 312 152 313 
rect 152 1 153 2 
rect 152 3 153 4 
rect 152 8 153 9 
rect 152 18 153 19 
rect 152 20 153 21 
rect 152 23 153 24 
rect 152 25 153 26 
rect 152 26 153 27 
rect 152 27 153 28 
rect 152 33 153 34 
rect 152 34 153 35 
rect 152 36 153 37 
rect 152 38 153 39 
rect 152 40 153 41 
rect 152 41 153 42 
rect 152 42 153 43 
rect 152 43 153 44 
rect 152 44 153 45 
rect 152 45 153 46 
rect 152 46 153 47 
rect 152 47 153 48 
rect 152 48 153 49 
rect 152 50 153 51 
rect 152 51 153 52 
rect 152 52 153 53 
rect 152 53 153 54 
rect 152 54 153 55 
rect 152 55 153 56 
rect 152 56 153 57 
rect 152 57 153 58 
rect 152 58 153 59 
rect 152 59 153 60 
rect 152 60 153 61 
rect 152 61 153 62 
rect 152 62 153 63 
rect 152 63 153 64 
rect 152 64 153 65 
rect 152 65 153 66 
rect 152 66 153 67 
rect 152 67 153 68 
rect 152 68 153 69 
rect 152 69 153 70 
rect 152 70 153 71 
rect 152 71 153 72 
rect 152 72 153 73 
rect 152 73 153 74 
rect 152 74 153 75 
rect 152 75 153 76 
rect 152 76 153 77 
rect 152 77 153 78 
rect 152 78 153 79 
rect 152 79 153 80 
rect 152 80 153 81 
rect 152 81 153 82 
rect 152 82 153 83 
rect 152 83 153 84 
rect 152 84 153 85 
rect 152 85 153 86 
rect 152 86 153 87 
rect 152 87 153 88 
rect 152 88 153 89 
rect 152 89 153 90 
rect 152 90 153 91 
rect 152 91 153 92 
rect 152 92 153 93 
rect 152 93 153 94 
rect 152 94 153 95 
rect 152 95 153 96 
rect 152 96 153 97 
rect 152 97 153 98 
rect 152 98 153 99 
rect 152 99 153 100 
rect 152 100 153 101 
rect 152 101 153 102 
rect 152 102 153 103 
rect 152 103 153 104 
rect 152 104 153 105 
rect 152 105 153 106 
rect 152 106 153 107 
rect 152 107 153 108 
rect 152 108 153 109 
rect 152 109 153 110 
rect 152 110 153 111 
rect 152 111 153 112 
rect 152 112 153 113 
rect 152 113 153 114 
rect 152 114 153 115 
rect 152 118 153 119 
rect 152 129 153 130 
rect 152 130 153 131 
rect 152 131 153 132 
rect 152 132 153 133 
rect 152 133 153 134 
rect 152 136 153 137 
rect 152 145 153 146 
rect 152 146 153 147 
rect 152 147 153 148 
rect 152 148 153 149 
rect 152 149 153 150 
rect 152 150 153 151 
rect 152 151 153 152 
rect 152 153 153 154 
rect 152 154 153 155 
rect 152 155 153 156 
rect 152 156 153 157 
rect 152 157 153 158 
rect 152 158 153 159 
rect 152 159 153 160 
rect 152 161 153 162 
rect 152 165 153 166 
rect 152 166 153 167 
rect 152 169 153 170 
rect 152 170 153 171 
rect 152 171 153 172 
rect 152 172 153 173 
rect 152 173 153 174 
rect 152 174 153 175 
rect 152 175 153 176 
rect 152 176 153 177 
rect 152 177 153 178 
rect 152 178 153 179 
rect 152 179 153 180 
rect 152 180 153 181 
rect 152 181 153 182 
rect 152 182 153 183 
rect 152 183 153 184 
rect 152 184 153 185 
rect 152 187 153 188 
rect 152 193 153 194 
rect 152 194 153 195 
rect 152 195 153 196 
rect 152 196 153 197 
rect 152 197 153 198 
rect 152 198 153 199 
rect 152 199 153 200 
rect 152 200 153 201 
rect 152 201 153 202 
rect 152 202 153 203 
rect 152 203 153 204 
rect 152 204 153 205 
rect 152 205 153 206 
rect 152 206 153 207 
rect 152 207 153 208 
rect 152 208 153 209 
rect 152 209 153 210 
rect 152 210 153 211 
rect 152 211 153 212 
rect 152 212 153 213 
rect 152 213 153 214 
rect 152 214 153 215 
rect 152 215 153 216 
rect 152 216 153 217 
rect 152 217 153 218 
rect 152 218 153 219 
rect 152 219 153 220 
rect 152 220 153 221 
rect 152 221 153 222 
rect 152 222 153 223 
rect 152 223 153 224 
rect 152 224 153 225 
rect 152 226 153 227 
rect 152 233 153 234 
rect 152 234 153 235 
rect 152 235 153 236 
rect 152 236 153 237 
rect 152 237 153 238 
rect 152 238 153 239 
rect 152 239 153 240 
rect 152 240 153 241 
rect 152 243 153 244 
rect 152 244 153 245 
rect 152 245 153 246 
rect 152 246 153 247 
rect 152 247 153 248 
rect 152 248 153 249 
rect 152 249 153 250 
rect 152 250 153 251 
rect 152 251 153 252 
rect 152 252 153 253 
rect 152 253 153 254 
rect 152 254 153 255 
rect 152 255 153 256 
rect 152 256 153 257 
rect 152 257 153 258 
rect 152 258 153 259 
rect 152 259 153 260 
rect 152 260 153 261 
rect 152 261 153 262 
rect 152 262 153 263 
rect 152 263 153 264 
rect 152 267 153 268 
rect 152 268 153 269 
rect 152 273 153 274 
rect 152 275 153 276 
rect 152 276 153 277 
rect 152 278 153 279 
rect 152 279 153 280 
rect 152 280 153 281 
rect 152 281 153 282 
rect 152 282 153 283 
rect 152 283 153 284 
rect 152 284 153 285 
rect 152 285 153 286 
rect 152 286 153 287 
rect 152 287 153 288 
rect 152 288 153 289 
rect 152 290 153 291 
rect 152 293 153 294 
rect 152 305 153 306 
rect 152 308 153 309 
rect 152 310 153 311 
rect 152 312 153 313 
rect 153 1 154 2 
rect 153 3 154 4 
rect 153 8 154 9 
rect 153 17 154 18 
rect 153 18 154 19 
rect 153 20 154 21 
rect 153 23 154 24 
rect 153 25 154 26 
rect 153 33 154 34 
rect 153 36 154 37 
rect 153 38 154 39 
rect 153 40 154 41 
rect 153 50 154 51 
rect 153 118 154 119 
rect 153 129 154 130 
rect 153 134 154 135 
rect 153 136 154 137 
rect 153 145 154 146 
rect 153 152 154 153 
rect 153 153 154 154 
rect 153 161 154 162 
rect 153 165 154 166 
rect 153 184 154 185 
rect 153 193 154 194 
rect 153 226 154 227 
rect 153 232 154 233 
rect 153 233 154 234 
rect 153 263 154 264 
rect 153 267 154 268 
rect 153 273 154 274 
rect 153 275 154 276 
rect 153 278 154 279 
rect 153 289 154 290 
rect 153 290 154 291 
rect 153 293 154 294 
rect 153 305 154 306 
rect 153 308 154 309 
rect 153 310 154 311 
rect 153 312 154 313 
rect 154 1 155 2 
rect 154 3 155 4 
rect 154 8 155 9 
rect 154 17 155 18 
rect 154 20 155 21 
rect 154 23 155 24 
rect 154 33 155 34 
rect 154 36 155 37 
rect 154 38 155 39 
rect 154 40 155 41 
rect 154 50 155 51 
rect 154 53 155 54 
rect 154 54 155 55 
rect 154 55 155 56 
rect 154 66 155 67 
rect 154 69 155 70 
rect 154 71 155 72 
rect 154 98 155 99 
rect 154 99 155 100 
rect 154 100 155 101 
rect 154 101 155 102 
rect 154 102 155 103 
rect 154 103 155 104 
rect 154 104 155 105 
rect 154 118 155 119 
rect 154 129 155 130 
rect 154 131 155 132 
rect 154 134 155 135 
rect 154 136 155 137 
rect 154 145 155 146 
rect 154 152 155 153 
rect 154 161 155 162 
rect 154 165 155 166 
rect 154 184 155 185 
rect 154 193 155 194 
rect 154 210 155 211 
rect 154 211 155 212 
rect 154 212 155 213 
rect 154 213 155 214 
rect 154 214 155 215 
rect 154 215 155 216 
rect 154 226 155 227 
rect 154 232 155 233 
rect 154 244 155 245 
rect 154 245 155 246 
rect 154 258 155 259 
rect 154 263 155 264 
rect 154 267 155 268 
rect 154 273 155 274 
rect 154 275 155 276 
rect 154 278 155 279 
rect 154 280 155 281 
rect 154 289 155 290 
rect 154 293 155 294 
rect 154 305 155 306 
rect 154 308 155 309 
rect 154 310 155 311 
rect 154 312 155 313 
rect 155 1 156 2 
rect 155 3 156 4 
rect 155 8 156 9 
rect 155 17 156 18 
rect 155 20 156 21 
rect 155 23 156 24 
rect 155 33 156 34 
rect 155 36 156 37 
rect 155 38 156 39 
rect 155 40 156 41 
rect 155 50 156 51 
rect 155 55 156 56 
rect 155 66 156 67 
rect 155 69 156 70 
rect 155 71 156 72 
rect 155 104 156 105 
rect 155 118 156 119 
rect 155 129 156 130 
rect 155 131 156 132 
rect 155 134 156 135 
rect 155 136 156 137 
rect 155 145 156 146 
rect 155 152 156 153 
rect 155 161 156 162 
rect 155 165 156 166 
rect 155 184 156 185 
rect 155 193 156 194 
rect 155 210 156 211 
rect 155 226 156 227 
rect 155 232 156 233 
rect 155 244 156 245 
rect 155 248 156 249 
rect 155 258 156 259 
rect 155 263 156 264 
rect 155 273 156 274 
rect 155 275 156 276 
rect 155 278 156 279 
rect 155 280 156 281 
rect 155 289 156 290 
rect 155 293 156 294 
rect 155 305 156 306 
rect 155 308 156 309 
rect 155 310 156 311 
rect 155 312 156 313 
rect 156 1 157 2 
rect 156 3 157 4 
rect 156 8 157 9 
rect 156 17 157 18 
rect 156 20 157 21 
rect 156 23 157 24 
rect 156 33 157 34 
rect 156 36 157 37 
rect 156 38 157 39 
rect 156 40 157 41 
rect 156 50 157 51 
rect 156 53 157 54 
rect 156 55 157 56 
rect 156 66 157 67 
rect 156 69 157 70 
rect 156 71 157 72 
rect 156 104 157 105 
rect 156 118 157 119 
rect 156 129 157 130 
rect 156 131 157 132 
rect 156 134 157 135 
rect 156 136 157 137 
rect 156 145 157 146 
rect 156 152 157 153 
rect 156 161 157 162 
rect 156 165 157 166 
rect 156 184 157 185 
rect 156 193 157 194 
rect 156 210 157 211 
rect 156 226 157 227 
rect 156 232 157 233 
rect 156 244 157 245 
rect 156 248 157 249 
rect 156 258 157 259 
rect 156 263 157 264 
rect 156 273 157 274 
rect 156 275 157 276 
rect 156 278 157 279 
rect 156 280 157 281 
rect 156 289 157 290 
rect 156 293 157 294 
rect 156 305 157 306 
rect 156 308 157 309 
rect 156 310 157 311 
rect 156 312 157 313 
rect 157 1 158 2 
rect 157 3 158 4 
rect 157 8 158 9 
rect 157 17 158 18 
rect 157 20 158 21 
rect 157 23 158 24 
rect 157 33 158 34 
rect 157 36 158 37 
rect 157 38 158 39 
rect 157 40 158 41 
rect 157 50 158 51 
rect 157 53 158 54 
rect 157 55 158 56 
rect 157 66 158 67 
rect 157 69 158 70 
rect 157 71 158 72 
rect 157 104 158 105 
rect 157 118 158 119 
rect 157 129 158 130 
rect 157 131 158 132 
rect 157 134 158 135 
rect 157 136 158 137 
rect 157 145 158 146 
rect 157 152 158 153 
rect 157 161 158 162 
rect 157 162 158 163 
rect 157 165 158 166 
rect 157 184 158 185 
rect 157 193 158 194 
rect 157 210 158 211 
rect 157 226 158 227 
rect 157 232 158 233 
rect 157 244 158 245 
rect 157 248 158 249 
rect 157 258 158 259 
rect 157 263 158 264 
rect 157 273 158 274 
rect 157 275 158 276 
rect 157 278 158 279 
rect 157 280 158 281 
rect 157 289 158 290 
rect 157 293 158 294 
rect 157 305 158 306 
rect 157 308 158 309 
rect 157 310 158 311 
rect 157 312 158 313 
rect 158 1 159 2 
rect 158 3 159 4 
rect 158 8 159 9 
rect 158 17 159 18 
rect 158 20 159 21 
rect 158 23 159 24 
rect 158 33 159 34 
rect 158 36 159 37 
rect 158 38 159 39 
rect 158 40 159 41 
rect 158 50 159 51 
rect 158 53 159 54 
rect 158 55 159 56 
rect 158 66 159 67 
rect 158 69 159 70 
rect 158 71 159 72 
rect 158 104 159 105 
rect 158 118 159 119 
rect 158 129 159 130 
rect 158 131 159 132 
rect 158 134 159 135 
rect 158 136 159 137 
rect 158 145 159 146 
rect 158 152 159 153 
rect 158 162 159 163 
rect 158 165 159 166 
rect 158 184 159 185 
rect 158 193 159 194 
rect 158 210 159 211 
rect 158 226 159 227 
rect 158 232 159 233 
rect 158 244 159 245 
rect 158 248 159 249 
rect 158 258 159 259 
rect 158 263 159 264 
rect 158 273 159 274 
rect 158 275 159 276 
rect 158 278 159 279 
rect 158 280 159 281 
rect 158 289 159 290 
rect 158 293 159 294 
rect 158 305 159 306 
rect 158 308 159 309 
rect 158 310 159 311 
rect 158 312 159 313 
rect 159 1 160 2 
rect 159 3 160 4 
rect 159 8 160 9 
rect 159 11 160 12 
rect 159 17 160 18 
rect 159 20 160 21 
rect 159 23 160 24 
rect 159 33 160 34 
rect 159 36 160 37 
rect 159 38 160 39 
rect 159 40 160 41 
rect 159 46 160 47 
rect 159 50 160 51 
rect 159 53 160 54 
rect 159 55 160 56 
rect 159 66 160 67 
rect 159 69 160 70 
rect 159 71 160 72 
rect 159 118 160 119 
rect 159 129 160 130 
rect 159 131 160 132 
rect 159 134 160 135 
rect 159 136 160 137 
rect 159 139 160 140 
rect 159 145 160 146 
rect 159 152 160 153 
rect 159 162 160 163 
rect 159 165 160 166 
rect 159 184 160 185 
rect 159 190 160 191 
rect 159 193 160 194 
rect 159 210 160 211 
rect 159 219 160 220 
rect 159 226 160 227 
rect 159 232 160 233 
rect 159 238 160 239 
rect 159 244 160 245 
rect 159 248 160 249 
rect 159 251 160 252 
rect 159 258 160 259 
rect 159 263 160 264 
rect 159 270 160 271 
rect 159 273 160 274 
rect 159 275 160 276 
rect 159 278 160 279 
rect 159 280 160 281 
rect 159 286 160 287 
rect 159 289 160 290 
rect 159 293 160 294 
rect 159 305 160 306 
rect 159 308 160 309 
rect 159 310 160 311 
rect 159 312 160 313 
rect 160 1 161 2 
rect 160 3 161 4 
rect 160 8 161 9 
rect 160 11 161 12 
rect 160 16 161 17 
rect 160 17 161 18 
rect 160 20 161 21 
rect 160 23 161 24 
rect 160 32 161 33 
rect 160 33 161 34 
rect 160 36 161 37 
rect 160 38 161 39 
rect 160 40 161 41 
rect 160 46 161 47 
rect 160 50 161 51 
rect 160 53 161 54 
rect 160 55 161 56 
rect 160 66 161 67 
rect 160 69 161 70 
rect 160 71 161 72 
rect 160 97 161 98 
rect 160 98 161 99 
rect 160 99 161 100 
rect 160 100 161 101 
rect 160 101 161 102 
rect 160 102 161 103 
rect 160 103 161 104 
rect 160 104 161 105 
rect 160 118 161 119 
rect 160 128 161 129 
rect 160 129 161 130 
rect 160 131 161 132 
rect 160 134 161 135 
rect 160 136 161 137 
rect 160 139 161 140 
rect 160 145 161 146 
rect 160 152 161 153 
rect 160 162 161 163 
rect 160 165 161 166 
rect 160 184 161 185 
rect 160 185 161 186 
rect 160 190 161 191 
rect 160 192 161 193 
rect 160 193 161 194 
rect 160 210 161 211 
rect 160 219 161 220 
rect 160 226 161 227 
rect 160 232 161 233 
rect 160 238 161 239 
rect 160 240 161 241 
rect 160 241 161 242 
rect 160 242 161 243 
rect 160 243 161 244 
rect 160 244 161 245 
rect 160 248 161 249 
rect 160 251 161 252 
rect 160 258 161 259 
rect 160 263 161 264 
rect 160 270 161 271 
rect 160 273 161 274 
rect 160 275 161 276 
rect 160 278 161 279 
rect 160 280 161 281 
rect 160 281 161 282 
rect 160 286 161 287 
rect 160 288 161 289 
rect 160 289 161 290 
rect 160 293 161 294 
rect 160 305 161 306 
rect 160 308 161 309 
rect 160 310 161 311 
rect 160 312 161 313 
rect 161 1 162 2 
rect 161 3 162 4 
rect 161 8 162 9 
rect 161 11 162 12 
rect 161 12 162 13 
rect 161 13 162 14 
rect 161 14 162 15 
rect 161 15 162 16 
rect 161 16 162 17 
rect 161 20 162 21 
rect 161 23 162 24 
rect 161 25 162 26 
rect 161 26 162 27 
rect 161 27 162 28 
rect 161 28 162 29 
rect 161 29 162 30 
rect 161 30 162 31 
rect 161 31 162 32 
rect 161 32 162 33 
rect 161 36 162 37 
rect 161 38 162 39 
rect 161 40 162 41 
rect 161 46 162 47 
rect 161 47 162 48 
rect 161 48 162 49 
rect 161 50 162 51 
rect 161 53 162 54 
rect 161 55 162 56 
rect 161 66 162 67 
rect 161 69 162 70 
rect 161 71 162 72 
rect 161 75 162 76 
rect 161 76 162 77 
rect 161 77 162 78 
rect 161 78 162 79 
rect 161 79 162 80 
rect 161 80 162 81 
rect 161 81 162 82 
rect 161 82 162 83 
rect 161 83 162 84 
rect 161 84 162 85 
rect 161 85 162 86 
rect 161 86 162 87 
rect 161 87 162 88 
rect 161 88 162 89 
rect 161 89 162 90 
rect 161 90 162 91 
rect 161 91 162 92 
rect 161 92 162 93 
rect 161 93 162 94 
rect 161 94 162 95 
rect 161 97 162 98 
rect 161 104 162 105 
rect 161 105 162 106 
rect 161 106 162 107 
rect 161 107 162 108 
rect 161 108 162 109 
rect 161 109 162 110 
rect 161 110 162 111 
rect 161 111 162 112 
rect 161 112 162 113 
rect 161 113 162 114 
rect 161 114 162 115 
rect 161 115 162 116 
rect 161 118 162 119 
rect 161 120 162 121 
rect 161 121 162 122 
rect 161 122 162 123 
rect 161 123 162 124 
rect 161 124 162 125 
rect 161 125 162 126 
rect 161 126 162 127 
rect 161 127 162 128 
rect 161 128 162 129 
rect 161 130 162 131 
rect 161 131 162 132 
rect 161 134 162 135 
rect 161 136 162 137 
rect 161 139 162 140 
rect 161 145 162 146 
rect 161 152 162 153 
rect 161 162 162 163 
rect 161 185 162 186 
rect 161 186 162 187 
rect 161 187 162 188 
rect 161 188 162 189 
rect 161 190 162 191 
rect 161 191 162 192 
rect 161 192 162 193 
rect 161 201 162 202 
rect 161 202 162 203 
rect 161 203 162 204 
rect 161 204 162 205 
rect 161 205 162 206 
rect 161 206 162 207 
rect 161 207 162 208 
rect 161 208 162 209 
rect 161 209 162 210 
rect 161 210 162 211 
rect 161 219 162 220 
rect 161 226 162 227 
rect 161 232 162 233 
rect 161 238 162 239 
rect 161 239 162 240 
rect 161 240 162 241 
rect 161 248 162 249 
rect 161 251 162 252 
rect 161 258 162 259 
rect 161 259 162 260 
rect 161 260 162 261 
rect 161 261 162 262 
rect 161 263 162 264 
rect 161 270 162 271 
rect 161 273 162 274 
rect 161 275 162 276 
rect 161 278 162 279 
rect 161 281 162 282 
rect 161 282 162 283 
rect 161 283 162 284 
rect 161 284 162 285 
rect 161 285 162 286 
rect 161 286 162 287 
rect 161 288 162 289 
rect 161 293 162 294 
rect 161 305 162 306 
rect 161 308 162 309 
rect 161 310 162 311 
rect 161 312 162 313 
rect 162 1 163 2 
rect 162 3 163 4 
rect 162 8 163 9 
rect 162 18 163 19 
rect 162 20 163 21 
rect 162 23 163 24 
rect 162 25 163 26 
rect 162 36 163 37 
rect 162 38 163 39 
rect 162 40 163 41 
rect 162 50 163 51 
rect 162 53 163 54 
rect 162 55 163 56 
rect 162 66 163 67 
rect 162 69 163 70 
rect 162 71 163 72 
rect 162 75 163 76 
rect 162 94 163 95 
rect 162 95 163 96 
rect 162 97 163 98 
rect 162 118 163 119 
rect 162 129 163 130 
rect 162 130 163 131 
rect 162 134 163 135 
rect 162 136 163 137 
rect 162 145 163 146 
rect 162 152 163 153 
rect 162 162 163 163 
rect 162 163 163 164 
rect 162 164 163 165 
rect 162 165 163 166 
rect 162 166 163 167 
rect 162 167 163 168 
rect 162 188 163 189 
rect 162 189 163 190 
rect 162 219 163 220 
rect 162 226 163 227 
rect 162 232 163 233 
rect 162 246 163 247 
rect 162 248 163 249 
rect 162 251 163 252 
rect 162 261 163 262 
rect 162 263 163 264 
rect 162 270 163 271 
rect 162 273 163 274 
rect 162 275 163 276 
rect 162 278 163 279 
rect 162 287 163 288 
rect 162 288 163 289 
rect 162 293 163 294 
rect 162 305 163 306 
rect 162 308 163 309 
rect 162 310 163 311 
rect 162 312 163 313 
rect 163 1 164 2 
rect 163 3 164 4 
rect 163 8 164 9 
rect 163 18 164 19 
rect 163 20 164 21 
rect 163 23 164 24 
rect 163 25 164 26 
rect 163 36 164 37 
rect 163 38 164 39 
rect 163 40 164 41 
rect 163 50 164 51 
rect 163 53 164 54 
rect 163 55 164 56 
rect 163 66 164 67 
rect 163 69 164 70 
rect 163 71 164 72 
rect 163 75 164 76 
rect 163 90 164 91 
rect 163 91 164 92 
rect 163 92 164 93 
rect 163 93 164 94 
rect 163 95 164 96 
rect 163 97 164 98 
rect 163 118 164 119 
rect 163 126 164 127 
rect 163 127 164 128 
rect 163 128 164 129 
rect 163 129 164 130 
rect 163 134 164 135 
rect 163 136 164 137 
rect 163 145 164 146 
rect 163 152 164 153 
rect 163 167 164 168 
rect 163 189 164 190 
rect 163 190 164 191 
rect 163 191 164 192 
rect 163 192 164 193 
rect 163 193 164 194 
rect 163 194 164 195 
rect 163 195 164 196 
rect 163 196 164 197 
rect 163 197 164 198 
rect 163 198 164 199 
rect 163 199 164 200 
rect 163 200 164 201 
rect 163 201 164 202 
rect 163 202 164 203 
rect 163 203 164 204 
rect 163 204 164 205 
rect 163 205 164 206 
rect 163 206 164 207 
rect 163 207 164 208 
rect 163 208 164 209 
rect 163 209 164 210 
rect 163 210 164 211 
rect 163 211 164 212 
rect 163 212 164 213 
rect 163 213 164 214 
rect 163 214 164 215 
rect 163 215 164 216 
rect 163 216 164 217 
rect 163 219 164 220 
rect 163 226 164 227 
rect 163 232 164 233 
rect 163 246 164 247 
rect 163 248 164 249 
rect 163 251 164 252 
rect 163 261 164 262 
rect 163 263 164 264 
rect 163 270 164 271 
rect 163 273 164 274 
rect 163 275 164 276 
rect 163 278 164 279 
rect 163 280 164 281 
rect 163 281 164 282 
rect 163 282 164 283 
rect 163 283 164 284 
rect 163 284 164 285 
rect 163 285 164 286 
rect 163 286 164 287 
rect 163 287 164 288 
rect 163 293 164 294 
rect 163 305 164 306 
rect 163 308 164 309 
rect 163 310 164 311 
rect 163 312 164 313 
rect 164 1 165 2 
rect 164 3 165 4 
rect 164 8 165 9 
rect 164 16 165 17 
rect 164 18 165 19 
rect 164 20 165 21 
rect 164 23 165 24 
rect 164 36 165 37 
rect 164 38 165 39 
rect 164 40 165 41 
rect 164 50 165 51 
rect 164 53 165 54 
rect 164 55 165 56 
rect 164 66 165 67 
rect 164 69 165 70 
rect 164 71 165 72 
rect 164 75 165 76 
rect 164 90 165 91 
rect 164 97 165 98 
rect 164 99 165 100 
rect 164 100 165 101 
rect 164 101 165 102 
rect 164 102 165 103 
rect 164 103 165 104 
rect 164 104 165 105 
rect 164 105 165 106 
rect 164 106 165 107 
rect 164 107 165 108 
rect 164 108 165 109 
rect 164 109 165 110 
rect 164 110 165 111 
rect 164 111 165 112 
rect 164 112 165 113 
rect 164 113 165 114 
rect 164 114 165 115 
rect 164 115 165 116 
rect 164 118 165 119 
rect 164 126 165 127 
rect 164 134 165 135 
rect 164 136 165 137 
rect 164 138 165 139 
rect 164 139 165 140 
rect 164 140 165 141 
rect 164 141 165 142 
rect 164 142 165 143 
rect 164 143 165 144 
rect 164 145 165 146 
rect 164 152 165 153 
rect 164 167 165 168 
rect 164 216 165 217 
rect 164 219 165 220 
rect 164 226 165 227 
rect 164 230 165 231 
rect 164 232 165 233 
rect 164 246 165 247 
rect 164 248 165 249 
rect 164 259 165 260 
rect 164 261 165 262 
rect 164 263 165 264 
rect 164 270 165 271 
rect 164 273 165 274 
rect 164 275 165 276 
rect 164 278 165 279 
rect 164 280 165 281 
rect 164 293 165 294 
rect 164 305 165 306 
rect 164 308 165 309 
rect 164 310 165 311 
rect 164 312 165 313 
rect 165 1 166 2 
rect 165 3 166 4 
rect 165 8 166 9 
rect 165 16 166 17 
rect 165 18 166 19 
rect 165 20 166 21 
rect 165 23 166 24 
rect 165 36 166 37 
rect 165 38 166 39 
rect 165 40 166 41 
rect 165 50 166 51 
rect 165 53 166 54 
rect 165 55 166 56 
rect 165 66 166 67 
rect 165 69 166 70 
rect 165 71 166 72 
rect 165 75 166 76 
rect 165 90 166 91 
rect 165 97 166 98 
rect 165 115 166 116 
rect 165 118 166 119 
rect 165 126 166 127 
rect 165 134 166 135 
rect 165 136 166 137 
rect 165 143 166 144 
rect 165 145 166 146 
rect 165 152 166 153 
rect 165 154 166 155 
rect 165 155 166 156 
rect 165 156 166 157 
rect 165 157 166 158 
rect 165 158 166 159 
rect 165 159 166 160 
rect 165 160 166 161 
rect 165 161 166 162 
rect 165 162 166 163 
rect 165 163 166 164 
rect 165 165 166 166 
rect 165 167 166 168 
rect 165 169 166 170 
rect 165 170 166 171 
rect 165 171 166 172 
rect 165 172 166 173 
rect 165 173 166 174 
rect 165 174 166 175 
rect 165 175 166 176 
rect 165 176 166 177 
rect 165 177 166 178 
rect 165 178 166 179 
rect 165 179 166 180 
rect 165 180 166 181 
rect 165 181 166 182 
rect 165 182 166 183 
rect 165 183 166 184 
rect 165 184 166 185 
rect 165 185 166 186 
rect 165 186 166 187 
rect 165 187 166 188 
rect 165 188 166 189 
rect 165 189 166 190 
rect 165 190 166 191 
rect 165 191 166 192 
rect 165 192 166 193 
rect 165 193 166 194 
rect 165 194 166 195 
rect 165 197 166 198 
rect 165 199 166 200 
rect 165 200 166 201 
rect 165 212 166 213 
rect 165 213 166 214 
rect 165 216 166 217 
rect 165 219 166 220 
rect 165 226 166 227 
rect 165 230 166 231 
rect 165 232 166 233 
rect 165 246 166 247 
rect 165 248 166 249 
rect 165 259 166 260 
rect 165 261 166 262 
rect 165 263 166 264 
rect 165 270 166 271 
rect 165 273 166 274 
rect 165 275 166 276 
rect 165 278 166 279 
rect 165 280 166 281 
rect 165 293 166 294 
rect 165 305 166 306 
rect 165 308 166 309 
rect 165 310 166 311 
rect 165 312 166 313 
rect 166 1 167 2 
rect 166 3 167 4 
rect 166 8 167 9 
rect 166 11 167 12 
rect 166 12 167 13 
rect 166 13 167 14 
rect 166 14 167 15 
rect 166 15 167 16 
rect 166 16 167 17 
rect 166 18 167 19 
rect 166 20 167 21 
rect 166 23 167 24 
rect 166 36 167 37 
rect 166 38 167 39 
rect 166 40 167 41 
rect 166 50 167 51 
rect 166 53 167 54 
rect 166 55 167 56 
rect 166 65 167 66 
rect 166 66 167 67 
rect 166 69 167 70 
rect 166 71 167 72 
rect 166 75 167 76 
rect 166 90 167 91 
rect 166 97 167 98 
rect 166 103 167 104 
rect 166 104 167 105 
rect 166 118 167 119 
rect 166 126 167 127 
rect 166 134 167 135 
rect 166 136 167 137 
rect 166 143 167 144 
rect 166 145 167 146 
rect 166 152 167 153 
rect 166 165 167 166 
rect 166 167 167 168 
rect 166 169 167 170 
rect 166 196 167 197 
rect 166 197 167 198 
rect 166 199 167 200 
rect 166 212 167 213 
rect 166 216 167 217 
rect 166 219 167 220 
rect 166 226 167 227 
rect 166 230 167 231 
rect 166 232 167 233 
rect 166 246 167 247 
rect 166 248 167 249 
rect 166 259 167 260 
rect 166 261 167 262 
rect 166 263 167 264 
rect 166 273 167 274 
rect 166 275 167 276 
rect 166 278 167 279 
rect 166 280 167 281 
rect 166 282 167 283 
rect 166 283 167 284 
rect 166 284 167 285 
rect 166 285 167 286 
rect 166 286 167 287 
rect 166 287 167 288 
rect 166 288 167 289 
rect 166 293 167 294 
rect 166 305 167 306 
rect 166 308 167 309 
rect 166 310 167 311 
rect 166 312 167 313 
rect 167 1 168 2 
rect 167 3 168 4 
rect 167 8 168 9 
rect 167 11 168 12 
rect 167 18 168 19 
rect 167 20 168 21 
rect 167 23 168 24 
rect 167 36 168 37 
rect 167 38 168 39 
rect 167 40 168 41 
rect 167 50 168 51 
rect 167 53 168 54 
rect 167 55 168 56 
rect 167 69 168 70 
rect 167 71 168 72 
rect 167 75 168 76 
rect 167 90 168 91 
rect 167 97 168 98 
rect 167 104 168 105 
rect 167 118 168 119 
rect 167 126 168 127 
rect 167 134 168 135 
rect 167 136 168 137 
rect 167 143 168 144 
rect 167 145 168 146 
rect 167 152 168 153 
rect 167 165 168 166 
rect 167 167 168 168 
rect 167 174 168 175 
rect 167 175 168 176 
rect 167 176 168 177 
rect 167 177 168 178 
rect 167 178 168 179 
rect 167 179 168 180 
rect 167 180 168 181 
rect 167 181 168 182 
rect 167 182 168 183 
rect 167 183 168 184 
rect 167 184 168 185 
rect 167 185 168 186 
rect 167 186 168 187 
rect 167 187 168 188 
rect 167 188 168 189 
rect 167 189 168 190 
rect 167 190 168 191 
rect 167 191 168 192 
rect 167 192 168 193 
rect 167 193 168 194 
rect 167 194 168 195 
rect 167 195 168 196 
rect 167 196 168 197 
rect 167 198 168 199 
rect 167 199 168 200 
rect 167 212 168 213 
rect 167 216 168 217 
rect 167 219 168 220 
rect 167 226 168 227 
rect 167 230 168 231 
rect 167 232 168 233 
rect 167 246 168 247 
rect 167 248 168 249 
rect 167 259 168 260 
rect 167 261 168 262 
rect 167 263 168 264 
rect 167 273 168 274 
rect 167 275 168 276 
rect 167 278 168 279 
rect 167 280 168 281 
rect 167 288 168 289 
rect 167 293 168 294 
rect 167 305 168 306 
rect 167 308 168 309 
rect 167 310 168 311 
rect 167 312 168 313 
rect 168 1 169 2 
rect 168 3 169 4 
rect 168 8 169 9 
rect 168 11 169 12 
rect 168 18 169 19 
rect 168 20 169 21 
rect 168 23 169 24 
rect 168 36 169 37 
rect 168 38 169 39 
rect 168 40 169 41 
rect 168 50 169 51 
rect 168 53 169 54 
rect 168 55 169 56 
rect 168 59 169 60 
rect 168 60 169 61 
rect 168 61 169 62 
rect 168 62 169 63 
rect 168 63 169 64 
rect 168 64 169 65 
rect 168 65 169 66 
rect 168 66 169 67 
rect 168 67 169 68 
rect 168 68 169 69 
rect 168 69 169 70 
rect 168 71 169 72 
rect 168 75 169 76 
rect 168 89 169 90 
rect 168 90 169 91 
rect 168 97 169 98 
rect 168 104 169 105 
rect 168 107 169 108 
rect 168 108 169 109 
rect 168 109 169 110 
rect 168 110 169 111 
rect 168 111 169 112 
rect 168 112 169 113 
rect 168 118 169 119 
rect 168 126 169 127 
rect 168 134 169 135 
rect 168 136 169 137 
rect 168 143 169 144 
rect 168 145 169 146 
rect 168 152 169 153 
rect 168 155 169 156 
rect 168 156 169 157 
rect 168 157 169 158 
rect 168 158 169 159 
rect 168 159 169 160 
rect 168 160 169 161 
rect 168 165 169 166 
rect 168 167 169 168 
rect 168 174 169 175 
rect 168 197 169 198 
rect 168 198 169 199 
rect 168 212 169 213 
rect 168 216 169 217 
rect 168 219 169 220 
rect 168 226 169 227 
rect 168 230 169 231 
rect 168 232 169 233 
rect 168 246 169 247 
rect 168 248 169 249 
rect 168 259 169 260 
rect 168 261 169 262 
rect 168 263 169 264 
rect 168 273 169 274 
rect 168 275 169 276 
rect 168 278 169 279 
rect 168 280 169 281 
rect 168 282 169 283 
rect 168 283 169 284 
rect 168 288 169 289 
rect 168 293 169 294 
rect 168 305 169 306 
rect 168 308 169 309 
rect 168 310 169 311 
rect 168 312 169 313 
rect 169 1 170 2 
rect 169 3 170 4 
rect 169 8 170 9 
rect 169 11 170 12 
rect 169 18 170 19 
rect 169 20 170 21 
rect 169 23 170 24 
rect 169 36 170 37 
rect 169 38 170 39 
rect 169 40 170 41 
rect 169 50 170 51 
rect 169 53 170 54 
rect 169 55 170 56 
rect 169 59 170 60 
rect 169 71 170 72 
rect 169 75 170 76 
rect 169 88 170 89 
rect 169 89 170 90 
rect 169 97 170 98 
rect 169 104 170 105 
rect 169 107 170 108 
rect 169 112 170 113 
rect 169 113 170 114 
rect 169 118 170 119 
rect 169 126 170 127 
rect 169 134 170 135 
rect 169 136 170 137 
rect 169 145 170 146 
rect 169 152 170 153 
rect 169 155 170 156 
rect 169 160 170 161 
rect 169 161 170 162 
rect 169 165 170 166 
rect 169 167 170 168 
rect 169 174 170 175 
rect 169 197 170 198 
rect 169 212 170 213 
rect 169 216 170 217 
rect 169 226 170 227 
rect 169 230 170 231 
rect 169 232 170 233 
rect 169 246 170 247 
rect 169 248 170 249 
rect 169 257 170 258 
rect 169 258 170 259 
rect 169 259 170 260 
rect 169 261 170 262 
rect 169 263 170 264 
rect 169 273 170 274 
rect 169 275 170 276 
rect 169 278 170 279 
rect 169 280 170 281 
rect 169 283 170 284 
rect 169 288 170 289 
rect 169 289 170 290 
rect 169 293 170 294 
rect 169 305 170 306 
rect 169 308 170 309 
rect 169 310 170 311 
rect 169 312 170 313 
rect 170 1 171 2 
rect 170 3 171 4 
rect 170 8 171 9 
rect 170 11 171 12 
rect 170 18 171 19 
rect 170 20 171 21 
rect 170 23 171 24 
rect 170 36 171 37 
rect 170 38 171 39 
rect 170 40 171 41 
rect 170 50 171 51 
rect 170 53 171 54 
rect 170 55 171 56 
rect 170 59 171 60 
rect 170 66 171 67 
rect 170 67 171 68 
rect 170 68 171 69 
rect 170 69 171 70 
rect 170 71 171 72 
rect 170 75 171 76 
rect 170 88 171 89 
rect 170 97 171 98 
rect 170 104 171 105 
rect 170 107 171 108 
rect 170 113 171 114 
rect 170 114 171 115 
rect 170 115 171 116 
rect 170 118 171 119 
rect 170 126 171 127 
rect 170 134 171 135 
rect 170 136 171 137 
rect 170 145 171 146 
rect 170 152 171 153 
rect 170 155 171 156 
rect 170 161 171 162 
rect 170 165 171 166 
rect 170 167 171 168 
rect 170 174 171 175 
rect 170 197 171 198 
rect 170 212 171 213 
rect 170 216 171 217 
rect 170 226 171 227 
rect 170 230 171 231 
rect 170 232 171 233 
rect 170 246 171 247 
rect 170 248 171 249 
rect 170 257 171 258 
rect 170 261 171 262 
rect 170 263 171 264 
rect 170 273 171 274 
rect 170 275 171 276 
rect 170 278 171 279 
rect 170 280 171 281 
rect 170 283 171 284 
rect 170 289 171 290 
rect 170 293 171 294 
rect 170 305 171 306 
rect 170 308 171 309 
rect 170 310 171 311 
rect 170 312 171 313 
rect 171 1 172 2 
rect 171 3 172 4 
rect 171 8 172 9 
rect 171 18 172 19 
rect 171 20 172 21 
rect 171 23 172 24 
rect 171 36 172 37 
rect 171 38 172 39 
rect 171 40 172 41 
rect 171 50 172 51 
rect 171 53 172 54 
rect 171 55 172 56 
rect 171 69 172 70 
rect 171 71 172 72 
rect 171 88 172 89 
rect 171 97 172 98 
rect 171 104 172 105 
rect 171 115 172 116 
rect 171 118 172 119 
rect 171 134 172 135 
rect 171 136 172 137 
rect 171 145 172 146 
rect 171 152 172 153 
rect 171 161 172 162 
rect 171 165 172 166 
rect 171 167 172 168 
rect 171 197 172 198 
rect 171 212 172 213 
rect 171 216 172 217 
rect 171 226 172 227 
rect 171 230 172 231 
rect 171 232 172 233 
rect 171 246 172 247 
rect 171 248 172 249 
rect 171 257 172 258 
rect 171 261 172 262 
rect 171 263 172 264 
rect 171 273 172 274 
rect 171 275 172 276 
rect 171 278 172 279 
rect 171 280 172 281 
rect 171 289 172 290 
rect 171 293 172 294 
rect 171 305 172 306 
rect 171 308 172 309 
rect 171 310 172 311 
rect 171 312 172 313 
rect 172 1 173 2 
rect 172 3 173 4 
rect 172 8 173 9 
rect 172 18 173 19 
rect 172 20 173 21 
rect 172 23 173 24 
rect 172 36 173 37 
rect 172 38 173 39 
rect 172 40 173 41 
rect 172 50 173 51 
rect 172 53 173 54 
rect 172 55 173 56 
rect 172 69 173 70 
rect 172 71 173 72 
rect 172 88 173 89 
rect 172 97 173 98 
rect 172 104 173 105 
rect 172 115 173 116 
rect 172 118 173 119 
rect 172 134 173 135 
rect 172 136 173 137 
rect 172 145 173 146 
rect 172 152 173 153 
rect 172 161 173 162 
rect 172 165 173 166 
rect 172 167 173 168 
rect 172 197 173 198 
rect 172 212 173 213 
rect 172 216 173 217 
rect 172 226 173 227 
rect 172 230 173 231 
rect 172 232 173 233 
rect 172 246 173 247 
rect 172 248 173 249 
rect 172 257 173 258 
rect 172 261 173 262 
rect 172 263 173 264 
rect 172 273 173 274 
rect 172 275 173 276 
rect 172 278 173 279 
rect 172 280 173 281 
rect 172 289 173 290 
rect 172 293 173 294 
rect 172 305 173 306 
rect 172 308 173 309 
rect 172 310 173 311 
rect 172 312 173 313 
rect 173 1 174 2 
rect 173 3 174 4 
rect 173 8 174 9 
rect 173 18 174 19 
rect 173 20 174 21 
rect 173 23 174 24 
rect 173 36 174 37 
rect 173 38 174 39 
rect 173 40 174 41 
rect 173 50 174 51 
rect 173 53 174 54 
rect 173 55 174 56 
rect 173 69 174 70 
rect 173 71 174 72 
rect 173 88 174 89 
rect 173 97 174 98 
rect 173 104 174 105 
rect 173 115 174 116 
rect 173 118 174 119 
rect 173 134 174 135 
rect 173 136 174 137 
rect 173 145 174 146 
rect 173 152 174 153 
rect 173 161 174 162 
rect 173 165 174 166 
rect 173 167 174 168 
rect 173 197 174 198 
rect 173 212 174 213 
rect 173 216 174 217 
rect 173 226 174 227 
rect 173 230 174 231 
rect 173 232 174 233 
rect 173 246 174 247 
rect 173 248 174 249 
rect 173 257 174 258 
rect 173 261 174 262 
rect 173 263 174 264 
rect 173 273 174 274 
rect 173 275 174 276 
rect 173 278 174 279 
rect 173 280 174 281 
rect 173 289 174 290 
rect 173 293 174 294 
rect 173 305 174 306 
rect 173 308 174 309 
rect 173 310 174 311 
rect 173 312 174 313 
rect 174 1 175 2 
rect 174 3 175 4 
rect 174 8 175 9 
rect 174 18 175 19 
rect 174 20 175 21 
rect 174 23 175 24 
rect 174 36 175 37 
rect 174 38 175 39 
rect 174 40 175 41 
rect 174 50 175 51 
rect 174 53 175 54 
rect 174 55 175 56 
rect 174 69 175 70 
rect 174 71 175 72 
rect 174 88 175 89 
rect 174 97 175 98 
rect 174 104 175 105 
rect 174 115 175 116 
rect 174 118 175 119 
rect 174 134 175 135 
rect 174 136 175 137 
rect 174 145 175 146 
rect 174 152 175 153 
rect 174 161 175 162 
rect 174 165 175 166 
rect 174 167 175 168 
rect 174 197 175 198 
rect 174 212 175 213 
rect 174 216 175 217 
rect 174 226 175 227 
rect 174 230 175 231 
rect 174 232 175 233 
rect 174 246 175 247 
rect 174 248 175 249 
rect 174 257 175 258 
rect 174 261 175 262 
rect 174 263 175 264 
rect 174 273 175 274 
rect 174 275 175 276 
rect 174 278 175 279 
rect 174 280 175 281 
rect 174 289 175 290 
rect 174 293 175 294 
rect 174 305 175 306 
rect 174 308 175 309 
rect 174 310 175 311 
rect 174 312 175 313 
rect 175 1 176 2 
rect 175 3 176 4 
rect 175 8 176 9 
rect 175 11 176 12 
rect 175 18 176 19 
rect 175 20 176 21 
rect 175 23 176 24 
rect 175 30 176 31 
rect 175 36 176 37 
rect 175 38 176 39 
rect 175 40 176 41 
rect 175 50 176 51 
rect 175 53 176 54 
rect 175 55 176 56 
rect 175 62 176 63 
rect 175 69 176 70 
rect 175 71 176 72 
rect 175 88 176 89 
rect 175 91 176 92 
rect 175 97 176 98 
rect 175 104 176 105 
rect 175 107 176 108 
rect 175 113 176 114 
rect 175 115 176 116 
rect 175 118 176 119 
rect 175 129 176 130 
rect 175 130 176 131 
rect 175 131 176 132 
rect 175 132 176 133 
rect 175 133 176 134 
rect 175 134 176 135 
rect 175 136 176 137 
rect 175 145 176 146 
rect 175 152 176 153 
rect 175 155 176 156 
rect 175 161 176 162 
rect 175 165 176 166 
rect 175 167 176 168 
rect 175 197 176 198 
rect 175 212 176 213 
rect 175 216 176 217 
rect 175 226 176 227 
rect 175 230 176 231 
rect 175 232 176 233 
rect 175 238 176 239 
rect 175 246 176 247 
rect 175 248 176 249 
rect 175 257 176 258 
rect 175 261 176 262 
rect 175 263 176 264 
rect 175 273 176 274 
rect 175 275 176 276 
rect 175 278 176 279 
rect 175 280 176 281 
rect 175 289 176 290 
rect 175 293 176 294 
rect 175 305 176 306 
rect 175 308 176 309 
rect 175 310 176 311 
rect 175 312 176 313 
rect 176 1 177 2 
rect 176 3 177 4 
rect 176 8 177 9 
rect 176 11 177 12 
rect 176 18 177 19 
rect 176 20 177 21 
rect 176 23 177 24 
rect 176 30 177 31 
rect 176 32 177 33 
rect 176 33 177 34 
rect 176 34 177 35 
rect 176 36 177 37 
rect 176 38 177 39 
rect 176 50 177 51 
rect 176 53 177 54 
rect 176 55 177 56 
rect 176 62 177 63 
rect 176 69 177 70 
rect 176 71 177 72 
rect 176 88 177 89 
rect 176 91 177 92 
rect 176 97 177 98 
rect 176 104 177 105 
rect 176 107 177 108 
rect 176 112 177 113 
rect 176 113 177 114 
rect 176 115 177 116 
rect 176 118 177 119 
rect 176 120 177 121 
rect 176 121 177 122 
rect 176 128 177 129 
rect 176 129 177 130 
rect 176 136 177 137 
rect 176 137 177 138 
rect 176 145 177 146 
rect 176 152 177 153 
rect 176 155 177 156 
rect 176 161 177 162 
rect 176 165 177 166 
rect 176 167 177 168 
rect 176 208 177 209 
rect 176 209 177 210 
rect 176 210 177 211 
rect 176 211 177 212 
rect 176 212 177 213 
rect 176 216 177 217 
rect 176 217 177 218 
rect 176 226 177 227 
rect 176 230 177 231 
rect 176 232 177 233 
rect 176 238 177 239 
rect 176 246 177 247 
rect 176 248 177 249 
rect 176 249 177 250 
rect 176 256 177 257 
rect 176 257 177 258 
rect 176 261 177 262 
rect 176 263 177 264 
rect 176 272 177 273 
rect 176 273 177 274 
rect 176 275 177 276 
rect 176 278 177 279 
rect 176 280 177 281 
rect 176 289 177 290 
rect 176 293 177 294 
rect 176 294 177 295 
rect 176 295 177 296 
rect 176 296 177 297 
rect 176 297 177 298 
rect 176 305 177 306 
rect 176 308 177 309 
rect 176 310 177 311 
rect 176 312 177 313 
rect 177 1 178 2 
rect 177 3 178 4 
rect 177 8 178 9 
rect 177 11 178 12 
rect 177 12 178 13 
rect 177 13 178 14 
rect 177 14 178 15 
rect 177 15 178 16 
rect 177 17 178 18 
rect 177 18 178 19 
rect 177 20 178 21 
rect 177 23 178 24 
rect 177 25 178 26 
rect 177 30 178 31 
rect 177 31 178 32 
rect 177 32 178 33 
rect 177 36 178 37 
rect 177 38 178 39 
rect 177 47 178 48 
rect 177 48 178 49 
rect 177 50 178 51 
rect 177 53 178 54 
rect 177 55 178 56 
rect 177 57 178 58 
rect 177 58 178 59 
rect 177 59 178 60 
rect 177 60 178 61 
rect 177 61 178 62 
rect 177 62 178 63 
rect 177 71 178 72 
rect 177 73 178 74 
rect 177 74 178 75 
rect 177 87 178 88 
rect 177 88 178 89 
rect 177 91 178 92 
rect 177 92 178 93 
rect 177 93 178 94 
rect 177 94 178 95 
rect 177 97 178 98 
rect 177 104 178 105 
rect 177 107 178 108 
rect 177 108 178 109 
rect 177 109 178 110 
rect 177 110 178 111 
rect 177 111 178 112 
rect 177 112 178 113 
rect 177 115 178 116 
rect 177 118 178 119 
rect 177 121 178 122 
rect 177 122 178 123 
rect 177 123 178 124 
rect 177 124 178 125 
rect 177 125 178 126 
rect 177 126 178 127 
rect 177 127 178 128 
rect 177 128 178 129 
rect 177 137 178 138 
rect 177 145 178 146 
rect 177 147 178 148 
rect 177 148 178 149 
rect 177 149 178 150 
rect 177 150 178 151 
rect 177 151 178 152 
rect 177 152 178 153 
rect 177 155 178 156 
rect 177 161 178 162 
rect 177 165 178 166 
rect 177 167 178 168 
rect 177 169 178 170 
rect 177 170 178 171 
rect 177 171 178 172 
rect 177 172 178 173 
rect 177 173 178 174 
rect 177 174 178 175 
rect 177 175 178 176 
rect 177 176 178 177 
rect 177 177 178 178 
rect 177 178 178 179 
rect 177 179 178 180 
rect 177 180 178 181 
rect 177 181 178 182 
rect 177 182 178 183 
rect 177 183 178 184 
rect 177 184 178 185 
rect 177 185 178 186 
rect 177 186 178 187 
rect 177 187 178 188 
rect 177 188 178 189 
rect 177 189 178 190 
rect 177 190 178 191 
rect 177 191 178 192 
rect 177 192 178 193 
rect 177 193 178 194 
rect 177 194 178 195 
rect 177 195 178 196 
rect 177 196 178 197 
rect 177 197 178 198 
rect 177 198 178 199 
rect 177 199 178 200 
rect 177 200 178 201 
rect 177 201 178 202 
rect 177 202 178 203 
rect 177 203 178 204 
rect 177 204 178 205 
rect 177 205 178 206 
rect 177 206 178 207 
rect 177 207 178 208 
rect 177 208 178 209 
rect 177 217 178 218 
rect 177 218 178 219 
rect 177 219 178 220 
rect 177 220 178 221 
rect 177 221 178 222 
rect 177 226 178 227 
rect 177 229 178 230 
rect 177 230 178 231 
rect 177 232 178 233 
rect 177 235 178 236 
rect 177 236 178 237 
rect 177 237 178 238 
rect 177 238 178 239 
rect 177 246 178 247 
rect 177 249 178 250 
rect 177 251 178 252 
rect 177 252 178 253 
rect 177 253 178 254 
rect 177 254 178 255 
rect 177 255 178 256 
rect 177 256 178 257 
rect 177 261 178 262 
rect 177 263 178 264 
rect 177 272 178 273 
rect 177 274 178 275 
rect 177 275 178 276 
rect 177 278 178 279 
rect 177 280 178 281 
rect 177 289 178 290 
rect 177 290 178 291 
rect 177 291 178 292 
rect 177 292 178 293 
rect 177 297 178 298 
rect 177 298 178 299 
rect 177 305 178 306 
rect 177 308 178 309 
rect 177 310 178 311 
rect 177 312 178 313 
rect 178 1 179 2 
rect 178 3 179 4 
rect 178 8 179 9 
rect 178 15 179 16 
rect 178 17 179 18 
rect 178 20 179 21 
rect 178 23 179 24 
rect 178 25 179 26 
rect 178 36 179 37 
rect 178 38 179 39 
rect 178 47 179 48 
rect 178 50 179 51 
rect 178 53 179 54 
rect 178 55 179 56 
rect 178 71 179 72 
rect 178 74 179 75 
rect 178 87 179 88 
rect 178 97 179 98 
rect 178 104 179 105 
rect 178 115 179 116 
rect 178 118 179 119 
rect 178 137 179 138 
rect 178 145 179 146 
rect 178 147 179 148 
rect 178 155 179 156 
rect 178 161 179 162 
rect 178 165 179 166 
rect 178 167 179 168 
rect 178 210 179 211 
rect 178 221 179 222 
rect 178 226 179 227 
rect 178 229 179 230 
rect 178 232 179 233 
rect 178 235 179 236 
rect 178 246 179 247 
rect 178 249 179 250 
rect 178 251 179 252 
rect 178 263 179 264 
rect 178 272 179 273 
rect 178 274 179 275 
rect 178 278 179 279 
rect 178 280 179 281 
rect 178 282 179 283 
rect 178 292 179 293 
rect 178 298 179 299 
rect 178 305 179 306 
rect 178 308 179 309 
rect 178 310 179 311 
rect 178 312 179 313 
rect 179 1 180 2 
rect 179 3 180 4 
rect 179 8 180 9 
rect 179 15 180 16 
rect 179 17 180 18 
rect 179 20 180 21 
rect 179 23 180 24 
rect 179 25 180 26 
rect 179 36 180 37 
rect 179 38 180 39 
rect 179 47 180 48 
rect 179 50 180 51 
rect 179 53 180 54 
rect 179 55 180 56 
rect 179 66 180 67 
rect 179 67 180 68 
rect 179 68 180 69 
rect 179 69 180 70 
rect 179 71 180 72 
rect 179 74 180 75 
rect 179 77 180 78 
rect 179 78 180 79 
rect 179 79 180 80 
rect 179 80 180 81 
rect 179 81 180 82 
rect 179 82 180 83 
rect 179 83 180 84 
rect 179 84 180 85 
rect 179 87 180 88 
rect 179 97 180 98 
rect 179 104 180 105 
rect 179 115 180 116 
rect 179 118 180 119 
rect 179 137 180 138 
rect 179 145 180 146 
rect 179 147 180 148 
rect 179 155 180 156 
rect 179 161 180 162 
rect 179 165 180 166 
rect 179 167 180 168 
rect 179 194 180 195 
rect 179 210 180 211 
rect 179 221 180 222 
rect 179 226 180 227 
rect 179 229 180 230 
rect 179 232 180 233 
rect 179 235 180 236 
rect 179 246 180 247 
rect 179 249 180 250 
rect 179 251 180 252 
rect 179 263 180 264 
rect 179 272 180 273 
rect 179 274 180 275 
rect 179 278 180 279 
rect 179 280 180 281 
rect 179 282 180 283 
rect 179 292 180 293 
rect 179 298 180 299 
rect 179 305 180 306 
rect 179 308 180 309 
rect 179 310 180 311 
rect 179 312 180 313 
rect 180 1 181 2 
rect 180 3 181 4 
rect 180 8 181 9 
rect 180 15 181 16 
rect 180 17 181 18 
rect 180 20 181 21 
rect 180 23 181 24 
rect 180 25 181 26 
rect 180 36 181 37 
rect 180 38 181 39 
rect 180 47 181 48 
rect 180 50 181 51 
rect 180 53 181 54 
rect 180 55 181 56 
rect 180 71 181 72 
rect 180 74 181 75 
rect 180 84 181 85 
rect 180 85 181 86 
rect 180 87 181 88 
rect 180 97 181 98 
rect 180 104 181 105 
rect 180 115 181 116 
rect 180 118 181 119 
rect 180 137 181 138 
rect 180 145 181 146 
rect 180 147 181 148 
rect 180 155 181 156 
rect 180 161 181 162 
rect 180 165 181 166 
rect 180 167 181 168 
rect 180 194 181 195 
rect 180 210 181 211 
rect 180 221 181 222 
rect 180 226 181 227 
rect 180 229 181 230 
rect 180 232 181 233 
rect 180 235 181 236 
rect 180 246 181 247 
rect 180 249 181 250 
rect 180 263 181 264 
rect 180 272 181 273 
rect 180 274 181 275 
rect 180 278 181 279 
rect 180 280 181 281 
rect 180 282 181 283 
rect 180 292 181 293 
rect 180 293 181 294 
rect 180 298 181 299 
rect 180 305 181 306 
rect 180 308 181 309 
rect 180 310 181 311 
rect 180 312 181 313 
rect 181 1 182 2 
rect 181 3 182 4 
rect 181 8 182 9 
rect 181 15 182 16 
rect 181 17 182 18 
rect 181 20 182 21 
rect 181 21 182 22 
rect 181 23 182 24 
rect 181 25 182 26 
rect 181 26 182 27 
rect 181 27 182 28 
rect 181 28 182 29 
rect 181 29 182 30 
rect 181 30 182 31 
rect 181 31 182 32 
rect 181 32 182 33 
rect 181 36 182 37 
rect 181 38 182 39 
rect 181 43 182 44 
rect 181 44 182 45 
rect 181 45 182 46 
rect 181 46 182 47 
rect 181 47 182 48 
rect 181 50 182 51 
rect 181 53 182 54 
rect 181 55 182 56 
rect 181 56 182 57 
rect 181 57 182 58 
rect 181 58 182 59 
rect 181 59 182 60 
rect 181 60 182 61 
rect 181 61 182 62 
rect 181 62 182 63 
rect 181 63 182 64 
rect 181 64 182 65 
rect 181 65 182 66 
rect 181 66 182 67 
rect 181 67 182 68 
rect 181 68 182 69 
rect 181 69 182 70 
rect 181 71 182 72 
rect 181 74 182 75 
rect 181 75 182 76 
rect 181 76 182 77 
rect 181 77 182 78 
rect 181 78 182 79 
rect 181 79 182 80 
rect 181 80 182 81 
rect 181 81 182 82 
rect 181 82 182 83 
rect 181 83 182 84 
rect 181 85 182 86 
rect 181 87 182 88 
rect 181 97 182 98 
rect 181 104 182 105 
rect 181 105 182 106 
rect 181 106 182 107 
rect 181 107 182 108 
rect 181 108 182 109 
rect 181 109 182 110 
rect 181 110 182 111 
rect 181 115 182 116 
rect 181 118 182 119 
rect 181 137 182 138 
rect 181 138 182 139 
rect 181 139 182 140 
rect 181 140 182 141 
rect 181 141 182 142 
rect 181 142 182 143 
rect 181 145 182 146 
rect 181 147 182 148 
rect 181 155 182 156 
rect 181 161 182 162 
rect 181 165 182 166 
rect 181 167 182 168 
rect 181 168 182 169 
rect 181 177 182 178 
rect 181 178 182 179 
rect 181 179 182 180 
rect 181 180 182 181 
rect 181 181 182 182 
rect 181 182 182 183 
rect 181 183 182 184 
rect 181 184 182 185 
rect 181 185 182 186 
rect 181 186 182 187 
rect 181 187 182 188 
rect 181 188 182 189 
rect 181 189 182 190 
rect 181 190 182 191 
rect 181 191 182 192 
rect 181 192 182 193 
rect 181 193 182 194 
rect 181 194 182 195 
rect 181 206 182 207 
rect 181 207 182 208 
rect 181 208 182 209 
rect 181 209 182 210 
rect 181 210 182 211 
rect 181 221 182 222 
rect 181 222 182 223 
rect 181 225 182 226 
rect 181 226 182 227 
rect 181 229 182 230 
rect 181 232 182 233 
rect 181 235 182 236 
rect 181 241 182 242 
rect 181 242 182 243 
rect 181 243 182 244 
rect 181 244 182 245 
rect 181 245 182 246 
rect 181 246 182 247 
rect 181 249 182 250 
rect 181 250 182 251 
rect 181 251 182 252 
rect 181 252 182 253 
rect 181 253 182 254 
rect 181 254 182 255 
rect 181 255 182 256 
rect 181 256 182 257 
rect 181 257 182 258 
rect 181 258 182 259 
rect 181 259 182 260 
rect 181 260 182 261 
rect 181 263 182 264 
rect 181 264 182 265 
rect 181 272 182 273 
rect 181 274 182 275 
rect 181 277 182 278 
rect 181 278 182 279 
rect 181 280 182 281 
rect 181 282 182 283 
rect 181 283 182 284 
rect 181 284 182 285 
rect 181 285 182 286 
rect 181 286 182 287 
rect 181 287 182 288 
rect 181 288 182 289 
rect 181 289 182 290 
rect 181 290 182 291 
rect 181 291 182 292 
rect 181 293 182 294 
rect 181 298 182 299 
rect 181 299 182 300 
rect 181 305 182 306 
rect 181 307 182 308 
rect 181 308 182 309 
rect 181 310 182 311 
rect 181 312 182 313 
rect 182 1 183 2 
rect 182 3 183 4 
rect 182 8 183 9 
rect 182 15 183 16 
rect 182 17 183 18 
rect 182 21 183 22 
rect 182 23 183 24 
rect 182 32 183 33 
rect 182 36 183 37 
rect 182 38 183 39 
rect 182 43 183 44 
rect 182 50 183 51 
rect 182 53 183 54 
rect 182 54 183 55 
rect 182 69 183 70 
rect 182 71 183 72 
rect 182 83 183 84 
rect 182 85 183 86 
rect 182 87 183 88 
rect 182 97 183 98 
rect 182 110 183 111 
rect 182 115 183 116 
rect 182 118 183 119 
rect 182 142 183 143 
rect 182 145 183 146 
rect 182 147 183 148 
rect 182 152 183 153 
rect 182 153 183 154 
rect 182 154 183 155 
rect 182 155 183 156 
rect 182 161 183 162 
rect 182 165 183 166 
rect 182 168 183 169 
rect 182 177 183 178 
rect 182 206 183 207 
rect 182 222 183 223 
rect 182 225 183 226 
rect 182 229 183 230 
rect 182 232 183 233 
rect 182 235 183 236 
rect 182 241 183 242 
rect 182 260 183 261 
rect 182 264 183 265 
rect 182 272 183 273 
rect 182 274 183 275 
rect 182 277 183 278 
rect 182 279 183 280 
rect 182 280 183 281 
rect 182 291 183 292 
rect 182 293 183 294 
rect 182 299 183 300 
rect 182 305 183 306 
rect 182 307 183 308 
rect 182 309 183 310 
rect 182 310 183 311 
rect 182 312 183 313 
rect 183 1 184 2 
rect 183 3 184 4 
rect 183 8 184 9 
rect 183 15 184 16 
rect 183 17 184 18 
rect 183 21 184 22 
rect 183 23 184 24 
rect 183 32 184 33 
rect 183 33 184 34 
rect 183 34 184 35 
rect 183 36 184 37 
rect 183 38 184 39 
rect 183 43 184 44 
rect 183 50 184 51 
rect 183 54 184 55 
rect 183 55 184 56 
rect 183 56 184 57 
rect 183 57 184 58 
rect 183 58 184 59 
rect 183 59 184 60 
rect 183 60 184 61 
rect 183 61 184 62 
rect 183 62 184 63 
rect 183 63 184 64 
rect 183 64 184 65 
rect 183 65 184 66 
rect 183 66 184 67 
rect 183 69 184 70 
rect 183 71 184 72 
rect 183 87 184 88 
rect 183 97 184 98 
rect 183 110 184 111 
rect 183 115 184 116 
rect 183 118 184 119 
rect 183 142 184 143 
rect 183 145 184 146 
rect 183 147 184 148 
rect 183 151 184 152 
rect 183 152 184 153 
rect 183 161 184 162 
rect 183 163 184 164 
rect 183 165 184 166 
rect 183 168 184 169 
rect 183 177 184 178 
rect 183 206 184 207 
rect 183 222 184 223 
rect 183 225 184 226 
rect 183 229 184 230 
rect 183 232 184 233 
rect 183 241 184 242 
rect 183 243 184 244 
rect 183 244 184 245 
rect 183 245 184 246 
rect 183 246 184 247 
rect 183 247 184 248 
rect 183 248 184 249 
rect 183 249 184 250 
rect 183 250 184 251 
rect 183 251 184 252 
rect 183 252 184 253 
rect 183 253 184 254 
rect 183 254 184 255 
rect 183 255 184 256 
rect 183 256 184 257 
rect 183 257 184 258 
rect 183 258 184 259 
rect 183 260 184 261 
rect 183 262 184 263 
rect 183 264 184 265 
rect 183 272 184 273 
rect 183 277 184 278 
rect 183 279 184 280 
rect 183 291 184 292 
rect 183 293 184 294 
rect 183 299 184 300 
rect 183 305 184 306 
rect 183 307 184 308 
rect 183 309 184 310 
rect 183 311 184 312 
rect 183 312 184 313 
rect 184 1 185 2 
rect 184 3 185 4 
rect 184 8 185 9 
rect 184 15 185 16 
rect 184 17 185 18 
rect 184 21 185 22 
rect 184 23 185 24 
rect 184 30 185 31 
rect 184 31 185 32 
rect 184 36 185 37 
rect 184 38 185 39 
rect 184 41 185 42 
rect 184 42 185 43 
rect 184 43 185 44 
rect 184 50 185 51 
rect 184 52 185 53 
rect 184 66 185 67 
rect 184 69 185 70 
rect 184 71 185 72 
rect 184 75 185 76 
rect 184 76 185 77 
rect 184 77 185 78 
rect 184 78 185 79 
rect 184 79 185 80 
rect 184 80 185 81 
rect 184 81 185 82 
rect 184 82 185 83 
rect 184 83 185 84 
rect 184 84 185 85 
rect 184 85 185 86 
rect 184 86 185 87 
rect 184 87 185 88 
rect 184 91 185 92 
rect 184 92 185 93 
rect 184 93 185 94 
rect 184 94 185 95 
rect 184 95 185 96 
rect 184 97 185 98 
rect 184 110 185 111 
rect 184 113 185 114 
rect 184 115 185 116 
rect 184 118 185 119 
rect 184 121 185 122 
rect 184 122 185 123 
rect 184 123 185 124 
rect 184 124 185 125 
rect 184 125 185 126 
rect 184 126 185 127 
rect 184 127 185 128 
rect 184 128 185 129 
rect 184 129 185 130 
rect 184 137 185 138 
rect 184 138 185 139 
rect 184 139 185 140 
rect 184 140 185 141 
rect 184 142 185 143 
rect 184 145 185 146 
rect 184 147 185 148 
rect 184 150 185 151 
rect 184 151 185 152 
rect 184 153 185 154 
rect 184 154 185 155 
rect 184 155 185 156 
rect 184 156 185 157 
rect 184 157 185 158 
rect 184 158 185 159 
rect 184 161 185 162 
rect 184 163 185 164 
rect 184 165 185 166 
rect 184 168 185 169 
rect 184 177 185 178 
rect 184 180 185 181 
rect 184 181 185 182 
rect 184 182 185 183 
rect 184 183 185 184 
rect 184 184 185 185 
rect 184 185 185 186 
rect 184 186 185 187 
rect 184 187 185 188 
rect 184 188 185 189 
rect 184 189 185 190 
rect 184 190 185 191 
rect 184 191 185 192 
rect 184 192 185 193 
rect 184 193 185 194 
rect 184 194 185 195 
rect 184 195 185 196 
rect 184 196 185 197 
rect 184 197 185 198 
rect 184 198 185 199 
rect 184 199 185 200 
rect 184 200 185 201 
rect 184 201 185 202 
rect 184 202 185 203 
rect 184 203 185 204 
rect 184 204 185 205 
rect 184 205 185 206 
rect 184 206 185 207 
rect 184 222 185 223 
rect 184 225 185 226 
rect 184 227 185 228 
rect 184 228 185 229 
rect 184 229 185 230 
rect 184 232 185 233 
rect 184 241 185 242 
rect 184 258 185 259 
rect 184 260 185 261 
rect 184 262 185 263 
rect 184 264 185 265 
rect 184 267 185 268 
rect 184 272 185 273 
rect 184 277 185 278 
rect 184 279 185 280 
rect 184 291 185 292 
rect 184 293 185 294 
rect 184 299 185 300 
rect 184 305 185 306 
rect 184 307 185 308 
rect 184 309 185 310 
rect 184 311 185 312 
rect 185 1 186 2 
rect 185 3 186 4 
rect 185 8 186 9 
rect 185 17 186 18 
rect 185 21 186 22 
rect 185 23 186 24 
rect 185 30 186 31 
rect 185 36 186 37 
rect 185 38 186 39 
rect 185 40 186 41 
rect 185 41 186 42 
rect 185 50 186 51 
rect 185 52 186 53 
rect 185 54 186 55 
rect 185 55 186 56 
rect 185 56 186 57 
rect 185 66 186 67 
rect 185 69 186 70 
rect 185 71 186 72 
rect 185 75 186 76 
rect 185 91 186 92 
rect 185 97 186 98 
rect 185 110 186 111 
rect 185 113 186 114 
rect 185 115 186 116 
rect 185 118 186 119 
rect 185 129 186 130 
rect 185 130 186 131 
rect 185 131 186 132 
rect 185 132 186 133 
rect 185 133 186 134 
rect 185 134 186 135 
rect 185 135 186 136 
rect 185 136 186 137 
rect 185 137 186 138 
rect 185 142 186 143 
rect 185 145 186 146 
rect 185 147 186 148 
rect 185 150 186 151 
rect 185 152 186 153 
rect 185 153 186 154 
rect 185 158 186 159 
rect 185 161 186 162 
rect 185 163 186 164 
rect 185 165 186 166 
rect 185 168 186 169 
rect 185 177 186 178 
rect 185 222 186 223 
rect 185 225 186 226 
rect 185 232 186 233 
rect 185 241 186 242 
rect 185 257 186 258 
rect 185 260 186 261 
rect 185 262 186 263 
rect 185 264 186 265 
rect 185 267 186 268 
rect 185 272 186 273 
rect 185 273 186 274 
rect 185 277 186 278 
rect 185 279 186 280 
rect 185 291 186 292 
rect 185 293 186 294 
rect 185 299 186 300 
rect 185 305 186 306 
rect 185 307 186 308 
rect 185 309 186 310 
rect 185 311 186 312 
rect 186 1 187 2 
rect 186 3 187 4 
rect 186 8 187 9 
rect 186 17 187 18 
rect 186 18 187 19 
rect 186 21 187 22 
rect 186 23 187 24 
rect 186 30 187 31 
rect 186 36 187 37 
rect 186 38 187 39 
rect 186 40 187 41 
rect 186 50 187 51 
rect 186 52 187 53 
rect 186 54 187 55 
rect 186 66 187 67 
rect 186 69 187 70 
rect 186 71 187 72 
rect 186 75 187 76 
rect 186 91 187 92 
rect 186 97 187 98 
rect 186 110 187 111 
rect 186 113 187 114 
rect 186 115 187 116 
rect 186 118 187 119 
rect 186 142 187 143 
rect 186 145 187 146 
rect 186 147 187 148 
rect 186 150 187 151 
rect 186 152 187 153 
rect 186 158 187 159 
rect 186 161 187 162 
rect 186 163 187 164 
rect 186 165 187 166 
rect 186 168 187 169 
rect 186 177 187 178 
rect 186 222 187 223 
rect 186 225 187 226 
rect 186 227 187 228 
rect 186 228 187 229 
rect 186 229 187 230 
rect 186 230 187 231 
rect 186 232 187 233 
rect 186 241 187 242 
rect 186 257 187 258 
rect 186 260 187 261 
rect 186 262 187 263 
rect 186 264 187 265 
rect 186 267 187 268 
rect 186 273 187 274 
rect 186 277 187 278 
rect 186 279 187 280 
rect 186 291 187 292 
rect 186 293 187 294 
rect 186 299 187 300 
rect 186 305 187 306 
rect 186 307 187 308 
rect 186 309 187 310 
rect 186 311 187 312 
rect 187 1 188 2 
rect 187 3 188 4 
rect 187 8 188 9 
rect 187 18 188 19 
rect 187 21 188 22 
rect 187 23 188 24 
rect 187 36 188 37 
rect 187 38 188 39 
rect 187 40 188 41 
rect 187 50 188 51 
rect 187 52 188 53 
rect 187 54 188 55 
rect 187 66 188 67 
rect 187 69 188 70 
rect 187 71 188 72 
rect 187 97 188 98 
rect 187 113 188 114 
rect 187 115 188 116 
rect 187 118 188 119 
rect 187 145 188 146 
rect 187 147 188 148 
rect 187 150 188 151 
rect 187 152 188 153 
rect 187 161 188 162 
rect 187 163 188 164 
rect 187 165 188 166 
rect 187 168 188 169 
rect 187 177 188 178 
rect 187 225 188 226 
rect 187 227 188 228 
rect 187 232 188 233 
rect 187 241 188 242 
rect 187 257 188 258 
rect 187 260 188 261 
rect 187 262 188 263 
rect 187 264 188 265 
rect 187 273 188 274 
rect 187 277 188 278 
rect 187 279 188 280 
rect 187 291 188 292 
rect 187 293 188 294 
rect 187 305 188 306 
rect 187 307 188 308 
rect 187 309 188 310 
rect 187 311 188 312 
rect 188 1 189 2 
rect 188 3 189 4 
rect 188 8 189 9 
rect 188 18 189 19 
rect 188 21 189 22 
rect 188 23 189 24 
rect 188 36 189 37 
rect 188 38 189 39 
rect 188 40 189 41 
rect 188 50 189 51 
rect 188 52 189 53 
rect 188 54 189 55 
rect 188 66 189 67 
rect 188 69 189 70 
rect 188 71 189 72 
rect 188 97 189 98 
rect 188 113 189 114 
rect 188 115 189 116 
rect 188 118 189 119 
rect 188 145 189 146 
rect 188 147 189 148 
rect 188 150 189 151 
rect 188 152 189 153 
rect 188 161 189 162 
rect 188 163 189 164 
rect 188 165 189 166 
rect 188 168 189 169 
rect 188 177 189 178 
rect 188 225 189 226 
rect 188 227 189 228 
rect 188 232 189 233 
rect 188 241 189 242 
rect 188 257 189 258 
rect 188 260 189 261 
rect 188 262 189 263 
rect 188 264 189 265 
rect 188 273 189 274 
rect 188 277 189 278 
rect 188 279 189 280 
rect 188 291 189 292 
rect 188 293 189 294 
rect 188 305 189 306 
rect 188 307 189 308 
rect 188 309 189 310 
rect 188 311 189 312 
rect 189 1 190 2 
rect 189 3 190 4 
rect 189 8 190 9 
rect 189 18 190 19 
rect 189 21 190 22 
rect 189 23 190 24 
rect 189 36 190 37 
rect 189 38 190 39 
rect 189 40 190 41 
rect 189 50 190 51 
rect 189 52 190 53 
rect 189 54 190 55 
rect 189 66 190 67 
rect 189 69 190 70 
rect 189 71 190 72 
rect 189 97 190 98 
rect 189 113 190 114 
rect 189 115 190 116 
rect 189 118 190 119 
rect 189 145 190 146 
rect 189 147 190 148 
rect 189 150 190 151 
rect 189 152 190 153 
rect 189 161 190 162 
rect 189 163 190 164 
rect 189 165 190 166 
rect 189 168 190 169 
rect 189 177 190 178 
rect 189 225 190 226 
rect 189 227 190 228 
rect 189 232 190 233 
rect 189 241 190 242 
rect 189 257 190 258 
rect 189 260 190 261 
rect 189 262 190 263 
rect 189 264 190 265 
rect 189 273 190 274 
rect 189 277 190 278 
rect 189 279 190 280 
rect 189 291 190 292 
rect 189 293 190 294 
rect 189 305 190 306 
rect 189 307 190 308 
rect 189 309 190 310 
rect 189 311 190 312 
rect 190 1 191 2 
rect 190 3 191 4 
rect 190 8 191 9 
rect 190 18 191 19 
rect 190 21 191 22 
rect 190 23 191 24 
rect 190 36 191 37 
rect 190 38 191 39 
rect 190 40 191 41 
rect 190 50 191 51 
rect 190 52 191 53 
rect 190 54 191 55 
rect 190 66 191 67 
rect 190 69 191 70 
rect 190 71 191 72 
rect 190 97 191 98 
rect 190 113 191 114 
rect 190 115 191 116 
rect 190 118 191 119 
rect 190 145 191 146 
rect 190 147 191 148 
rect 190 150 191 151 
rect 190 152 191 153 
rect 190 161 191 162 
rect 190 163 191 164 
rect 190 165 191 166 
rect 190 168 191 169 
rect 190 177 191 178 
rect 190 225 191 226 
rect 190 227 191 228 
rect 190 232 191 233 
rect 190 241 191 242 
rect 190 257 191 258 
rect 190 260 191 261 
rect 190 262 191 263 
rect 190 264 191 265 
rect 190 273 191 274 
rect 190 277 191 278 
rect 190 279 191 280 
rect 190 291 191 292 
rect 190 293 191 294 
rect 190 305 191 306 
rect 190 307 191 308 
rect 190 309 191 310 
rect 190 311 191 312 
rect 191 1 192 2 
rect 191 3 192 4 
rect 191 8 192 9 
rect 191 18 192 19 
rect 191 19 192 20 
rect 191 21 192 22 
rect 191 23 192 24 
rect 191 27 192 28 
rect 191 36 192 37 
rect 191 38 192 39 
rect 191 40 192 41 
rect 191 46 192 47 
rect 191 50 192 51 
rect 191 52 192 53 
rect 191 54 192 55 
rect 191 62 192 63 
rect 191 66 192 67 
rect 191 69 192 70 
rect 191 71 192 72 
rect 191 75 192 76 
rect 191 78 192 79 
rect 191 94 192 95 
rect 191 97 192 98 
rect 191 113 192 114 
rect 191 115 192 116 
rect 191 118 192 119 
rect 191 145 192 146 
rect 191 147 192 148 
rect 191 150 192 151 
rect 191 152 192 153 
rect 191 161 192 162 
rect 191 163 192 164 
rect 191 165 192 166 
rect 191 168 192 169 
rect 191 177 192 178 
rect 191 225 192 226 
rect 191 227 192 228 
rect 191 232 192 233 
rect 191 241 192 242 
rect 191 257 192 258 
rect 191 260 192 261 
rect 191 262 192 263 
rect 191 264 192 265 
rect 191 273 192 274 
rect 191 277 192 278 
rect 191 279 192 280 
rect 191 291 192 292 
rect 191 293 192 294 
rect 191 299 192 300 
rect 191 305 192 306 
rect 191 307 192 308 
rect 191 309 192 310 
rect 191 311 192 312 
rect 192 1 193 2 
rect 192 3 193 4 
rect 192 8 193 9 
rect 192 19 193 20 
rect 192 20 193 21 
rect 192 23 193 24 
rect 192 27 193 28 
rect 192 32 193 33 
rect 192 33 193 34 
rect 192 36 193 37 
rect 192 38 193 39 
rect 192 40 193 41 
rect 192 46 193 47 
rect 192 50 193 51 
rect 192 52 193 53 
rect 192 54 193 55 
rect 192 62 193 63 
rect 192 66 193 67 
rect 192 69 193 70 
rect 192 71 193 72 
rect 192 75 193 76 
rect 192 78 193 79 
rect 192 94 193 95 
rect 192 97 193 98 
rect 192 112 193 113 
rect 192 113 193 114 
rect 192 115 193 116 
rect 192 118 193 119 
rect 192 144 193 145 
rect 192 145 193 146 
rect 192 147 193 148 
rect 192 150 193 151 
rect 192 152 193 153 
rect 192 153 193 154 
rect 192 161 193 162 
rect 192 165 193 166 
rect 192 168 193 169 
rect 192 169 193 170 
rect 192 176 193 177 
rect 192 177 193 178 
rect 192 224 193 225 
rect 192 225 193 226 
rect 192 227 193 228 
rect 192 232 193 233 
rect 192 240 193 241 
rect 192 241 193 242 
rect 192 256 193 257 
rect 192 257 193 258 
rect 192 260 193 261 
rect 192 262 193 263 
rect 192 264 193 265 
rect 192 265 193 266 
rect 192 273 193 274 
rect 192 299 193 300 
rect 192 305 193 306 
rect 192 307 193 308 
rect 192 309 193 310 
rect 192 311 193 312 
rect 193 1 194 2 
rect 193 3 194 4 
rect 193 8 194 9 
rect 193 17 194 18 
rect 193 18 194 19 
rect 193 20 194 21 
rect 193 21 194 22 
rect 193 23 194 24 
rect 193 25 194 26 
rect 193 26 194 27 
rect 193 27 194 28 
rect 193 32 194 33 
rect 193 36 194 37 
rect 193 40 194 41 
rect 193 43 194 44 
rect 193 44 194 45 
rect 193 45 194 46 
rect 193 46 194 47 
rect 193 50 194 51 
rect 193 52 194 53 
rect 193 54 194 55 
rect 193 62 194 63 
rect 193 63 194 64 
rect 193 64 194 65 
rect 193 66 194 67 
rect 193 71 194 72 
rect 193 73 194 74 
rect 193 75 194 76 
rect 193 76 194 77 
rect 193 78 194 79 
rect 193 79 194 80 
rect 193 80 194 81 
rect 193 81 194 82 
rect 193 82 194 83 
rect 193 83 194 84 
rect 193 84 194 85 
rect 193 85 194 86 
rect 193 86 194 87 
rect 193 87 194 88 
rect 193 88 194 89 
rect 193 89 194 90 
rect 193 90 194 91 
rect 193 91 194 92 
rect 193 94 194 95 
rect 193 97 194 98 
rect 193 99 194 100 
rect 193 100 194 101 
rect 193 101 194 102 
rect 193 102 194 103 
rect 193 103 194 104 
rect 193 104 194 105 
rect 193 105 194 106 
rect 193 106 194 107 
rect 193 107 194 108 
rect 193 108 194 109 
rect 193 109 194 110 
rect 193 110 194 111 
rect 193 111 194 112 
rect 193 112 194 113 
rect 193 115 194 116 
rect 193 118 194 119 
rect 193 120 194 121 
rect 193 121 194 122 
rect 193 122 194 123 
rect 193 123 194 124 
rect 193 124 194 125 
rect 193 125 194 126 
rect 193 126 194 127 
rect 193 127 194 128 
rect 193 128 194 129 
rect 193 129 194 130 
rect 193 130 194 131 
rect 193 131 194 132 
rect 193 132 194 133 
rect 193 133 194 134 
rect 193 134 194 135 
rect 193 135 194 136 
rect 193 136 194 137 
rect 193 137 194 138 
rect 193 138 194 139 
rect 193 139 194 140 
rect 193 140 194 141 
rect 193 141 194 142 
rect 193 142 194 143 
rect 193 143 194 144 
rect 193 144 194 145 
rect 193 147 194 148 
rect 193 150 194 151 
rect 193 151 194 152 
rect 193 153 194 154 
rect 193 161 194 162 
rect 193 165 194 166 
rect 193 169 194 170 
rect 193 170 194 171 
rect 193 171 194 172 
rect 193 173 194 174 
rect 193 174 194 175 
rect 193 175 194 176 
rect 193 176 194 177 
rect 193 182 194 183 
rect 193 183 194 184 
rect 193 184 194 185 
rect 193 185 194 186 
rect 193 186 194 187 
rect 193 187 194 188 
rect 193 188 194 189 
rect 193 189 194 190 
rect 193 190 194 191 
rect 193 191 194 192 
rect 193 192 194 193 
rect 193 193 194 194 
rect 193 194 194 195 
rect 193 195 194 196 
rect 193 196 194 197 
rect 193 197 194 198 
rect 193 198 194 199 
rect 193 199 194 200 
rect 193 200 194 201 
rect 193 201 194 202 
rect 193 202 194 203 
rect 193 203 194 204 
rect 193 204 194 205 
rect 193 205 194 206 
rect 193 206 194 207 
rect 193 207 194 208 
rect 193 208 194 209 
rect 193 209 194 210 
rect 193 210 194 211 
rect 193 211 194 212 
rect 193 212 194 213 
rect 193 213 194 214 
rect 193 214 194 215 
rect 193 215 194 216 
rect 193 216 194 217 
rect 193 217 194 218 
rect 193 218 194 219 
rect 193 219 194 220 
rect 193 220 194 221 
rect 193 221 194 222 
rect 193 222 194 223 
rect 193 223 194 224 
rect 193 224 194 225 
rect 193 226 194 227 
rect 193 227 194 228 
rect 193 232 194 233 
rect 193 234 194 235 
rect 193 235 194 236 
rect 193 236 194 237 
rect 193 237 194 238 
rect 193 238 194 239 
rect 193 239 194 240 
rect 193 240 194 241 
rect 193 242 194 243 
rect 193 243 194 244 
rect 193 244 194 245 
rect 193 245 194 246 
rect 193 246 194 247 
rect 193 247 194 248 
rect 193 248 194 249 
rect 193 249 194 250 
rect 193 250 194 251 
rect 193 251 194 252 
rect 193 252 194 253 
rect 193 253 194 254 
rect 193 254 194 255 
rect 193 255 194 256 
rect 193 256 194 257 
rect 193 260 194 261 
rect 193 265 194 266 
rect 193 266 194 267 
rect 193 267 194 268 
rect 193 268 194 269 
rect 193 269 194 270 
rect 193 270 194 271 
rect 193 271 194 272 
rect 193 273 194 274 
rect 193 276 194 277 
rect 193 277 194 278 
rect 193 278 194 279 
rect 193 279 194 280 
rect 193 280 194 281 
rect 193 281 194 282 
rect 193 282 194 283 
rect 193 283 194 284 
rect 193 284 194 285 
rect 193 285 194 286 
rect 193 286 194 287 
rect 193 287 194 288 
rect 193 288 194 289 
rect 193 289 194 290 
rect 193 290 194 291 
rect 193 291 194 292 
rect 193 292 194 293 
rect 193 293 194 294 
rect 193 294 194 295 
rect 193 295 194 296 
rect 193 296 194 297 
rect 193 297 194 298 
rect 193 298 194 299 
rect 193 299 194 300 
rect 193 305 194 306 
rect 193 307 194 308 
rect 193 309 194 310 
rect 193 311 194 312 
rect 194 1 195 2 
rect 194 3 195 4 
rect 194 8 195 9 
rect 194 18 195 19 
rect 194 21 195 22 
rect 194 23 195 24 
rect 194 32 195 33 
rect 194 36 195 37 
rect 194 40 195 41 
rect 194 50 195 51 
rect 194 52 195 53 
rect 194 54 195 55 
rect 194 66 195 67 
rect 194 68 195 69 
rect 194 71 195 72 
rect 194 73 195 74 
rect 194 76 195 77 
rect 194 77 195 78 
rect 194 94 195 95 
rect 194 97 195 98 
rect 194 99 195 100 
rect 194 115 195 116 
rect 194 118 195 119 
rect 194 147 195 148 
rect 194 153 195 154 
rect 194 161 195 162 
rect 194 163 195 164 
rect 194 165 195 166 
rect 194 171 195 172 
rect 194 182 195 183 
rect 194 225 195 226 
rect 194 226 195 227 
rect 194 228 195 229 
rect 194 230 195 231 
rect 194 232 195 233 
rect 194 241 195 242 
rect 194 242 195 243 
rect 194 260 195 261 
rect 194 273 195 274 
rect 194 303 195 304 
rect 194 305 195 306 
rect 194 308 195 309 
rect 194 309 195 310 
rect 194 311 195 312 
rect 195 1 196 2 
rect 195 3 196 4 
rect 195 8 196 9 
rect 195 18 196 19 
rect 195 21 196 22 
rect 195 23 196 24 
rect 195 32 196 33 
rect 195 36 196 37 
rect 195 40 196 41 
rect 195 50 196 51 
rect 195 52 196 53 
rect 195 54 196 55 
rect 195 66 196 67 
rect 195 68 196 69 
rect 195 71 196 72 
rect 195 73 196 74 
rect 195 77 196 78 
rect 195 78 196 79 
rect 195 79 196 80 
rect 195 80 196 81 
rect 195 81 196 82 
rect 195 82 196 83 
rect 195 83 196 84 
rect 195 84 196 85 
rect 195 85 196 86 
rect 195 86 196 87 
rect 195 87 196 88 
rect 195 88 196 89 
rect 195 89 196 90 
rect 195 90 196 91 
rect 195 91 196 92 
rect 195 92 196 93 
rect 195 94 196 95 
rect 195 97 196 98 
rect 195 115 196 116 
rect 195 118 196 119 
rect 195 147 196 148 
rect 195 153 196 154 
rect 195 161 196 162 
rect 195 163 196 164 
rect 195 165 196 166 
rect 195 171 196 172 
rect 195 182 196 183 
rect 195 185 196 186 
rect 195 186 196 187 
rect 195 192 196 193 
rect 195 193 196 194 
rect 195 194 196 195 
rect 195 195 196 196 
rect 195 196 196 197 
rect 195 197 196 198 
rect 195 198 196 199 
rect 195 199 196 200 
rect 195 200 196 201 
rect 195 201 196 202 
rect 195 202 196 203 
rect 195 203 196 204 
rect 195 204 196 205 
rect 195 205 196 206 
rect 195 206 196 207 
rect 195 207 196 208 
rect 195 208 196 209 
rect 195 209 196 210 
rect 195 210 196 211 
rect 195 211 196 212 
rect 195 212 196 213 
rect 195 213 196 214 
rect 195 214 196 215 
rect 195 215 196 216 
rect 195 216 196 217 
rect 195 217 196 218 
rect 195 218 196 219 
rect 195 219 196 220 
rect 195 220 196 221 
rect 195 221 196 222 
rect 195 222 196 223 
rect 195 223 196 224 
rect 195 224 196 225 
rect 195 225 196 226 
rect 195 228 196 229 
rect 195 230 196 231 
rect 195 232 196 233 
rect 195 234 196 235 
rect 195 235 196 236 
rect 195 236 196 237 
rect 195 237 196 238 
rect 195 238 196 239 
rect 195 239 196 240 
rect 195 240 196 241 
rect 195 241 196 242 
rect 195 264 196 265 
rect 195 265 196 266 
rect 195 266 196 267 
rect 195 267 196 268 
rect 195 268 196 269 
rect 195 269 196 270 
rect 195 270 196 271 
rect 195 273 196 274 
rect 195 275 196 276 
rect 195 276 196 277 
rect 195 277 196 278 
rect 195 278 196 279 
rect 195 279 196 280 
rect 195 280 196 281 
rect 195 281 196 282 
rect 195 282 196 283 
rect 195 283 196 284 
rect 195 284 196 285 
rect 195 285 196 286 
rect 195 286 196 287 
rect 195 287 196 288 
rect 195 288 196 289 
rect 195 293 196 294 
rect 195 294 196 295 
rect 195 295 196 296 
rect 195 296 196 297 
rect 195 297 196 298 
rect 195 298 196 299 
rect 195 299 196 300 
rect 195 300 196 301 
rect 195 301 196 302 
rect 195 302 196 303 
rect 195 303 196 304 
rect 195 305 196 306 
rect 195 308 196 309 
rect 195 310 196 311 
rect 195 311 196 312 
rect 196 1 197 2 
rect 196 3 197 4 
rect 196 8 197 9 
rect 196 18 197 19 
rect 196 21 197 22 
rect 196 23 197 24 
rect 196 32 197 33 
rect 196 36 197 37 
rect 196 40 197 41 
rect 196 50 197 51 
rect 196 52 197 53 
rect 196 54 197 55 
rect 196 66 197 67 
rect 196 68 197 69 
rect 196 71 197 72 
rect 196 73 197 74 
rect 196 94 197 95 
rect 196 97 197 98 
rect 196 115 197 116 
rect 196 118 197 119 
rect 196 147 197 148 
rect 196 153 197 154 
rect 196 161 197 162 
rect 196 163 197 164 
rect 196 165 197 166 
rect 196 171 197 172 
rect 196 182 197 183 
rect 196 186 197 187 
rect 196 187 197 188 
rect 196 188 197 189 
rect 196 189 197 190 
rect 196 190 197 191 
rect 196 191 197 192 
rect 196 192 197 193 
rect 196 228 197 229 
rect 196 230 197 231 
rect 196 232 197 233 
rect 196 234 197 235 
rect 196 242 197 243 
rect 196 243 197 244 
rect 196 244 197 245 
rect 196 245 197 246 
rect 196 246 197 247 
rect 196 247 197 248 
rect 196 248 197 249 
rect 196 249 197 250 
rect 196 250 197 251 
rect 196 251 197 252 
rect 196 252 197 253 
rect 196 253 197 254 
rect 196 254 197 255 
rect 196 255 197 256 
rect 196 256 197 257 
rect 196 257 197 258 
rect 196 258 197 259 
rect 196 259 197 260 
rect 196 260 197 261 
rect 196 261 197 262 
rect 196 262 197 263 
rect 196 264 197 265 
rect 196 273 197 274 
rect 196 275 197 276 
rect 196 293 197 294 
rect 196 305 197 306 
rect 196 308 197 309 
rect 196 310 197 311 
rect 197 1 198 2 
rect 197 3 198 4 
rect 197 8 198 9 
rect 197 18 198 19 
rect 197 21 198 22 
rect 197 23 198 24 
rect 197 32 198 33 
rect 197 36 198 37 
rect 197 40 198 41 
rect 197 50 198 51 
rect 197 52 198 53 
rect 197 54 198 55 
rect 197 66 198 67 
rect 197 68 198 69 
rect 197 71 198 72 
rect 197 73 198 74 
rect 197 82 198 83 
rect 197 94 198 95 
rect 197 97 198 98 
rect 197 100 198 101 
rect 197 115 198 116 
rect 197 118 198 119 
rect 197 147 198 148 
rect 197 153 198 154 
rect 197 161 198 162 
rect 197 163 198 164 
rect 197 165 198 166 
rect 197 171 198 172 
rect 197 182 198 183 
rect 197 193 198 194 
rect 197 194 198 195 
rect 197 195 198 196 
rect 197 196 198 197 
rect 197 197 198 198 
rect 197 198 198 199 
rect 197 199 198 200 
rect 197 200 198 201 
rect 197 201 198 202 
rect 197 202 198 203 
rect 197 203 198 204 
rect 197 204 198 205 
rect 197 205 198 206 
rect 197 206 198 207 
rect 197 207 198 208 
rect 197 208 198 209 
rect 197 209 198 210 
rect 197 210 198 211 
rect 197 211 198 212 
rect 197 212 198 213 
rect 197 213 198 214 
rect 197 214 198 215 
rect 197 215 198 216 
rect 197 216 198 217 
rect 197 217 198 218 
rect 197 218 198 219 
rect 197 219 198 220 
rect 197 220 198 221 
rect 197 221 198 222 
rect 197 222 198 223 
rect 197 223 198 224 
rect 197 224 198 225 
rect 197 225 198 226 
rect 197 226 198 227 
rect 197 228 198 229 
rect 197 230 198 231 
rect 197 232 198 233 
rect 197 242 198 243 
rect 197 264 198 265 
rect 197 273 198 274 
rect 197 275 198 276 
rect 197 293 198 294 
rect 197 305 198 306 
rect 197 308 198 309 
rect 197 310 198 311 
rect 198 1 199 2 
rect 198 3 199 4 
rect 198 8 199 9 
rect 198 18 199 19 
rect 198 21 199 22 
rect 198 23 199 24 
rect 198 32 199 33 
rect 198 36 199 37 
rect 198 40 199 41 
rect 198 50 199 51 
rect 198 52 199 53 
rect 198 54 199 55 
rect 198 66 199 67 
rect 198 68 199 69 
rect 198 71 199 72 
rect 198 73 199 74 
rect 198 82 199 83 
rect 198 94 199 95 
rect 198 97 199 98 
rect 198 100 199 101 
rect 198 103 199 104 
rect 198 104 199 105 
rect 198 105 199 106 
rect 198 106 199 107 
rect 198 107 199 108 
rect 198 108 199 109 
rect 198 109 199 110 
rect 198 110 199 111 
rect 198 111 199 112 
rect 198 112 199 113 
rect 198 113 199 114 
rect 198 115 199 116 
rect 198 118 199 119 
rect 198 147 199 148 
rect 198 153 199 154 
rect 198 161 199 162 
rect 198 163 199 164 
rect 198 165 199 166 
rect 198 171 199 172 
rect 198 182 199 183 
rect 198 184 199 185 
rect 198 185 199 186 
rect 198 186 199 187 
rect 198 187 199 188 
rect 198 188 199 189 
rect 198 189 199 190 
rect 198 190 199 191 
rect 198 191 199 192 
rect 198 192 199 193 
rect 198 193 199 194 
rect 198 228 199 229 
rect 198 230 199 231 
rect 198 232 199 233 
rect 198 242 199 243 
rect 198 247 199 248 
rect 198 259 199 260 
rect 198 264 199 265 
rect 198 273 199 274 
rect 198 275 199 276 
rect 198 293 199 294 
rect 198 305 199 306 
rect 198 308 199 309 
rect 198 310 199 311 
rect 199 1 200 2 
rect 199 3 200 4 
rect 199 8 200 9 
rect 199 18 200 19 
rect 199 21 200 22 
rect 199 23 200 24 
rect 199 32 200 33 
rect 199 36 200 37 
rect 199 40 200 41 
rect 199 50 200 51 
rect 199 52 200 53 
rect 199 54 200 55 
rect 199 66 200 67 
rect 199 68 200 69 
rect 199 71 200 72 
rect 199 73 200 74 
rect 199 82 200 83 
rect 199 94 200 95 
rect 199 97 200 98 
rect 199 100 200 101 
rect 199 103 200 104 
rect 199 113 200 114 
rect 199 115 200 116 
rect 199 118 200 119 
rect 199 147 200 148 
rect 199 153 200 154 
rect 199 163 200 164 
rect 199 165 200 166 
rect 199 171 200 172 
rect 199 182 200 183 
rect 199 184 200 185 
rect 199 227 200 228 
rect 199 228 200 229 
rect 199 230 200 231 
rect 199 232 200 233 
rect 199 242 200 243 
rect 199 244 200 245 
rect 199 245 200 246 
rect 199 247 200 248 
rect 199 259 200 260 
rect 199 264 200 265 
rect 199 273 200 274 
rect 199 275 200 276 
rect 199 293 200 294 
rect 199 305 200 306 
rect 199 308 200 309 
rect 199 310 200 311 
rect 200 1 201 2 
rect 200 3 201 4 
rect 200 8 201 9 
rect 200 18 201 19 
rect 200 21 201 22 
rect 200 23 201 24 
rect 200 27 201 28 
rect 200 28 201 29 
rect 200 29 201 30 
rect 200 30 201 31 
rect 200 31 201 32 
rect 200 32 201 33 
rect 200 36 201 37 
rect 200 40 201 41 
rect 200 50 201 51 
rect 200 52 201 53 
rect 200 54 201 55 
rect 200 66 201 67 
rect 200 68 201 69 
rect 200 71 201 72 
rect 200 73 201 74 
rect 200 74 201 75 
rect 200 75 201 76 
rect 200 82 201 83 
rect 200 89 201 90 
rect 200 90 201 91 
rect 200 91 201 92 
rect 200 92 201 93 
rect 200 93 201 94 
rect 200 94 201 95 
rect 200 97 201 98 
rect 200 100 201 101 
rect 200 113 201 114 
rect 200 115 201 116 
rect 200 118 201 119 
rect 200 123 201 124 
rect 200 124 201 125 
rect 200 125 201 126 
rect 200 126 201 127 
rect 200 127 201 128 
rect 200 128 201 129 
rect 200 129 201 130 
rect 200 130 201 131 
rect 200 131 201 132 
rect 200 132 201 133 
rect 200 133 201 134 
rect 200 134 201 135 
rect 200 135 201 136 
rect 200 136 201 137 
rect 200 137 201 138 
rect 200 138 201 139 
rect 200 139 201 140 
rect 200 140 201 141 
rect 200 141 201 142 
rect 200 142 201 143 
rect 200 143 201 144 
rect 200 144 201 145 
rect 200 145 201 146 
rect 200 146 201 147 
rect 200 147 201 148 
rect 200 153 201 154 
rect 200 155 201 156 
rect 200 156 201 157 
rect 200 157 201 158 
rect 200 158 201 159 
rect 200 159 201 160 
rect 200 160 201 161 
rect 200 161 201 162 
rect 200 162 201 163 
rect 200 163 201 164 
rect 200 165 201 166 
rect 200 171 201 172 
rect 200 182 201 183 
rect 200 184 201 185 
rect 200 219 201 220 
rect 200 220 201 221 
rect 200 221 201 222 
rect 200 222 201 223 
rect 200 223 201 224 
rect 200 224 201 225 
rect 200 225 201 226 
rect 200 226 201 227 
rect 200 227 201 228 
rect 200 229 201 230 
rect 200 230 201 231 
rect 200 232 201 233 
rect 200 242 201 243 
rect 200 245 201 246 
rect 200 247 201 248 
rect 200 259 201 260 
rect 200 264 201 265 
rect 200 273 201 274 
rect 200 275 201 276 
rect 200 293 201 294 
rect 200 297 201 298 
rect 200 298 201 299 
rect 200 299 201 300 
rect 200 300 201 301 
rect 200 301 201 302 
rect 200 302 201 303 
rect 200 305 201 306 
rect 200 308 201 309 
rect 200 310 201 311 
rect 201 1 202 2 
rect 201 3 202 4 
rect 201 8 202 9 
rect 201 18 202 19 
rect 201 21 202 22 
rect 201 23 202 24 
rect 201 27 202 28 
rect 201 36 202 37 
rect 201 40 202 41 
rect 201 50 202 51 
rect 201 52 202 53 
rect 201 54 202 55 
rect 201 66 202 67 
rect 201 68 202 69 
rect 201 71 202 72 
rect 201 75 202 76 
rect 201 82 202 83 
rect 201 88 202 89 
rect 201 89 202 90 
rect 201 97 202 98 
rect 201 100 202 101 
rect 201 113 202 114 
rect 201 115 202 116 
rect 201 118 202 119 
rect 201 123 202 124 
rect 201 152 202 153 
rect 201 153 202 154 
rect 201 155 202 156 
rect 201 165 202 166 
rect 201 171 202 172 
rect 201 182 202 183 
rect 201 184 202 185 
rect 201 219 202 220 
rect 201 229 202 230 
rect 201 232 202 233 
rect 201 242 202 243 
rect 201 245 202 246 
rect 201 247 202 248 
rect 201 259 202 260 
rect 201 262 202 263 
rect 201 263 202 264 
rect 201 264 202 265 
rect 201 273 202 274 
rect 201 275 202 276 
rect 201 293 202 294 
rect 201 296 202 297 
rect 201 297 202 298 
rect 201 302 202 303 
rect 201 305 202 306 
rect 201 308 202 309 
rect 201 310 202 311 
rect 202 1 203 2 
rect 202 3 203 4 
rect 202 8 203 9 
rect 202 18 203 19 
rect 202 21 203 22 
rect 202 23 203 24 
rect 202 27 203 28 
rect 202 36 203 37 
rect 202 40 203 41 
rect 202 50 203 51 
rect 202 52 203 53 
rect 202 54 203 55 
rect 202 66 203 67 
rect 202 68 203 69 
rect 202 71 203 72 
rect 202 75 203 76 
rect 202 82 203 83 
rect 202 88 203 89 
rect 202 97 203 98 
rect 202 100 203 101 
rect 202 113 203 114 
rect 202 115 203 116 
rect 202 118 203 119 
rect 202 123 203 124 
rect 202 152 203 153 
rect 202 155 203 156 
rect 202 165 203 166 
rect 202 171 203 172 
rect 202 182 203 183 
rect 202 184 203 185 
rect 202 219 203 220 
rect 202 229 203 230 
rect 202 232 203 233 
rect 202 242 203 243 
rect 202 245 203 246 
rect 202 247 203 248 
rect 202 259 203 260 
rect 202 262 203 263 
rect 202 273 203 274 
rect 202 275 203 276 
rect 202 289 203 290 
rect 202 290 203 291 
rect 202 291 203 292 
rect 202 292 203 293 
rect 202 293 203 294 
rect 202 295 203 296 
rect 202 296 203 297 
rect 202 302 203 303 
rect 202 305 203 306 
rect 202 308 203 309 
rect 202 310 203 311 
rect 203 1 204 2 
rect 203 3 204 4 
rect 203 8 204 9 
rect 203 18 204 19 
rect 203 21 204 22 
rect 203 23 204 24 
rect 203 36 204 37 
rect 203 40 204 41 
rect 203 50 204 51 
rect 203 52 204 53 
rect 203 54 204 55 
rect 203 66 204 67 
rect 203 68 204 69 
rect 203 71 204 72 
rect 203 82 204 83 
rect 203 88 204 89 
rect 203 97 204 98 
rect 203 100 204 101 
rect 203 113 204 114 
rect 203 115 204 116 
rect 203 118 204 119 
rect 203 152 204 153 
rect 203 165 204 166 
rect 203 182 204 183 
rect 203 184 204 185 
rect 203 229 204 230 
rect 203 232 204 233 
rect 203 242 204 243 
rect 203 245 204 246 
rect 203 247 204 248 
rect 203 259 204 260 
rect 203 262 204 263 
rect 203 273 204 274 
rect 203 275 204 276 
rect 203 289 204 290 
rect 203 294 204 295 
rect 203 295 204 296 
rect 203 305 204 306 
rect 203 308 204 309 
rect 203 310 204 311 
rect 204 1 205 2 
rect 204 3 205 4 
rect 204 8 205 9 
rect 204 18 205 19 
rect 204 21 205 22 
rect 204 23 205 24 
rect 204 36 205 37 
rect 204 40 205 41 
rect 204 50 205 51 
rect 204 52 205 53 
rect 204 54 205 55 
rect 204 66 205 67 
rect 204 68 205 69 
rect 204 71 205 72 
rect 204 82 205 83 
rect 204 88 205 89 
rect 204 97 205 98 
rect 204 100 205 101 
rect 204 113 205 114 
rect 204 115 205 116 
rect 204 118 205 119 
rect 204 152 205 153 
rect 204 165 205 166 
rect 204 182 205 183 
rect 204 184 205 185 
rect 204 229 205 230 
rect 204 232 205 233 
rect 204 242 205 243 
rect 204 245 205 246 
rect 204 247 205 248 
rect 204 259 205 260 
rect 204 262 205 263 
rect 204 264 205 265 
rect 204 273 205 274 
rect 204 275 205 276 
rect 204 289 205 290 
rect 204 291 205 292 
rect 204 292 205 293 
rect 204 293 205 294 
rect 204 294 205 295 
rect 204 305 205 306 
rect 204 308 205 309 
rect 204 310 205 311 
rect 205 1 206 2 
rect 205 3 206 4 
rect 205 8 206 9 
rect 205 18 206 19 
rect 205 21 206 22 
rect 205 23 206 24 
rect 205 36 206 37 
rect 205 40 206 41 
rect 205 50 206 51 
rect 205 52 206 53 
rect 205 54 206 55 
rect 205 66 206 67 
rect 205 68 206 69 
rect 205 71 206 72 
rect 205 82 206 83 
rect 205 88 206 89 
rect 205 97 206 98 
rect 205 100 206 101 
rect 205 113 206 114 
rect 205 115 206 116 
rect 205 118 206 119 
rect 205 152 206 153 
rect 205 165 206 166 
rect 205 182 206 183 
rect 205 184 206 185 
rect 205 229 206 230 
rect 205 232 206 233 
rect 205 242 206 243 
rect 205 245 206 246 
rect 205 247 206 248 
rect 205 257 206 258 
rect 205 258 206 259 
rect 205 259 206 260 
rect 205 262 206 263 
rect 205 264 206 265 
rect 205 273 206 274 
rect 205 275 206 276 
rect 205 289 206 290 
rect 205 291 206 292 
rect 205 305 206 306 
rect 205 308 206 309 
rect 205 310 206 311 
rect 206 1 207 2 
rect 206 3 207 4 
rect 206 8 207 9 
rect 206 18 207 19 
rect 206 21 207 22 
rect 206 23 207 24 
rect 206 36 207 37 
rect 206 40 207 41 
rect 206 50 207 51 
rect 206 52 207 53 
rect 206 54 207 55 
rect 206 66 207 67 
rect 206 68 207 69 
rect 206 71 207 72 
rect 206 82 207 83 
rect 206 87 207 88 
rect 206 88 207 89 
rect 206 97 207 98 
rect 206 100 207 101 
rect 206 113 207 114 
rect 206 115 207 116 
rect 206 118 207 119 
rect 206 145 207 146 
rect 206 146 207 147 
rect 206 147 207 148 
rect 206 148 207 149 
rect 206 149 207 150 
rect 206 150 207 151 
rect 206 151 207 152 
rect 206 152 207 153 
rect 206 165 207 166 
rect 206 182 207 183 
rect 206 184 207 185 
rect 206 229 207 230 
rect 206 232 207 233 
rect 206 242 207 243 
rect 206 245 207 246 
rect 206 247 207 248 
rect 206 257 207 258 
rect 206 262 207 263 
rect 206 264 207 265 
rect 206 273 207 274 
rect 206 275 207 276 
rect 206 289 207 290 
rect 206 291 207 292 
rect 206 305 207 306 
rect 206 308 207 309 
rect 206 310 207 311 
rect 207 1 208 2 
rect 207 3 208 4 
rect 207 8 208 9 
rect 207 18 208 19 
rect 207 21 208 22 
rect 207 23 208 24 
rect 207 36 208 37 
rect 207 40 208 41 
rect 207 50 208 51 
rect 207 52 208 53 
rect 207 54 208 55 
rect 207 62 208 63 
rect 207 66 208 67 
rect 207 68 208 69 
rect 207 71 208 72 
rect 207 82 208 83 
rect 207 87 208 88 
rect 207 97 208 98 
rect 207 100 208 101 
rect 207 113 208 114 
rect 207 115 208 116 
rect 207 118 208 119 
rect 207 145 208 146 
rect 207 165 208 166 
rect 207 182 208 183 
rect 207 184 208 185 
rect 207 229 208 230 
rect 207 232 208 233 
rect 207 235 208 236 
rect 207 242 208 243 
rect 207 245 208 246 
rect 207 247 208 248 
rect 207 257 208 258 
rect 207 262 208 263 
rect 207 264 208 265 
rect 207 273 208 274 
rect 207 289 208 290 
rect 207 291 208 292 
rect 207 305 208 306 
rect 207 308 208 309 
rect 207 310 208 311 
rect 208 1 209 2 
rect 208 3 209 4 
rect 208 8 209 9 
rect 208 18 209 19 
rect 208 21 209 22 
rect 208 23 209 24 
rect 208 36 209 37 
rect 208 40 209 41 
rect 208 50 209 51 
rect 208 52 209 53 
rect 208 54 209 55 
rect 208 62 209 63 
rect 208 66 209 67 
rect 208 68 209 69 
rect 208 71 209 72 
rect 208 82 209 83 
rect 208 87 209 88 
rect 208 97 209 98 
rect 208 100 209 101 
rect 208 113 209 114 
rect 208 115 209 116 
rect 208 118 209 119 
rect 208 144 209 145 
rect 208 145 209 146 
rect 208 165 209 166 
rect 208 182 209 183 
rect 208 184 209 185 
rect 208 229 209 230 
rect 208 232 209 233 
rect 208 235 209 236 
rect 208 242 209 243 
rect 208 245 209 246 
rect 208 247 209 248 
rect 208 257 209 258 
rect 208 262 209 263 
rect 208 264 209 265 
rect 208 273 209 274 
rect 208 289 209 290 
rect 208 291 209 292 
rect 208 305 209 306 
rect 208 308 209 309 
rect 208 310 209 311 
rect 209 1 210 2 
rect 209 3 210 4 
rect 209 8 210 9 
rect 209 18 210 19 
rect 209 21 210 22 
rect 209 23 210 24 
rect 209 36 210 37 
rect 209 40 210 41 
rect 209 50 210 51 
rect 209 52 210 53 
rect 209 54 210 55 
rect 209 61 210 62 
rect 209 62 210 63 
rect 209 66 210 67 
rect 209 68 210 69 
rect 209 71 210 72 
rect 209 82 210 83 
rect 209 87 210 88 
rect 209 97 210 98 
rect 209 100 210 101 
rect 209 113 210 114 
rect 209 115 210 116 
rect 209 118 210 119 
rect 209 143 210 144 
rect 209 144 210 145 
rect 209 182 210 183 
rect 209 229 210 230 
rect 209 232 210 233 
rect 209 235 210 236 
rect 209 242 210 243 
rect 209 245 210 246 
rect 209 247 210 248 
rect 209 257 210 258 
rect 209 262 210 263 
rect 209 264 210 265 
rect 209 273 210 274 
rect 209 289 210 290 
rect 209 291 210 292 
rect 209 305 210 306 
rect 209 308 210 309 
rect 209 310 210 311 
rect 210 1 211 2 
rect 210 3 211 4 
rect 210 8 211 9 
rect 210 18 211 19 
rect 210 21 211 22 
rect 210 23 211 24 
rect 210 36 211 37 
rect 210 40 211 41 
rect 210 49 211 50 
rect 210 50 211 51 
rect 210 52 211 53 
rect 210 54 211 55 
rect 210 61 211 62 
rect 210 66 211 67 
rect 210 68 211 69 
rect 210 71 211 72 
rect 210 82 211 83 
rect 210 83 211 84 
rect 210 84 211 85 
rect 210 87 211 88 
rect 210 97 211 98 
rect 210 100 211 101 
rect 210 101 211 102 
rect 210 102 211 103 
rect 210 103 211 104 
rect 210 104 211 105 
rect 210 113 211 114 
rect 210 115 211 116 
rect 210 116 211 117 
rect 210 118 211 119 
rect 210 143 211 144 
rect 210 145 211 146 
rect 210 146 211 147 
rect 210 147 211 148 
rect 210 148 211 149 
rect 210 149 211 150 
rect 210 150 211 151 
rect 210 151 211 152 
rect 210 152 211 153 
rect 210 153 211 154 
rect 210 154 211 155 
rect 210 155 211 156 
rect 210 156 211 157 
rect 210 157 211 158 
rect 210 158 211 159 
rect 210 159 211 160 
rect 210 160 211 161 
rect 210 161 211 162 
rect 210 162 211 163 
rect 210 163 211 164 
rect 210 164 211 165 
rect 210 165 211 166 
rect 210 166 211 167 
rect 210 167 211 168 
rect 210 168 211 169 
rect 210 169 211 170 
rect 210 170 211 171 
rect 210 171 211 172 
rect 210 172 211 173 
rect 210 173 211 174 
rect 210 174 211 175 
rect 210 175 211 176 
rect 210 176 211 177 
rect 210 177 211 178 
rect 210 178 211 179 
rect 210 179 211 180 
rect 210 180 211 181 
rect 210 181 211 182 
rect 210 182 211 183 
rect 210 184 211 185 
rect 210 185 211 186 
rect 210 186 211 187 
rect 210 187 211 188 
rect 210 188 211 189 
rect 210 189 211 190 
rect 210 190 211 191 
rect 210 191 211 192 
rect 210 192 211 193 
rect 210 193 211 194 
rect 210 194 211 195 
rect 210 195 211 196 
rect 210 196 211 197 
rect 210 197 211 198 
rect 210 198 211 199 
rect 210 199 211 200 
rect 210 200 211 201 
rect 210 201 211 202 
rect 210 202 211 203 
rect 210 203 211 204 
rect 210 204 211 205 
rect 210 205 211 206 
rect 210 206 211 207 
rect 210 207 211 208 
rect 210 208 211 209 
rect 210 209 211 210 
rect 210 210 211 211 
rect 210 211 211 212 
rect 210 212 211 213 
rect 210 213 211 214 
rect 210 214 211 215 
rect 210 215 211 216 
rect 210 216 211 217 
rect 210 217 211 218 
rect 210 218 211 219 
rect 210 219 211 220 
rect 210 220 211 221 
rect 210 221 211 222 
rect 210 222 211 223 
rect 210 223 211 224 
rect 210 224 211 225 
rect 210 225 211 226 
rect 210 226 211 227 
rect 210 227 211 228 
rect 210 228 211 229 
rect 210 229 211 230 
rect 210 232 211 233 
rect 210 235 211 236 
rect 210 236 211 237 
rect 210 237 211 238 
rect 210 238 211 239 
rect 210 239 211 240 
rect 210 241 211 242 
rect 210 242 211 243 
rect 210 245 211 246 
rect 210 247 211 248 
rect 210 248 211 249 
rect 210 249 211 250 
rect 210 250 211 251 
rect 210 251 211 252 
rect 210 252 211 253 
rect 210 253 211 254 
rect 210 254 211 255 
rect 210 255 211 256 
rect 210 257 211 258 
rect 210 262 211 263 
rect 210 264 211 265 
rect 210 273 211 274 
rect 210 276 211 277 
rect 210 277 211 278 
rect 210 278 211 279 
rect 210 279 211 280 
rect 210 280 211 281 
rect 210 281 211 282 
rect 210 282 211 283 
rect 210 283 211 284 
rect 210 284 211 285 
rect 210 285 211 286 
rect 210 286 211 287 
rect 210 287 211 288 
rect 210 288 211 289 
rect 210 289 211 290 
rect 210 291 211 292 
rect 210 293 211 294 
rect 210 294 211 295 
rect 210 295 211 296 
rect 210 296 211 297 
rect 210 297 211 298 
rect 210 298 211 299 
rect 210 299 211 300 
rect 210 300 211 301 
rect 210 301 211 302 
rect 210 302 211 303 
rect 210 305 211 306 
rect 210 307 211 308 
rect 210 308 211 309 
rect 210 310 211 311 
rect 211 1 212 2 
rect 211 3 212 4 
rect 211 8 212 9 
rect 211 18 212 19 
rect 211 21 212 22 
rect 211 23 212 24 
rect 211 36 212 37 
rect 211 40 212 41 
rect 211 49 212 50 
rect 211 52 212 53 
rect 211 54 212 55 
rect 211 61 212 62 
rect 211 66 212 67 
rect 211 68 212 69 
rect 211 71 212 72 
rect 211 84 212 85 
rect 211 87 212 88 
rect 211 97 212 98 
rect 211 104 212 105 
rect 211 113 212 114 
rect 211 114 212 115 
rect 211 116 212 117 
rect 211 118 212 119 
rect 211 143 212 144 
rect 211 145 212 146 
rect 211 183 212 184 
rect 211 184 212 185 
rect 211 232 212 233 
rect 211 239 212 240 
rect 211 241 212 242 
rect 211 245 212 246 
rect 211 246 212 247 
rect 211 255 212 256 
rect 211 257 212 258 
rect 211 262 212 263 
rect 211 264 212 265 
rect 211 268 212 269 
rect 211 269 212 270 
rect 211 270 212 271 
rect 211 271 212 272 
rect 211 273 212 274 
rect 211 276 212 277 
rect 211 290 212 291 
rect 211 291 212 292 
rect 211 293 212 294 
rect 211 305 212 306 
rect 211 309 212 310 
rect 211 310 212 311 
rect 212 1 213 2 
rect 212 3 213 4 
rect 212 8 213 9 
rect 212 18 213 19 
rect 212 21 213 22 
rect 212 23 213 24 
rect 212 36 213 37 
rect 212 40 213 41 
rect 212 49 213 50 
rect 212 52 213 53 
rect 212 54 213 55 
rect 212 61 213 62 
rect 212 66 213 67 
rect 212 68 213 69 
rect 212 71 213 72 
rect 212 84 213 85 
rect 212 87 213 88 
rect 212 97 213 98 
rect 212 104 213 105 
rect 212 114 213 115 
rect 212 116 213 117 
rect 212 118 213 119 
rect 212 143 213 144 
rect 212 145 213 146 
rect 212 148 213 149 
rect 212 149 213 150 
rect 212 150 213 151 
rect 212 151 213 152 
rect 212 152 213 153 
rect 212 153 213 154 
rect 212 154 213 155 
rect 212 155 213 156 
rect 212 156 213 157 
rect 212 157 213 158 
rect 212 158 213 159 
rect 212 159 213 160 
rect 212 160 213 161 
rect 212 161 213 162 
rect 212 162 213 163 
rect 212 163 213 164 
rect 212 164 213 165 
rect 212 165 213 166 
rect 212 166 213 167 
rect 212 167 213 168 
rect 212 168 213 169 
rect 212 169 213 170 
rect 212 170 213 171 
rect 212 171 213 172 
rect 212 172 213 173 
rect 212 173 213 174 
rect 212 174 213 175 
rect 212 175 213 176 
rect 212 176 213 177 
rect 212 177 213 178 
rect 212 178 213 179 
rect 212 179 213 180 
rect 212 180 213 181 
rect 212 181 213 182 
rect 212 182 213 183 
rect 212 183 213 184 
rect 212 232 213 233 
rect 212 239 213 240 
rect 212 241 213 242 
rect 212 243 213 244 
rect 212 244 213 245 
rect 212 246 213 247 
rect 212 247 213 248 
rect 212 248 213 249 
rect 212 249 213 250 
rect 212 250 213 251 
rect 212 251 213 252 
rect 212 252 213 253 
rect 212 253 213 254 
rect 212 255 213 256 
rect 212 257 213 258 
rect 212 262 213 263 
rect 212 264 213 265 
rect 212 268 213 269 
rect 212 273 213 274 
rect 212 276 213 277 
rect 212 279 213 280 
rect 212 285 213 286 
rect 212 286 213 287 
rect 212 287 213 288 
rect 212 288 213 289 
rect 212 289 213 290 
rect 212 290 213 291 
rect 212 293 213 294 
rect 212 305 213 306 
rect 212 307 213 308 
rect 212 308 213 309 
rect 212 309 213 310 
rect 213 1 214 2 
rect 213 3 214 4 
rect 213 8 214 9 
rect 213 18 214 19 
rect 213 21 214 22 
rect 213 23 214 24 
rect 213 36 214 37 
rect 213 40 214 41 
rect 213 49 214 50 
rect 213 52 214 53 
rect 213 54 214 55 
rect 213 61 214 62 
rect 213 66 214 67 
rect 213 68 214 69 
rect 213 71 214 72 
rect 213 84 214 85 
rect 213 87 214 88 
rect 213 97 214 98 
rect 213 104 214 105 
rect 213 114 214 115 
rect 213 116 214 117 
rect 213 118 214 119 
rect 213 143 214 144 
rect 213 145 214 146 
rect 213 148 214 149 
rect 213 232 214 233 
rect 213 239 214 240 
rect 213 241 214 242 
rect 213 244 214 245 
rect 213 245 214 246 
rect 213 255 214 256 
rect 213 257 214 258 
rect 213 262 214 263 
rect 213 264 214 265 
rect 213 268 214 269 
rect 213 273 214 274 
rect 213 276 214 277 
rect 213 279 214 280 
rect 213 280 214 281 
rect 213 281 214 282 
rect 213 282 214 283 
rect 213 283 214 284 
rect 213 284 214 285 
rect 213 285 214 286 
rect 213 293 214 294 
rect 213 305 214 306 
rect 213 307 214 308 
rect 214 1 215 2 
rect 214 3 215 4 
rect 214 8 215 9 
rect 214 18 215 19 
rect 214 21 215 22 
rect 214 23 215 24 
rect 214 36 215 37 
rect 214 40 215 41 
rect 214 49 215 50 
rect 214 52 215 53 
rect 214 54 215 55 
rect 214 61 215 62 
rect 214 66 215 67 
rect 214 68 215 69 
rect 214 71 215 72 
rect 214 84 215 85 
rect 214 87 215 88 
rect 214 97 215 98 
rect 214 104 215 105 
rect 214 114 215 115 
rect 214 116 215 117 
rect 214 118 215 119 
rect 214 143 215 144 
rect 214 145 215 146 
rect 214 148 215 149 
rect 214 151 215 152 
rect 214 152 215 153 
rect 214 155 215 156 
rect 214 156 215 157 
rect 214 157 215 158 
rect 214 158 215 159 
rect 214 159 215 160 
rect 214 160 215 161 
rect 214 164 215 165 
rect 214 165 215 166 
rect 214 166 215 167 
rect 214 167 215 168 
rect 214 168 215 169 
rect 214 169 215 170 
rect 214 170 215 171 
rect 214 171 215 172 
rect 214 172 215 173 
rect 214 173 215 174 
rect 214 174 215 175 
rect 214 175 215 176 
rect 214 176 215 177 
rect 214 177 215 178 
rect 214 178 215 179 
rect 214 179 215 180 
rect 214 180 215 181 
rect 214 181 215 182 
rect 214 182 215 183 
rect 214 183 215 184 
rect 214 184 215 185 
rect 214 185 215 186 
rect 214 186 215 187 
rect 214 187 215 188 
rect 214 188 215 189 
rect 214 189 215 190 
rect 214 190 215 191 
rect 214 191 215 192 
rect 214 192 215 193 
rect 214 193 215 194 
rect 214 194 215 195 
rect 214 195 215 196 
rect 214 196 215 197 
rect 214 197 215 198 
rect 214 198 215 199 
rect 214 199 215 200 
rect 214 200 215 201 
rect 214 201 215 202 
rect 214 202 215 203 
rect 214 203 215 204 
rect 214 204 215 205 
rect 214 205 215 206 
rect 214 206 215 207 
rect 214 207 215 208 
rect 214 208 215 209 
rect 214 209 215 210 
rect 214 210 215 211 
rect 214 211 215 212 
rect 214 212 215 213 
rect 214 213 215 214 
rect 214 214 215 215 
rect 214 215 215 216 
rect 214 216 215 217 
rect 214 217 215 218 
rect 214 218 215 219 
rect 214 219 215 220 
rect 214 220 215 221 
rect 214 221 215 222 
rect 214 222 215 223 
rect 214 223 215 224 
rect 214 224 215 225 
rect 214 225 215 226 
rect 214 226 215 227 
rect 214 227 215 228 
rect 214 228 215 229 
rect 214 229 215 230 
rect 214 230 215 231 
rect 214 232 215 233 
rect 214 239 215 240 
rect 214 241 215 242 
rect 214 245 215 246 
rect 214 246 215 247 
rect 214 247 215 248 
rect 214 248 215 249 
rect 214 249 215 250 
rect 214 250 215 251 
rect 214 251 215 252 
rect 214 252 215 253 
rect 214 255 215 256 
rect 214 257 215 258 
rect 214 262 215 263 
rect 214 264 215 265 
rect 214 266 215 267 
rect 214 267 215 268 
rect 214 268 215 269 
rect 214 273 215 274 
rect 214 276 215 277 
rect 214 293 215 294 
rect 214 305 215 306 
rect 214 307 215 308 
rect 215 1 216 2 
rect 215 3 216 4 
rect 215 8 216 9 
rect 215 18 216 19 
rect 215 21 216 22 
rect 215 23 216 24 
rect 215 36 216 37 
rect 215 40 216 41 
rect 215 49 216 50 
rect 215 52 216 53 
rect 215 54 216 55 
rect 215 61 216 62 
rect 215 66 216 67 
rect 215 68 216 69 
rect 215 71 216 72 
rect 215 84 216 85 
rect 215 87 216 88 
rect 215 97 216 98 
rect 215 104 216 105 
rect 215 116 216 117 
rect 215 118 216 119 
rect 215 143 216 144 
rect 215 145 216 146 
rect 215 148 216 149 
rect 215 152 216 153 
rect 215 155 216 156 
rect 215 232 216 233 
rect 215 239 216 240 
rect 215 241 216 242 
rect 215 243 216 244 
rect 215 255 216 256 
rect 215 257 216 258 
rect 215 262 216 263 
rect 215 264 216 265 
rect 215 273 216 274 
rect 215 276 216 277 
rect 215 293 216 294 
rect 215 305 216 306 
rect 215 307 216 308 
rect 215 309 216 310 
rect 216 1 217 2 
rect 216 3 217 4 
rect 216 8 217 9 
rect 216 18 217 19 
rect 216 21 217 22 
rect 216 23 217 24 
rect 216 36 217 37 
rect 216 40 217 41 
rect 216 49 217 50 
rect 216 52 217 53 
rect 216 54 217 55 
rect 216 57 217 58 
rect 216 58 217 59 
rect 216 59 217 60 
rect 216 60 217 61 
rect 216 61 217 62 
rect 216 66 217 67 
rect 216 68 217 69 
rect 216 71 217 72 
rect 216 84 217 85 
rect 216 87 217 88 
rect 216 97 217 98 
rect 216 104 217 105 
rect 216 114 217 115 
rect 216 116 217 117 
rect 216 118 217 119 
rect 216 121 217 122 
rect 216 122 217 123 
rect 216 123 217 124 
rect 216 124 217 125 
rect 216 125 217 126 
rect 216 126 217 127 
rect 216 127 217 128 
rect 216 128 217 129 
rect 216 129 217 130 
rect 216 137 217 138 
rect 216 138 217 139 
rect 216 139 217 140 
rect 216 140 217 141 
rect 216 141 217 142 
rect 216 142 217 143 
rect 216 143 217 144 
rect 216 145 217 146 
rect 216 148 217 149 
rect 216 152 217 153 
rect 216 155 217 156 
rect 216 168 217 169 
rect 216 169 217 170 
rect 216 170 217 171 
rect 216 171 217 172 
rect 216 172 217 173 
rect 216 173 217 174 
rect 216 174 217 175 
rect 216 175 217 176 
rect 216 176 217 177 
rect 216 177 217 178 
rect 216 178 217 179 
rect 216 179 217 180 
rect 216 180 217 181 
rect 216 181 217 182 
rect 216 182 217 183 
rect 216 183 217 184 
rect 216 184 217 185 
rect 216 185 217 186 
rect 216 186 217 187 
rect 216 187 217 188 
rect 216 188 217 189 
rect 216 189 217 190 
rect 216 190 217 191 
rect 216 191 217 192 
rect 216 192 217 193 
rect 216 193 217 194 
rect 216 194 217 195 
rect 216 195 217 196 
rect 216 196 217 197 
rect 216 201 217 202 
rect 216 202 217 203 
rect 216 203 217 204 
rect 216 232 217 233 
rect 216 239 217 240 
rect 216 241 217 242 
rect 216 243 217 244 
rect 216 244 217 245 
rect 216 245 217 246 
rect 216 246 217 247 
rect 216 247 217 248 
rect 216 248 217 249 
rect 216 249 217 250 
rect 216 250 217 251 
rect 216 251 217 252 
rect 216 255 217 256 
rect 216 257 217 258 
rect 216 262 217 263 
rect 216 264 217 265 
rect 216 273 217 274 
rect 216 276 217 277 
rect 216 293 217 294 
rect 216 297 217 298 
rect 216 298 217 299 
rect 216 299 217 300 
rect 216 305 217 306 
rect 216 307 217 308 
rect 216 309 217 310 
rect 217 1 218 2 
rect 217 3 218 4 
rect 217 8 218 9 
rect 217 18 218 19 
rect 217 21 218 22 
rect 217 23 218 24 
rect 217 36 218 37 
rect 217 40 218 41 
rect 217 49 218 50 
rect 217 52 218 53 
rect 217 54 218 55 
rect 217 56 218 57 
rect 217 57 218 58 
rect 217 66 218 67 
rect 217 68 218 69 
rect 217 71 218 72 
rect 217 84 218 85 
rect 217 87 218 88 
rect 217 97 218 98 
rect 217 104 218 105 
rect 217 114 218 115 
rect 217 116 218 117 
rect 217 118 218 119 
rect 217 129 218 130 
rect 217 130 218 131 
rect 217 131 218 132 
rect 217 132 218 133 
rect 217 133 218 134 
rect 217 134 218 135 
rect 217 135 218 136 
rect 217 136 218 137 
rect 217 137 218 138 
rect 217 145 218 146 
rect 217 148 218 149 
rect 217 152 218 153 
rect 217 155 218 156 
rect 217 168 218 169 
rect 217 200 218 201 
rect 217 201 218 202 
rect 217 203 218 204 
rect 217 232 218 233 
rect 217 241 218 242 
rect 217 251 218 252 
rect 217 257 218 258 
rect 217 262 218 263 
rect 217 264 218 265 
rect 217 273 218 274 
rect 217 276 218 277 
rect 217 293 218 294 
rect 217 295 218 296 
rect 217 296 218 297 
rect 217 297 218 298 
rect 217 299 218 300 
rect 217 305 218 306 
rect 217 307 218 308 
rect 217 309 218 310 
rect 218 1 219 2 
rect 218 3 219 4 
rect 218 8 219 9 
rect 218 18 219 19 
rect 218 21 219 22 
rect 218 23 219 24 
rect 218 36 219 37 
rect 218 40 219 41 
rect 218 49 219 50 
rect 218 52 219 53 
rect 218 54 219 55 
rect 218 56 219 57 
rect 218 66 219 67 
rect 218 68 219 69 
rect 218 71 219 72 
rect 218 84 219 85 
rect 218 87 219 88 
rect 218 97 219 98 
rect 218 104 219 105 
rect 218 114 219 115 
rect 218 116 219 117 
rect 218 118 219 119 
rect 218 145 219 146 
rect 218 148 219 149 
rect 218 152 219 153 
rect 218 155 219 156 
rect 218 168 219 169 
rect 218 200 219 201 
rect 218 203 219 204 
rect 218 232 219 233 
rect 218 241 219 242 
rect 218 251 219 252 
rect 218 257 219 258 
rect 218 262 219 263 
rect 218 264 219 265 
rect 218 273 219 274 
rect 218 276 219 277 
rect 218 289 219 290 
rect 218 290 219 291 
rect 218 291 219 292 
rect 218 292 219 293 
rect 218 293 219 294 
rect 218 299 219 300 
rect 218 305 219 306 
rect 218 307 219 308 
rect 218 309 219 310 
rect 219 1 220 2 
rect 219 3 220 4 
rect 219 8 220 9 
rect 219 18 220 19 
rect 219 21 220 22 
rect 219 23 220 24 
rect 219 36 220 37 
rect 219 40 220 41 
rect 219 49 220 50 
rect 219 52 220 53 
rect 219 54 220 55 
rect 219 56 220 57 
rect 219 66 220 67 
rect 219 68 220 69 
rect 219 71 220 72 
rect 219 84 220 85 
rect 219 87 220 88 
rect 219 97 220 98 
rect 219 104 220 105 
rect 219 114 220 115 
rect 219 116 220 117 
rect 219 118 220 119 
rect 219 145 220 146 
rect 219 148 220 149 
rect 219 152 220 153 
rect 219 168 220 169 
rect 219 200 220 201 
rect 219 232 220 233 
rect 219 241 220 242 
rect 219 257 220 258 
rect 219 262 220 263 
rect 219 264 220 265 
rect 219 273 220 274 
rect 219 276 220 277 
rect 219 289 220 290 
rect 219 305 220 306 
rect 219 307 220 308 
rect 219 309 220 310 
rect 220 1 221 2 
rect 220 3 221 4 
rect 220 8 221 9 
rect 220 18 221 19 
rect 220 21 221 22 
rect 220 23 221 24 
rect 220 36 221 37 
rect 220 40 221 41 
rect 220 49 221 50 
rect 220 52 221 53 
rect 220 54 221 55 
rect 220 56 221 57 
rect 220 66 221 67 
rect 220 68 221 69 
rect 220 71 221 72 
rect 220 84 221 85 
rect 220 87 221 88 
rect 220 97 221 98 
rect 220 104 221 105 
rect 220 114 221 115 
rect 220 116 221 117 
rect 220 118 221 119 
rect 220 145 221 146 
rect 220 148 221 149 
rect 220 152 221 153 
rect 220 168 221 169 
rect 220 200 221 201 
rect 220 232 221 233 
rect 220 241 221 242 
rect 220 257 221 258 
rect 220 262 221 263 
rect 220 264 221 265 
rect 220 273 221 274 
rect 220 276 221 277 
rect 220 289 221 290 
rect 220 292 221 293 
rect 220 293 221 294 
rect 220 305 221 306 
rect 220 307 221 308 
rect 220 309 221 310 
rect 221 1 222 2 
rect 221 3 222 4 
rect 221 8 222 9 
rect 221 18 222 19 
rect 221 21 222 22 
rect 221 23 222 24 
rect 221 36 222 37 
rect 221 40 222 41 
rect 221 49 222 50 
rect 221 52 222 53 
rect 221 54 222 55 
rect 221 56 222 57 
rect 221 66 222 67 
rect 221 68 222 69 
rect 221 71 222 72 
rect 221 84 222 85 
rect 221 87 222 88 
rect 221 97 222 98 
rect 221 104 222 105 
rect 221 114 222 115 
rect 221 116 222 117 
rect 221 118 222 119 
rect 221 145 222 146 
rect 221 148 222 149 
rect 221 152 222 153 
rect 221 168 222 169 
rect 221 200 222 201 
rect 221 232 222 233 
rect 221 241 222 242 
rect 221 257 222 258 
rect 221 262 222 263 
rect 221 264 222 265 
rect 221 273 222 274 
rect 221 276 222 277 
rect 221 289 222 290 
rect 221 293 222 294 
rect 221 305 222 306 
rect 221 307 222 308 
rect 221 309 222 310 
rect 222 1 223 2 
rect 222 3 223 4 
rect 222 8 223 9 
rect 222 18 223 19 
rect 222 21 223 22 
rect 222 23 223 24 
rect 222 36 223 37 
rect 222 40 223 41 
rect 222 49 223 50 
rect 222 52 223 53 
rect 222 54 223 55 
rect 222 56 223 57 
rect 222 66 223 67 
rect 222 68 223 69 
rect 222 71 223 72 
rect 222 87 223 88 
rect 222 97 223 98 
rect 222 104 223 105 
rect 222 114 223 115 
rect 222 116 223 117 
rect 222 118 223 119 
rect 222 145 223 146 
rect 222 148 223 149 
rect 222 152 223 153 
rect 222 168 223 169 
rect 222 200 223 201 
rect 222 232 223 233 
rect 222 241 223 242 
rect 222 257 223 258 
rect 222 262 223 263 
rect 222 264 223 265 
rect 222 273 223 274 
rect 222 276 223 277 
rect 222 289 223 290 
rect 222 293 223 294 
rect 222 305 223 306 
rect 222 307 223 308 
rect 222 309 223 310 
rect 223 1 224 2 
rect 223 3 224 4 
rect 223 8 224 9 
rect 223 18 224 19 
rect 223 21 224 22 
rect 223 23 224 24 
rect 223 27 224 28 
rect 223 36 224 37 
rect 223 40 224 41 
rect 223 49 224 50 
rect 223 52 224 53 
rect 223 54 224 55 
rect 223 56 224 57 
rect 223 66 224 67 
rect 223 68 224 69 
rect 223 71 224 72 
rect 223 81 224 82 
rect 223 82 224 83 
rect 223 83 224 84 
rect 223 84 224 85 
rect 223 85 224 86 
rect 223 86 224 87 
rect 223 87 224 88 
rect 223 97 224 98 
rect 223 104 224 105 
rect 223 114 224 115 
rect 223 116 224 117 
rect 223 118 224 119 
rect 223 139 224 140 
rect 223 145 224 146 
rect 223 148 224 149 
rect 223 152 224 153 
rect 223 168 224 169 
rect 223 200 224 201 
rect 223 232 224 233 
rect 223 241 224 242 
rect 223 257 224 258 
rect 223 262 224 263 
rect 223 264 224 265 
rect 223 273 224 274 
rect 223 276 224 277 
rect 223 289 224 290 
rect 223 293 224 294 
rect 223 305 224 306 
rect 223 307 224 308 
rect 223 309 224 310 
rect 224 1 225 2 
rect 224 3 225 4 
rect 224 8 225 9 
rect 224 18 225 19 
rect 224 21 225 22 
rect 224 23 225 24 
rect 224 27 225 28 
rect 224 32 225 33 
rect 224 33 225 34 
rect 224 34 225 35 
rect 224 35 225 36 
rect 224 36 225 37 
rect 224 40 225 41 
rect 224 48 225 49 
rect 224 49 225 50 
rect 224 52 225 53 
rect 224 54 225 55 
rect 224 66 225 67 
rect 224 68 225 69 
rect 224 71 225 72 
rect 224 80 225 81 
rect 224 81 225 82 
rect 224 97 225 98 
rect 224 104 225 105 
rect 224 105 225 106 
rect 224 114 225 115 
rect 224 116 225 117 
rect 224 118 225 119 
rect 224 129 225 130 
rect 224 130 225 131 
rect 224 131 225 132 
rect 224 132 225 133 
rect 224 133 225 134 
rect 224 134 225 135 
rect 224 135 225 136 
rect 224 136 225 137 
rect 224 137 225 138 
rect 224 139 225 140 
rect 224 144 225 145 
rect 224 145 225 146 
rect 224 148 225 149 
rect 224 152 225 153 
rect 224 153 225 154 
rect 224 208 225 209 
rect 224 209 225 210 
rect 224 210 225 211 
rect 224 211 225 212 
rect 224 212 225 213 
rect 224 213 225 214 
rect 224 214 225 215 
rect 224 215 225 216 
rect 224 216 225 217 
rect 224 224 225 225 
rect 224 225 225 226 
rect 224 226 225 227 
rect 224 227 225 228 
rect 224 228 225 229 
rect 224 229 225 230 
rect 224 230 225 231 
rect 224 232 225 233 
rect 224 240 225 241 
rect 224 241 225 242 
rect 224 256 225 257 
rect 224 257 225 258 
rect 224 262 225 263 
rect 224 264 225 265 
rect 224 273 225 274 
rect 224 276 225 277 
rect 224 288 225 289 
rect 224 289 225 290 
rect 224 293 225 294 
rect 224 294 225 295 
rect 224 295 225 296 
rect 224 296 225 297 
rect 224 297 225 298 
rect 224 305 225 306 
rect 224 307 225 308 
rect 224 309 225 310 
rect 225 1 226 2 
rect 225 3 226 4 
rect 225 8 226 9 
rect 225 18 226 19 
rect 225 21 226 22 
rect 225 23 226 24 
rect 225 27 226 28 
rect 225 28 226 29 
rect 225 30 226 31 
rect 225 31 226 32 
rect 225 32 226 33 
rect 225 40 226 41 
rect 225 43 226 44 
rect 225 44 226 45 
rect 225 45 226 46 
rect 225 46 226 47 
rect 225 47 226 48 
rect 225 48 226 49 
rect 225 51 226 52 
rect 225 66 226 67 
rect 225 68 226 69 
rect 225 71 226 72 
rect 225 80 226 81 
rect 225 97 226 98 
rect 225 105 226 106 
rect 225 106 226 107 
rect 225 107 226 108 
rect 225 108 226 109 
rect 225 109 226 110 
rect 225 110 226 111 
rect 225 111 226 112 
rect 225 112 226 113 
rect 225 114 226 115 
rect 225 116 226 117 
rect 225 118 226 119 
rect 225 121 226 122 
rect 225 122 226 123 
rect 225 123 226 124 
rect 225 124 226 125 
rect 225 125 226 126 
rect 225 126 226 127 
rect 225 127 226 128 
rect 225 128 226 129 
rect 225 129 226 130 
rect 225 137 226 138 
rect 225 139 226 140 
rect 225 140 226 141 
rect 225 141 226 142 
rect 225 142 226 143 
rect 225 143 226 144 
rect 225 144 226 145 
rect 225 148 226 149 
rect 225 153 226 154 
rect 225 154 226 155 
rect 225 155 226 156 
rect 225 156 226 157 
rect 225 157 226 158 
rect 225 158 226 159 
rect 225 159 226 160 
rect 225 160 226 161 
rect 225 161 226 162 
rect 225 162 226 163 
rect 225 163 226 164 
rect 225 164 226 165 
rect 225 165 226 166 
rect 225 166 226 167 
rect 225 167 226 168 
rect 225 168 226 169 
rect 225 169 226 170 
rect 225 170 226 171 
rect 225 171 226 172 
rect 225 172 226 173 
rect 225 173 226 174 
rect 225 174 226 175 
rect 225 175 226 176 
rect 225 176 226 177 
rect 225 177 226 178 
rect 225 178 226 179 
rect 225 179 226 180 
rect 225 180 226 181 
rect 225 181 226 182 
rect 225 182 226 183 
rect 225 183 226 184 
rect 225 184 226 185 
rect 225 185 226 186 
rect 225 187 226 188 
rect 225 188 226 189 
rect 225 189 226 190 
rect 225 190 226 191 
rect 225 191 226 192 
rect 225 192 226 193 
rect 225 193 226 194 
rect 225 194 226 195 
rect 225 195 226 196 
rect 225 196 226 197 
rect 225 197 226 198 
rect 225 198 226 199 
rect 225 199 226 200 
rect 225 200 226 201 
rect 225 201 226 202 
rect 225 202 226 203 
rect 225 203 226 204 
rect 225 204 226 205 
rect 225 205 226 206 
rect 225 206 226 207 
rect 225 207 226 208 
rect 225 208 226 209 
rect 225 216 226 217 
rect 225 217 226 218 
rect 225 218 226 219 
rect 225 219 226 220 
rect 225 220 226 221 
rect 225 221 226 222 
rect 225 222 226 223 
rect 225 223 226 224 
rect 225 224 226 225 
rect 225 232 226 233 
rect 225 234 226 235 
rect 225 235 226 236 
rect 225 236 226 237 
rect 225 237 226 238 
rect 225 238 226 239 
rect 225 239 226 240 
rect 225 240 226 241 
rect 225 244 226 245 
rect 225 245 226 246 
rect 225 246 226 247 
rect 225 247 226 248 
rect 225 248 226 249 
rect 225 249 226 250 
rect 225 250 226 251 
rect 225 251 226 252 
rect 225 252 226 253 
rect 225 253 226 254 
rect 225 254 226 255 
rect 225 255 226 256 
rect 225 256 226 257 
rect 225 258 226 259 
rect 225 259 226 260 
rect 225 260 226 261 
rect 225 262 226 263 
rect 225 264 226 265 
rect 225 265 226 266 
rect 225 266 226 267 
rect 225 267 226 268 
rect 225 268 226 269 
rect 225 269 226 270 
rect 225 270 226 271 
rect 225 273 226 274 
rect 225 276 226 277 
rect 225 278 226 279 
rect 225 279 226 280 
rect 225 280 226 281 
rect 225 281 226 282 
rect 225 282 226 283 
rect 225 283 226 284 
rect 225 284 226 285 
rect 225 285 226 286 
rect 225 286 226 287 
rect 225 287 226 288 
rect 225 288 226 289 
rect 225 297 226 298 
rect 225 298 226 299 
rect 225 299 226 300 
rect 225 300 226 301 
rect 225 301 226 302 
rect 225 302 226 303 
rect 225 305 226 306 
rect 225 307 226 308 
rect 225 309 226 310 
rect 226 1 227 2 
rect 226 3 227 4 
rect 226 8 227 9 
rect 226 18 227 19 
rect 226 21 227 22 
rect 226 23 227 24 
rect 226 30 227 31 
rect 226 40 227 41 
rect 226 43 227 44 
rect 226 51 227 52 
rect 226 52 227 53 
rect 226 53 227 54 
rect 226 54 227 55 
rect 226 55 227 56 
rect 226 56 227 57 
rect 226 57 227 58 
rect 226 58 227 59 
rect 226 59 227 60 
rect 226 60 227 61 
rect 226 61 227 62 
rect 226 62 227 63 
rect 226 63 227 64 
rect 226 64 227 65 
rect 226 66 227 67 
rect 226 68 227 69 
rect 226 71 227 72 
rect 226 74 227 75 
rect 226 80 227 81 
rect 226 97 227 98 
rect 226 112 227 113 
rect 226 114 227 115 
rect 226 118 227 119 
rect 226 137 227 138 
rect 226 138 227 139 
rect 226 187 227 188 
rect 226 232 227 233 
rect 226 242 227 243 
rect 226 244 227 245 
rect 226 257 227 258 
rect 226 258 227 259 
rect 226 262 227 263 
rect 226 270 227 271 
rect 226 273 227 274 
rect 226 276 227 277 
rect 226 278 227 279 
rect 226 302 227 303 
rect 226 305 227 306 
rect 226 307 227 308 
rect 226 309 227 310 
rect 227 1 228 2 
rect 227 3 228 4 
rect 227 8 228 9 
rect 227 18 228 19 
rect 227 21 228 22 
rect 227 23 228 24 
rect 227 30 228 31 
rect 227 40 228 41 
rect 227 43 228 44 
rect 227 66 228 67 
rect 227 68 228 69 
rect 227 71 228 72 
rect 227 74 228 75 
rect 227 75 228 76 
rect 227 76 228 77 
rect 227 77 228 78 
rect 227 78 228 79 
rect 227 79 228 80 
rect 227 80 228 81 
rect 227 97 228 98 
rect 227 112 228 113 
rect 227 114 228 115 
rect 227 118 228 119 
rect 227 138 228 139 
rect 227 139 228 140 
rect 227 140 228 141 
rect 227 141 228 142 
rect 227 142 228 143 
rect 227 143 228 144 
rect 227 144 228 145 
rect 227 145 228 146 
rect 227 146 228 147 
rect 227 147 228 148 
rect 227 148 228 149 
rect 227 149 228 150 
rect 227 150 228 151 
rect 227 151 228 152 
rect 227 152 228 153 
rect 227 153 228 154 
rect 227 154 228 155 
rect 227 155 228 156 
rect 227 156 228 157 
rect 227 157 228 158 
rect 227 158 228 159 
rect 227 159 228 160 
rect 227 160 228 161 
rect 227 161 228 162 
rect 227 162 228 163 
rect 227 163 228 164 
rect 227 164 228 165 
rect 227 165 228 166 
rect 227 166 228 167 
rect 227 167 228 168 
rect 227 168 228 169 
rect 227 169 228 170 
rect 227 170 228 171 
rect 227 171 228 172 
rect 227 172 228 173 
rect 227 173 228 174 
rect 227 174 228 175 
rect 227 175 228 176 
rect 227 176 228 177 
rect 227 177 228 178 
rect 227 178 228 179 
rect 227 179 228 180 
rect 227 180 228 181 
rect 227 181 228 182 
rect 227 182 228 183 
rect 227 183 228 184 
rect 227 184 228 185 
rect 227 185 228 186 
rect 227 187 228 188 
rect 227 190 228 191 
rect 227 191 228 192 
rect 227 192 228 193 
rect 227 193 228 194 
rect 227 194 228 195 
rect 227 195 228 196 
rect 227 196 228 197 
rect 227 197 228 198 
rect 227 198 228 199 
rect 227 199 228 200 
rect 227 200 228 201 
rect 227 201 228 202 
rect 227 202 228 203 
rect 227 203 228 204 
rect 227 204 228 205 
rect 227 205 228 206 
rect 227 206 228 207 
rect 227 207 228 208 
rect 227 208 228 209 
rect 227 209 228 210 
rect 227 210 228 211 
rect 227 211 228 212 
rect 227 212 228 213 
rect 227 213 228 214 
rect 227 214 228 215 
rect 227 215 228 216 
rect 227 216 228 217 
rect 227 217 228 218 
rect 227 218 228 219 
rect 227 219 228 220 
rect 227 220 228 221 
rect 227 221 228 222 
rect 227 222 228 223 
rect 227 223 228 224 
rect 227 224 228 225 
rect 227 225 228 226 
rect 227 226 228 227 
rect 227 227 228 228 
rect 227 228 228 229 
rect 227 229 228 230 
rect 227 232 228 233 
rect 227 242 228 243 
rect 227 244 228 245 
rect 227 247 228 248 
rect 227 253 228 254 
rect 227 254 228 255 
rect 227 255 228 256 
rect 227 256 228 257 
rect 227 257 228 258 
rect 227 262 228 263 
rect 227 270 228 271 
rect 227 273 228 274 
rect 227 276 228 277 
rect 227 278 228 279 
rect 227 293 228 294 
rect 227 302 228 303 
rect 227 305 228 306 
rect 227 308 228 309 
rect 227 309 228 310 
rect 228 1 229 2 
rect 228 3 229 4 
rect 228 8 229 9 
rect 228 18 229 19 
rect 228 21 229 22 
rect 228 23 229 24 
rect 228 30 229 31 
rect 228 40 229 41 
rect 228 43 229 44 
rect 228 53 229 54 
rect 228 54 229 55 
rect 228 55 229 56 
rect 228 56 229 57 
rect 228 57 229 58 
rect 228 58 229 59 
rect 228 59 229 60 
rect 228 60 229 61 
rect 228 61 229 62 
rect 228 62 229 63 
rect 228 63 229 64 
rect 228 64 229 65 
rect 228 66 229 67 
rect 228 68 229 69 
rect 228 71 229 72 
rect 228 97 229 98 
rect 228 112 229 113 
rect 228 114 229 115 
rect 228 118 229 119 
rect 228 187 229 188 
rect 228 229 229 230 
rect 228 232 229 233 
rect 228 242 229 243 
rect 228 244 229 245 
rect 228 247 229 248 
rect 228 248 229 249 
rect 228 249 229 250 
rect 228 250 229 251 
rect 228 251 229 252 
rect 228 252 229 253 
rect 228 253 229 254 
rect 228 262 229 263 
rect 228 270 229 271 
rect 228 273 229 274 
rect 228 276 229 277 
rect 228 278 229 279 
rect 228 293 229 294 
rect 228 302 229 303 
rect 228 305 229 306 
rect 228 307 229 308 
rect 228 308 229 309 
rect 229 1 230 2 
rect 229 3 230 4 
rect 229 8 230 9 
rect 229 18 230 19 
rect 229 21 230 22 
rect 229 23 230 24 
rect 229 30 230 31 
rect 229 40 230 41 
rect 229 43 230 44 
rect 229 66 230 67 
rect 229 68 230 69 
rect 229 71 230 72 
rect 229 73 230 74 
rect 229 74 230 75 
rect 229 75 230 76 
rect 229 76 230 77 
rect 229 77 230 78 
rect 229 78 230 79 
rect 229 79 230 80 
rect 229 80 230 81 
rect 229 81 230 82 
rect 229 82 230 83 
rect 229 83 230 84 
rect 229 84 230 85 
rect 229 85 230 86 
rect 229 86 230 87 
rect 229 87 230 88 
rect 229 88 230 89 
rect 229 89 230 90 
rect 229 90 230 91 
rect 229 91 230 92 
rect 229 92 230 93 
rect 229 93 230 94 
rect 229 94 230 95 
rect 229 95 230 96 
rect 229 97 230 98 
rect 229 101 230 102 
rect 229 102 230 103 
rect 229 103 230 104 
rect 229 104 230 105 
rect 229 105 230 106 
rect 229 106 230 107 
rect 229 107 230 108 
rect 229 108 230 109 
rect 229 109 230 110 
rect 229 110 230 111 
rect 229 112 230 113 
rect 229 114 230 115 
rect 229 118 230 119 
rect 229 187 230 188 
rect 229 192 230 193 
rect 229 193 230 194 
rect 229 194 230 195 
rect 229 195 230 196 
rect 229 196 230 197 
rect 229 197 230 198 
rect 229 198 230 199 
rect 229 199 230 200 
rect 229 200 230 201 
rect 229 201 230 202 
rect 229 202 230 203 
rect 229 203 230 204 
rect 229 204 230 205 
rect 229 205 230 206 
rect 229 206 230 207 
rect 229 207 230 208 
rect 229 208 230 209 
rect 229 209 230 210 
rect 229 210 230 211 
rect 229 211 230 212 
rect 229 212 230 213 
rect 229 213 230 214 
rect 229 214 230 215 
rect 229 215 230 216 
rect 229 216 230 217 
rect 229 217 230 218 
rect 229 218 230 219 
rect 229 219 230 220 
rect 229 220 230 221 
rect 229 221 230 222 
rect 229 222 230 223 
rect 229 223 230 224 
rect 229 224 230 225 
rect 229 225 230 226 
rect 229 229 230 230 
rect 229 232 230 233 
rect 229 242 230 243 
rect 229 244 230 245 
rect 229 262 230 263 
rect 229 270 230 271 
rect 229 273 230 274 
rect 229 276 230 277 
rect 229 278 230 279 
rect 229 293 230 294 
rect 229 302 230 303 
rect 229 305 230 306 
rect 229 307 230 308 
rect 230 1 231 2 
rect 230 3 231 4 
rect 230 8 231 9 
rect 230 18 231 19 
rect 230 21 231 22 
rect 230 23 231 24 
rect 230 30 231 31 
rect 230 40 231 41 
rect 230 43 231 44 
rect 230 66 231 67 
rect 230 68 231 69 
rect 230 71 231 72 
rect 230 95 231 96 
rect 230 97 231 98 
rect 230 100 231 101 
rect 230 101 231 102 
rect 230 112 231 113 
rect 230 114 231 115 
rect 230 118 231 119 
rect 230 120 231 121 
rect 230 121 231 122 
rect 230 122 231 123 
rect 230 123 231 124 
rect 230 124 231 125 
rect 230 125 231 126 
rect 230 126 231 127 
rect 230 127 231 128 
rect 230 128 231 129 
rect 230 129 231 130 
rect 230 130 231 131 
rect 230 131 231 132 
rect 230 132 231 133 
rect 230 133 231 134 
rect 230 134 231 135 
rect 230 135 231 136 
rect 230 136 231 137 
rect 230 137 231 138 
rect 230 138 231 139 
rect 230 139 231 140 
rect 230 140 231 141 
rect 230 141 231 142 
rect 230 142 231 143 
rect 230 143 231 144 
rect 230 144 231 145 
rect 230 145 231 146 
rect 230 146 231 147 
rect 230 147 231 148 
rect 230 148 231 149 
rect 230 149 231 150 
rect 230 150 231 151 
rect 230 151 231 152 
rect 230 152 231 153 
rect 230 153 231 154 
rect 230 154 231 155 
rect 230 155 231 156 
rect 230 156 231 157 
rect 230 157 231 158 
rect 230 158 231 159 
rect 230 159 231 160 
rect 230 160 231 161 
rect 230 161 231 162 
rect 230 162 231 163 
rect 230 163 231 164 
rect 230 164 231 165 
rect 230 165 231 166 
rect 230 166 231 167 
rect 230 167 231 168 
rect 230 168 231 169 
rect 230 169 231 170 
rect 230 170 231 171 
rect 230 171 231 172 
rect 230 172 231 173 
rect 230 173 231 174 
rect 230 174 231 175 
rect 230 175 231 176 
rect 230 176 231 177 
rect 230 177 231 178 
rect 230 178 231 179 
rect 230 179 231 180 
rect 230 180 231 181 
rect 230 181 231 182 
rect 230 182 231 183 
rect 230 183 231 184 
rect 230 187 231 188 
rect 230 227 231 228 
rect 230 229 231 230 
rect 230 232 231 233 
rect 230 242 231 243 
rect 230 262 231 263 
rect 230 270 231 271 
rect 230 273 231 274 
rect 230 276 231 277 
rect 230 278 231 279 
rect 230 293 231 294 
rect 230 302 231 303 
rect 230 305 231 306 
rect 230 307 231 308 
rect 231 1 232 2 
rect 231 3 232 4 
rect 231 8 232 9 
rect 231 18 232 19 
rect 231 21 232 22 
rect 231 23 232 24 
rect 231 30 232 31 
rect 231 39 232 40 
rect 231 40 232 41 
rect 231 43 232 44 
rect 231 66 232 67 
rect 231 68 232 69 
rect 231 71 232 72 
rect 231 95 232 96 
rect 231 97 232 98 
rect 231 114 232 115 
rect 231 118 232 119 
rect 231 215 232 216 
rect 231 216 232 217 
rect 231 217 232 218 
rect 231 218 232 219 
rect 231 219 232 220 
rect 231 220 232 221 
rect 231 221 232 222 
rect 231 222 232 223 
rect 231 227 232 228 
rect 231 229 232 230 
rect 231 232 232 233 
rect 231 242 232 243 
rect 231 262 232 263 
rect 231 270 232 271 
rect 231 273 232 274 
rect 231 276 232 277 
rect 231 278 232 279 
rect 231 293 232 294 
rect 231 302 232 303 
rect 231 305 232 306 
rect 231 307 232 308 
rect 232 1 233 2 
rect 232 3 233 4 
rect 232 8 233 9 
rect 232 18 233 19 
rect 232 21 233 22 
rect 232 23 233 24 
rect 232 30 233 31 
rect 232 38 233 39 
rect 232 39 233 40 
rect 232 41 233 42 
rect 232 42 233 43 
rect 232 43 233 44 
rect 232 66 233 67 
rect 232 68 233 69 
rect 232 71 233 72 
rect 232 72 233 73 
rect 232 73 233 74 
rect 232 74 233 75 
rect 232 75 233 76 
rect 232 76 233 77 
rect 232 77 233 78 
rect 232 78 233 79 
rect 232 79 233 80 
rect 232 80 233 81 
rect 232 91 233 92 
rect 232 92 233 93 
rect 232 93 233 94 
rect 232 95 233 96 
rect 232 97 233 98 
rect 232 105 233 106 
rect 232 106 233 107 
rect 232 107 233 108 
rect 232 108 233 109 
rect 232 109 233 110 
rect 232 110 233 111 
rect 232 111 233 112 
rect 232 112 233 113 
rect 232 113 233 114 
rect 232 114 233 115 
rect 232 118 233 119 
rect 232 119 233 120 
rect 232 120 233 121 
rect 232 121 233 122 
rect 232 122 233 123 
rect 232 123 233 124 
rect 232 124 233 125 
rect 232 125 233 126 
rect 232 126 233 127 
rect 232 127 233 128 
rect 232 128 233 129 
rect 232 129 233 130 
rect 232 130 233 131 
rect 232 131 233 132 
rect 232 132 233 133 
rect 232 133 233 134 
rect 232 134 233 135 
rect 232 135 233 136 
rect 232 136 233 137 
rect 232 137 233 138 
rect 232 138 233 139 
rect 232 139 233 140 
rect 232 140 233 141 
rect 232 141 233 142 
rect 232 142 233 143 
rect 232 143 233 144 
rect 232 144 233 145 
rect 232 145 233 146 
rect 232 146 233 147 
rect 232 147 233 148 
rect 232 148 233 149 
rect 232 149 233 150 
rect 232 150 233 151 
rect 232 151 233 152 
rect 232 152 233 153 
rect 232 153 233 154 
rect 232 154 233 155 
rect 232 155 233 156 
rect 232 156 233 157 
rect 232 157 233 158 
rect 232 158 233 159 
rect 232 159 233 160 
rect 232 160 233 161 
rect 232 161 233 162 
rect 232 162 233 163 
rect 232 163 233 164 
rect 232 164 233 165 
rect 232 165 233 166 
rect 232 166 233 167 
rect 232 167 233 168 
rect 232 168 233 169 
rect 232 169 233 170 
rect 232 170 233 171 
rect 232 171 233 172 
rect 232 172 233 173 
rect 232 173 233 174 
rect 232 174 233 175 
rect 232 175 233 176 
rect 232 176 233 177 
rect 232 177 233 178 
rect 232 178 233 179 
rect 232 179 233 180 
rect 232 180 233 181 
rect 232 181 233 182 
rect 232 182 233 183 
rect 232 183 233 184 
rect 232 184 233 185 
rect 232 185 233 186 
rect 232 186 233 187 
rect 232 187 233 188 
rect 232 188 233 189 
rect 232 189 233 190 
rect 232 190 233 191 
rect 232 191 233 192 
rect 232 192 233 193 
rect 232 203 233 204 
rect 232 204 233 205 
rect 232 205 233 206 
rect 232 206 233 207 
rect 232 207 233 208 
rect 232 208 233 209 
rect 232 215 233 216 
rect 232 227 233 228 
rect 232 229 233 230 
rect 232 232 233 233 
rect 232 242 233 243 
rect 232 249 233 250 
rect 232 250 233 251 
rect 232 251 233 252 
rect 232 262 233 263 
rect 232 270 233 271 
rect 232 273 233 274 
rect 232 276 233 277 
rect 232 278 233 279 
rect 232 281 233 282 
rect 232 282 233 283 
rect 232 283 233 284 
rect 232 284 233 285 
rect 232 285 233 286 
rect 232 286 233 287 
rect 232 293 233 294 
rect 232 302 233 303 
rect 232 305 233 306 
rect 232 307 233 308 
rect 233 1 234 2 
rect 233 3 234 4 
rect 233 8 234 9 
rect 233 18 234 19 
rect 233 21 234 22 
rect 233 23 234 24 
rect 233 30 234 31 
rect 233 38 234 39 
rect 233 40 234 41 
rect 233 41 234 42 
rect 233 66 234 67 
rect 233 68 234 69 
rect 233 80 234 81 
rect 233 81 234 82 
rect 233 91 234 92 
rect 233 97 234 98 
rect 233 104 234 105 
rect 233 105 234 106 
rect 233 116 234 117 
rect 233 117 234 118 
rect 233 192 234 193 
rect 233 193 234 194 
rect 233 203 234 204 
rect 233 208 234 209 
rect 233 209 234 210 
rect 233 215 234 216 
rect 233 227 234 228 
rect 233 229 234 230 
rect 233 232 234 233 
rect 233 242 234 243 
rect 233 248 234 249 
rect 233 249 234 250 
rect 233 251 234 252 
rect 233 262 234 263 
rect 233 270 234 271 
rect 233 273 234 274 
rect 233 276 234 277 
rect 233 278 234 279 
rect 233 280 234 281 
rect 233 281 234 282 
rect 233 286 234 287 
rect 233 293 234 294 
rect 233 302 234 303 
rect 233 305 234 306 
rect 233 307 234 308 
rect 234 1 235 2 
rect 234 3 235 4 
rect 234 8 235 9 
rect 234 18 235 19 
rect 234 21 235 22 
rect 234 23 235 24 
rect 234 30 235 31 
rect 234 38 235 39 
rect 234 40 235 41 
rect 234 66 235 67 
rect 234 68 235 69 
rect 234 81 235 82 
rect 234 91 235 92 
rect 234 97 235 98 
rect 234 104 235 105 
rect 234 117 235 118 
rect 234 118 235 119 
rect 234 119 235 120 
rect 234 193 235 194 
rect 234 203 235 204 
rect 234 209 235 210 
rect 234 215 235 216 
rect 234 227 235 228 
rect 234 229 235 230 
rect 234 232 235 233 
rect 234 242 235 243 
rect 234 244 235 245 
rect 234 245 235 246 
rect 234 246 235 247 
rect 234 247 235 248 
rect 234 248 235 249 
rect 234 251 235 252 
rect 234 262 235 263 
rect 234 270 235 271 
rect 234 273 235 274 
rect 234 276 235 277 
rect 234 278 235 279 
rect 234 280 235 281 
rect 234 286 235 287 
rect 234 289 235 290 
rect 234 290 235 291 
rect 234 291 235 292 
rect 234 292 235 293 
rect 234 293 235 294 
rect 234 302 235 303 
rect 234 305 235 306 
rect 234 307 235 308 
rect 235 1 236 2 
rect 235 3 236 4 
rect 235 8 236 9 
rect 235 18 236 19 
rect 235 21 236 22 
rect 235 23 236 24 
rect 235 38 236 39 
rect 235 40 236 41 
rect 235 66 236 67 
rect 235 68 236 69 
rect 235 81 236 82 
rect 235 82 236 83 
rect 235 83 236 84 
rect 235 84 236 85 
rect 235 85 236 86 
rect 235 86 236 87 
rect 235 87 236 88 
rect 235 97 236 98 
rect 235 100 236 101 
rect 235 101 236 102 
rect 235 102 236 103 
rect 235 103 236 104 
rect 235 104 236 105 
rect 235 119 236 120 
rect 235 193 236 194 
rect 235 194 236 195 
rect 235 209 236 210 
rect 235 215 236 216 
rect 235 227 236 228 
rect 235 229 236 230 
rect 235 232 236 233 
rect 235 242 236 243 
rect 235 244 236 245 
rect 235 262 236 263 
rect 235 273 236 274 
rect 235 276 236 277 
rect 235 278 236 279 
rect 235 280 236 281 
rect 235 289 236 290 
rect 235 305 236 306 
rect 235 307 236 308 
rect 236 1 237 2 
rect 236 3 237 4 
rect 236 8 237 9 
rect 236 18 237 19 
rect 236 21 237 22 
rect 236 23 237 24 
rect 236 38 237 39 
rect 236 40 237 41 
rect 236 66 237 67 
rect 236 68 237 69 
rect 236 87 237 88 
rect 236 97 237 98 
rect 236 100 237 101 
rect 236 119 237 120 
rect 236 194 237 195 
rect 236 209 237 210 
rect 236 215 237 216 
rect 236 227 237 228 
rect 236 229 237 230 
rect 236 232 237 233 
rect 236 242 237 243 
rect 236 244 237 245 
rect 236 262 237 263 
rect 236 273 237 274 
rect 236 276 237 277 
rect 236 278 237 279 
rect 236 280 237 281 
rect 236 289 237 290 
rect 236 305 237 306 
rect 236 307 237 308 
rect 237 1 238 2 
rect 237 3 238 4 
rect 237 8 238 9 
rect 237 18 238 19 
rect 237 21 238 22 
rect 237 23 238 24 
rect 237 38 238 39 
rect 237 40 238 41 
rect 237 66 238 67 
rect 237 68 238 69 
rect 237 87 238 88 
rect 237 97 238 98 
rect 237 100 238 101 
rect 237 119 238 120 
rect 237 194 238 195 
rect 237 209 238 210 
rect 237 215 238 216 
rect 237 227 238 228 
rect 237 229 238 230 
rect 237 232 238 233 
rect 237 242 238 243 
rect 237 244 238 245 
rect 237 262 238 263 
rect 237 273 238 274 
rect 237 276 238 277 
rect 237 278 238 279 
rect 237 280 238 281 
rect 237 289 238 290 
rect 237 305 238 306 
rect 237 307 238 308 
rect 238 1 239 2 
rect 238 3 239 4 
rect 238 8 239 9 
rect 238 18 239 19 
rect 238 21 239 22 
rect 238 23 239 24 
rect 238 38 239 39 
rect 238 40 239 41 
rect 238 66 239 67 
rect 238 68 239 69 
rect 238 87 239 88 
rect 238 97 239 98 
rect 238 100 239 101 
rect 238 119 239 120 
rect 238 194 239 195 
rect 238 209 239 210 
rect 238 215 239 216 
rect 238 227 239 228 
rect 238 229 239 230 
rect 238 232 239 233 
rect 238 242 239 243 
rect 238 262 239 263 
rect 238 273 239 274 
rect 238 276 239 277 
rect 238 278 239 279 
rect 238 280 239 281 
rect 238 289 239 290 
rect 238 305 239 306 
rect 238 307 239 308 
rect 239 1 240 2 
rect 239 3 240 4 
rect 239 8 240 9 
rect 239 14 240 15 
rect 239 18 240 19 
rect 239 19 240 20 
rect 239 21 240 22 
rect 239 23 240 24 
rect 239 24 240 25 
rect 239 38 240 39 
rect 239 40 240 41 
rect 239 66 240 67 
rect 239 68 240 69 
rect 239 87 240 88 
rect 239 97 240 98 
rect 239 100 240 101 
rect 239 119 240 120 
rect 239 120 240 121 
rect 239 187 240 188 
rect 239 194 240 195 
rect 239 209 240 210 
rect 239 211 240 212 
rect 239 212 240 213 
rect 239 213 240 214 
rect 239 214 240 215 
rect 239 215 240 216 
rect 239 225 240 226 
rect 239 226 240 227 
rect 239 227 240 228 
rect 239 229 240 230 
rect 239 230 240 231 
rect 239 232 240 233 
rect 239 242 240 243 
rect 239 243 240 244 
rect 239 244 240 245 
rect 239 245 240 246 
rect 239 246 240 247 
rect 239 247 240 248 
rect 239 248 240 249 
rect 239 262 240 263 
rect 239 273 240 274 
rect 239 276 240 277 
rect 239 278 240 279 
rect 239 280 240 281 
rect 239 289 240 290 
rect 239 305 240 306 
rect 239 307 240 308 
rect 240 3 241 4 
rect 240 8 241 9 
rect 240 14 241 15 
rect 240 19 241 20 
rect 240 21 241 22 
rect 240 22 241 23 
rect 240 24 241 25 
rect 240 25 241 26 
rect 240 187 241 188 
rect 240 194 241 195 
rect 240 224 241 225 
rect 240 225 241 226 
rect 240 230 241 231 
rect 240 232 241 233 
rect 240 248 241 249 
rect 240 249 241 250 
rect 240 262 241 263 
rect 240 273 241 274 
rect 240 276 241 277 
rect 240 278 241 279 
rect 240 280 241 281 
rect 240 288 241 289 
rect 240 289 241 290 
rect 240 305 241 306 
rect 240 307 241 308 
rect 241 3 242 4 
rect 241 8 242 9 
rect 241 11 242 12 
rect 241 12 242 13 
rect 241 13 242 14 
rect 241 14 242 15 
rect 241 19 242 20 
rect 241 20 242 21 
rect 241 22 242 23 
rect 241 23 242 24 
rect 241 25 242 26 
rect 241 26 242 27 
rect 241 27 242 28 
rect 241 28 242 29 
rect 241 29 242 30 
rect 241 30 242 31 
rect 241 31 242 32 
rect 241 32 242 33 
rect 241 33 242 34 
rect 241 34 242 35 
rect 241 35 242 36 
rect 241 36 242 37 
rect 241 37 242 38 
rect 241 38 242 39 
rect 241 39 242 40 
rect 241 40 242 41 
rect 241 41 242 42 
rect 241 42 242 43 
rect 241 43 242 44 
rect 241 44 242 45 
rect 241 45 242 46 
rect 241 46 242 47 
rect 241 47 242 48 
rect 241 48 242 49 
rect 241 49 242 50 
rect 241 50 242 51 
rect 241 51 242 52 
rect 241 52 242 53 
rect 241 53 242 54 
rect 241 54 242 55 
rect 241 55 242 56 
rect 241 56 242 57 
rect 241 57 242 58 
rect 241 58 242 59 
rect 241 59 242 60 
rect 241 60 242 61 
rect 241 61 242 62 
rect 241 62 242 63 
rect 241 63 242 64 
rect 241 64 242 65 
rect 241 65 242 66 
rect 241 66 242 67 
rect 241 67 242 68 
rect 241 68 242 69 
rect 241 69 242 70 
rect 241 70 242 71 
rect 241 71 242 72 
rect 241 72 242 73 
rect 241 73 242 74 
rect 241 74 242 75 
rect 241 75 242 76 
rect 241 76 242 77 
rect 241 77 242 78 
rect 241 78 242 79 
rect 241 79 242 80 
rect 241 80 242 81 
rect 241 81 242 82 
rect 241 82 242 83 
rect 241 83 242 84 
rect 241 84 242 85 
rect 241 85 242 86 
rect 241 86 242 87 
rect 241 87 242 88 
rect 241 88 242 89 
rect 241 89 242 90 
rect 241 90 242 91 
rect 241 91 242 92 
rect 241 92 242 93 
rect 241 93 242 94 
rect 241 94 242 95 
rect 241 95 242 96 
rect 241 96 242 97 
rect 241 97 242 98 
rect 241 98 242 99 
rect 241 99 242 100 
rect 241 100 242 101 
rect 241 101 242 102 
rect 241 102 242 103 
rect 241 103 242 104 
rect 241 104 242 105 
rect 241 105 242 106 
rect 241 106 242 107 
rect 241 107 242 108 
rect 241 108 242 109 
rect 241 109 242 110 
rect 241 110 242 111 
rect 241 111 242 112 
rect 241 112 242 113 
rect 241 113 242 114 
rect 241 114 242 115 
rect 241 115 242 116 
rect 241 116 242 117 
rect 241 117 242 118 
rect 241 118 242 119 
rect 241 119 242 120 
rect 241 120 242 121 
rect 241 121 242 122 
rect 241 122 242 123 
rect 241 123 242 124 
rect 241 124 242 125 
rect 241 125 242 126 
rect 241 126 242 127 
rect 241 127 242 128 
rect 241 128 242 129 
rect 241 129 242 130 
rect 241 130 242 131 
rect 241 131 242 132 
rect 241 132 242 133 
rect 241 133 242 134 
rect 241 134 242 135 
rect 241 135 242 136 
rect 241 136 242 137 
rect 241 137 242 138 
rect 241 138 242 139 
rect 241 139 242 140 
rect 241 140 242 141 
rect 241 141 242 142 
rect 241 142 242 143 
rect 241 143 242 144 
rect 241 144 242 145 
rect 241 145 242 146 
rect 241 146 242 147 
rect 241 147 242 148 
rect 241 148 242 149 
rect 241 149 242 150 
rect 241 150 242 151 
rect 241 151 242 152 
rect 241 152 242 153 
rect 241 153 242 154 
rect 241 154 242 155 
rect 241 155 242 156 
rect 241 156 242 157 
rect 241 157 242 158 
rect 241 158 242 159 
rect 241 159 242 160 
rect 241 160 242 161 
rect 241 161 242 162 
rect 241 162 242 163 
rect 241 163 242 164 
rect 241 164 242 165 
rect 241 165 242 166 
rect 241 166 242 167 
rect 241 167 242 168 
rect 241 168 242 169 
rect 241 169 242 170 
rect 241 170 242 171 
rect 241 171 242 172 
rect 241 172 242 173 
rect 241 173 242 174 
rect 241 174 242 175 
rect 241 175 242 176 
rect 241 176 242 177 
rect 241 177 242 178 
rect 241 178 242 179 
rect 241 179 242 180 
rect 241 180 242 181 
rect 241 181 242 182 
rect 241 182 242 183 
rect 241 183 242 184 
rect 241 184 242 185 
rect 241 187 242 188 
rect 241 194 242 195 
rect 241 198 242 199 
rect 241 199 242 200 
rect 241 200 242 201 
rect 241 201 242 202 
rect 241 202 242 203 
rect 241 203 242 204 
rect 241 204 242 205 
rect 241 205 242 206 
rect 241 206 242 207 
rect 241 207 242 208 
rect 241 208 242 209 
rect 241 209 242 210 
rect 241 210 242 211 
rect 241 211 242 212 
rect 241 212 242 213 
rect 241 213 242 214 
rect 241 214 242 215 
rect 241 215 242 216 
rect 241 216 242 217 
rect 241 217 242 218 
rect 241 218 242 219 
rect 241 219 242 220 
rect 241 220 242 221 
rect 241 221 242 222 
rect 241 222 242 223 
rect 241 223 242 224 
rect 241 224 242 225 
rect 241 230 242 231 
rect 241 232 242 233 
rect 241 235 242 236 
rect 241 236 242 237 
rect 241 237 242 238 
rect 241 238 242 239 
rect 241 239 242 240 
rect 241 240 242 241 
rect 241 241 242 242 
rect 241 242 242 243 
rect 241 243 242 244 
rect 241 244 242 245 
rect 241 245 242 246 
rect 241 246 242 247 
rect 241 247 242 248 
rect 241 249 242 250 
rect 241 250 242 251 
rect 241 251 242 252 
rect 241 252 242 253 
rect 241 253 242 254 
rect 241 254 242 255 
rect 241 255 242 256 
rect 241 256 242 257 
rect 241 257 242 258 
rect 241 258 242 259 
rect 241 259 242 260 
rect 241 260 242 261 
rect 241 262 242 263 
rect 241 265 242 266 
rect 241 266 242 267 
rect 241 267 242 268 
rect 241 268 242 269 
rect 241 273 242 274 
rect 241 276 242 277 
rect 241 278 242 279 
rect 241 280 242 281 
rect 241 282 242 283 
rect 241 283 242 284 
rect 241 284 242 285 
rect 241 285 242 286 
rect 241 286 242 287 
rect 241 287 242 288 
rect 241 288 242 289 
rect 241 301 242 302 
rect 241 302 242 303 
rect 241 305 242 306 
rect 242 3 243 4 
rect 242 8 243 9 
rect 242 20 243 21 
rect 242 21 243 22 
rect 242 23 243 24 
rect 242 24 243 25 
rect 242 184 243 185 
rect 242 194 243 195 
rect 242 198 243 199 
rect 242 230 243 231 
rect 242 232 243 233 
rect 242 247 243 248 
rect 242 248 243 249 
rect 242 262 243 263 
rect 242 268 243 269 
rect 242 273 243 274 
rect 242 276 243 277 
rect 242 278 243 279 
rect 242 280 243 281 
rect 242 282 243 283 
rect 242 289 243 290 
rect 242 290 243 291 
rect 242 291 243 292 
rect 242 292 243 293 
rect 242 293 243 294 
rect 242 294 243 295 
rect 242 295 243 296 
rect 242 296 243 297 
rect 242 297 243 298 
rect 242 298 243 299 
rect 242 299 243 300 
rect 242 300 243 301 
rect 242 301 243 302 
rect 242 305 243 306 
rect 243 3 244 4 
rect 243 8 244 9 
rect 243 21 244 22 
rect 243 22 244 23 
rect 243 24 244 25 
rect 243 25 244 26 
rect 243 26 244 27 
rect 243 27 244 28 
rect 243 28 244 29 
rect 243 29 244 30 
rect 243 30 244 31 
rect 243 31 244 32 
rect 243 32 244 33 
rect 243 41 244 42 
rect 243 67 244 68 
rect 243 68 244 69 
rect 243 69 244 70 
rect 243 70 244 71 
rect 243 71 244 72 
rect 243 72 244 73 
rect 243 73 244 74 
rect 243 74 244 75 
rect 243 75 244 76 
rect 243 76 244 77 
rect 243 77 244 78 
rect 243 78 244 79 
rect 243 79 244 80 
rect 243 80 244 81 
rect 243 81 244 82 
rect 243 82 244 83 
rect 243 83 244 84 
rect 243 84 244 85 
rect 243 85 244 86 
rect 243 86 244 87 
rect 243 87 244 88 
rect 243 88 244 89 
rect 243 94 244 95 
rect 243 95 244 96 
rect 243 96 244 97 
rect 243 102 244 103 
rect 243 103 244 104 
rect 243 104 244 105 
rect 243 105 244 106 
rect 243 106 244 107 
rect 243 107 244 108 
rect 243 108 244 109 
rect 243 109 244 110 
rect 243 110 244 111 
rect 243 111 244 112 
rect 243 112 244 113 
rect 243 113 244 114 
rect 243 114 244 115 
rect 243 115 244 116 
rect 243 116 244 117 
rect 243 117 244 118 
rect 243 118 244 119 
rect 243 119 244 120 
rect 243 120 244 121 
rect 243 121 244 122 
rect 243 122 244 123 
rect 243 123 244 124 
rect 243 124 244 125 
rect 243 125 244 126 
rect 243 126 244 127 
rect 243 127 244 128 
rect 243 128 244 129 
rect 243 129 244 130 
rect 243 130 244 131 
rect 243 131 244 132 
rect 243 132 244 133 
rect 243 133 244 134 
rect 243 134 244 135 
rect 243 135 244 136 
rect 243 136 244 137 
rect 243 137 244 138 
rect 243 138 244 139 
rect 243 139 244 140 
rect 243 140 244 141 
rect 243 141 244 142 
rect 243 142 244 143 
rect 243 143 244 144 
rect 243 144 244 145 
rect 243 145 244 146 
rect 243 146 244 147 
rect 243 147 244 148 
rect 243 148 244 149 
rect 243 149 244 150 
rect 243 150 244 151 
rect 243 151 244 152 
rect 243 152 244 153 
rect 243 153 244 154 
rect 243 154 244 155 
rect 243 155 244 156 
rect 243 156 244 157 
rect 243 157 244 158 
rect 243 158 244 159 
rect 243 159 244 160 
rect 243 160 244 161 
rect 243 161 244 162 
rect 243 162 244 163 
rect 243 163 244 164 
rect 243 164 244 165 
rect 243 165 244 166 
rect 243 166 244 167 
rect 243 167 244 168 
rect 243 168 244 169 
rect 243 169 244 170 
rect 243 170 244 171 
rect 243 171 244 172 
rect 243 172 244 173 
rect 243 173 244 174 
rect 243 174 244 175 
rect 243 175 244 176 
rect 243 176 244 177 
rect 243 177 244 178 
rect 243 184 244 185 
rect 243 194 244 195 
rect 243 198 244 199 
rect 243 230 244 231 
rect 243 232 244 233 
rect 243 258 244 259 
rect 243 262 244 263 
rect 243 268 244 269 
rect 243 273 244 274 
rect 243 276 244 277 
rect 243 278 244 279 
rect 243 280 244 281 
rect 243 282 244 283 
rect 243 284 244 285 
rect 243 285 244 286 
rect 243 286 244 287 
rect 243 287 244 288 
rect 243 288 244 289 
rect 243 289 244 290 
rect 243 305 244 306 
rect 244 3 245 4 
rect 244 8 245 9 
rect 244 22 245 23 
rect 244 23 245 24 
rect 244 32 245 33 
rect 244 35 245 36 
rect 244 36 245 37 
rect 244 37 245 38 
rect 244 38 245 39 
rect 244 39 245 40 
rect 244 41 245 42 
rect 244 44 245 45 
rect 244 45 245 46 
rect 244 46 245 47 
rect 244 47 245 48 
rect 244 48 245 49 
rect 244 49 245 50 
rect 244 50 245 51 
rect 244 51 245 52 
rect 244 52 245 53 
rect 244 53 245 54 
rect 244 54 245 55 
rect 244 55 245 56 
rect 244 56 245 57 
rect 244 57 245 58 
rect 244 58 245 59 
rect 244 59 245 60 
rect 244 60 245 61 
rect 244 61 245 62 
rect 244 62 245 63 
rect 244 63 245 64 
rect 244 64 245 65 
rect 244 65 245 66 
rect 244 88 245 89 
rect 244 94 245 95 
rect 244 177 245 178 
rect 244 184 245 185 
rect 244 194 245 195 
rect 244 198 245 199 
rect 244 206 245 207 
rect 244 207 245 208 
rect 244 208 245 209 
rect 244 209 245 210 
rect 244 210 245 211 
rect 244 211 245 212 
rect 244 212 245 213 
rect 244 213 245 214 
rect 244 214 245 215 
rect 244 215 245 216 
rect 244 216 245 217 
rect 244 217 245 218 
rect 244 218 245 219 
rect 244 219 245 220 
rect 244 220 245 221 
rect 244 221 245 222 
rect 244 222 245 223 
rect 244 223 245 224 
rect 244 224 245 225 
rect 244 225 245 226 
rect 244 226 245 227 
rect 244 227 245 228 
rect 244 230 245 231 
rect 244 232 245 233 
rect 244 234 245 235 
rect 244 235 245 236 
rect 244 236 245 237 
rect 244 237 245 238 
rect 244 238 245 239 
rect 244 239 245 240 
rect 244 240 245 241 
rect 244 241 245 242 
rect 244 242 245 243 
rect 244 243 245 244 
rect 244 244 245 245 
rect 244 245 245 246 
rect 244 246 245 247 
rect 244 247 245 248 
rect 244 248 245 249 
rect 244 249 245 250 
rect 244 250 245 251 
rect 244 251 245 252 
rect 244 252 245 253 
rect 244 253 245 254 
rect 244 254 245 255 
rect 244 255 245 256 
rect 244 258 245 259 
rect 244 262 245 263 
rect 244 268 245 269 
rect 244 273 245 274 
rect 244 276 245 277 
rect 244 278 245 279 
rect 244 280 245 281 
rect 244 282 245 283 
rect 244 284 245 285 
rect 244 305 245 306 
rect 245 3 246 4 
rect 245 8 246 9 
rect 245 23 246 24 
rect 245 24 246 25 
rect 245 25 246 26 
rect 245 26 246 27 
rect 245 27 246 28 
rect 245 28 246 29 
rect 245 29 246 30 
rect 245 30 246 31 
rect 245 32 246 33 
rect 245 39 246 40 
rect 245 41 246 42 
rect 245 44 246 45 
rect 245 65 246 66 
rect 245 88 246 89 
rect 245 94 246 95 
rect 245 96 246 97 
rect 245 101 246 102 
rect 245 102 246 103 
rect 245 103 246 104 
rect 245 104 246 105 
rect 245 105 246 106 
rect 245 106 246 107 
rect 245 107 246 108 
rect 245 108 246 109 
rect 245 109 246 110 
rect 245 110 246 111 
rect 245 111 246 112 
rect 245 112 246 113 
rect 245 113 246 114 
rect 245 114 246 115 
rect 245 115 246 116 
rect 245 116 246 117 
rect 245 117 246 118 
rect 245 118 246 119 
rect 245 119 246 120 
rect 245 120 246 121 
rect 245 121 246 122 
rect 245 122 246 123 
rect 245 123 246 124 
rect 245 124 246 125 
rect 245 125 246 126 
rect 245 126 246 127 
rect 245 127 246 128 
rect 245 128 246 129 
rect 245 129 246 130 
rect 245 130 246 131 
rect 245 131 246 132 
rect 245 132 246 133 
rect 245 133 246 134 
rect 245 134 246 135 
rect 245 135 246 136 
rect 245 136 246 137 
rect 245 137 246 138 
rect 245 138 246 139 
rect 245 139 246 140 
rect 245 140 246 141 
rect 245 141 246 142 
rect 245 142 246 143 
rect 245 143 246 144 
rect 245 144 246 145 
rect 245 145 246 146 
rect 245 146 246 147 
rect 245 147 246 148 
rect 245 148 246 149 
rect 245 149 246 150 
rect 245 150 246 151 
rect 245 151 246 152 
rect 245 152 246 153 
rect 245 153 246 154 
rect 245 154 246 155 
rect 245 155 246 156 
rect 245 156 246 157 
rect 245 157 246 158 
rect 245 158 246 159 
rect 245 159 246 160 
rect 245 160 246 161 
rect 245 161 246 162 
rect 245 162 246 163 
rect 245 163 246 164 
rect 245 164 246 165 
rect 245 165 246 166 
rect 245 166 246 167 
rect 245 167 246 168 
rect 245 177 246 178 
rect 245 184 246 185 
rect 245 194 246 195 
rect 245 198 246 199 
rect 245 206 246 207 
rect 245 230 246 231 
rect 245 232 246 233 
rect 245 255 246 256 
rect 245 258 246 259 
rect 245 262 246 263 
rect 245 268 246 269 
rect 245 273 246 274 
rect 245 276 246 277 
rect 245 278 246 279 
rect 245 280 246 281 
rect 245 282 246 283 
rect 245 284 246 285 
rect 245 305 246 306 
rect 246 3 247 4 
rect 246 8 247 9 
rect 246 32 247 33 
rect 246 41 247 42 
rect 246 65 247 66 
rect 246 88 247 89 
rect 246 94 247 95 
rect 246 96 247 97 
rect 246 101 247 102 
rect 246 177 247 178 
rect 246 184 247 185 
rect 246 194 247 195 
rect 246 198 247 199 
rect 246 206 247 207 
rect 246 210 247 211 
rect 246 230 247 231 
rect 246 232 247 233 
rect 246 258 247 259 
rect 246 262 247 263 
rect 246 268 247 269 
rect 246 273 247 274 
rect 246 276 247 277 
rect 246 278 247 279 
rect 246 280 247 281 
rect 246 283 247 284 
rect 246 284 247 285 
rect 246 305 247 306 
rect 247 3 248 4 
rect 247 8 248 9 
rect 247 41 248 42 
rect 247 86 248 87 
rect 247 88 248 89 
rect 247 94 248 95 
rect 247 96 248 97 
rect 247 177 248 178 
rect 247 178 248 179 
rect 247 179 248 180 
rect 247 180 248 181 
rect 247 184 248 185 
rect 247 194 248 195 
rect 247 198 248 199 
rect 247 206 248 207 
rect 247 210 248 211 
rect 247 230 248 231 
rect 247 232 248 233 
rect 247 258 248 259 
rect 247 262 248 263 
rect 247 268 248 269 
rect 247 273 248 274 
rect 247 276 248 277 
rect 247 278 248 279 
rect 247 280 248 281 
rect 247 282 248 283 
rect 247 283 248 284 
rect 247 305 248 306 
rect 248 3 249 4 
rect 248 8 249 9 
rect 248 14 249 15 
rect 248 15 249 16 
rect 248 16 249 17 
rect 248 17 249 18 
rect 248 18 249 19 
rect 248 19 249 20 
rect 248 20 249 21 
rect 248 21 249 22 
rect 248 22 249 23 
rect 248 23 249 24 
rect 248 24 249 25 
rect 248 25 249 26 
rect 248 26 249 27 
rect 248 27 249 28 
rect 248 28 249 29 
rect 248 29 249 30 
rect 248 30 249 31 
rect 248 31 249 32 
rect 248 32 249 33 
rect 248 33 249 34 
rect 248 34 249 35 
rect 248 35 249 36 
rect 248 36 249 37 
rect 248 37 249 38 
rect 248 38 249 39 
rect 248 39 249 40 
rect 248 41 249 42 
rect 248 44 249 45 
rect 248 45 249 46 
rect 248 46 249 47 
rect 248 47 249 48 
rect 248 48 249 49 
rect 248 49 249 50 
rect 248 57 249 58 
rect 248 58 249 59 
rect 248 59 249 60 
rect 248 60 249 61 
rect 248 61 249 62 
rect 248 62 249 63 
rect 248 63 249 64 
rect 248 64 249 65 
rect 248 65 249 66 
rect 248 66 249 67 
rect 248 67 249 68 
rect 248 68 249 69 
rect 248 69 249 70 
rect 248 70 249 71 
rect 248 71 249 72 
rect 248 72 249 73 
rect 248 73 249 74 
rect 248 74 249 75 
rect 248 75 249 76 
rect 248 76 249 77 
rect 248 77 249 78 
rect 248 78 249 79 
rect 248 79 249 80 
rect 248 80 249 81 
rect 248 81 249 82 
rect 248 82 249 83 
rect 248 83 249 84 
rect 248 84 249 85 
rect 248 85 249 86 
rect 248 86 249 87 
rect 248 88 249 89 
rect 248 91 249 92 
rect 248 92 249 93 
rect 248 93 249 94 
rect 248 94 249 95 
rect 248 96 249 97 
rect 248 97 249 98 
rect 248 98 249 99 
rect 248 99 249 100 
rect 248 100 249 101 
rect 248 101 249 102 
rect 248 102 249 103 
rect 248 103 249 104 
rect 248 104 249 105 
rect 248 105 249 106 
rect 248 106 249 107 
rect 248 107 249 108 
rect 248 108 249 109 
rect 248 109 249 110 
rect 248 110 249 111 
rect 248 111 249 112 
rect 248 112 249 113 
rect 248 113 249 114 
rect 248 114 249 115 
rect 248 115 249 116 
rect 248 116 249 117 
rect 248 117 249 118 
rect 248 118 249 119 
rect 248 119 249 120 
rect 248 120 249 121 
rect 248 121 249 122 
rect 248 122 249 123 
rect 248 123 249 124 
rect 248 124 249 125 
rect 248 125 249 126 
rect 248 126 249 127 
rect 248 127 249 128 
rect 248 128 249 129 
rect 248 129 249 130 
rect 248 130 249 131 
rect 248 131 249 132 
rect 248 132 249 133 
rect 248 133 249 134 
rect 248 134 249 135 
rect 248 135 249 136 
rect 248 136 249 137 
rect 248 137 249 138 
rect 248 138 249 139 
rect 248 139 249 140 
rect 248 140 249 141 
rect 248 141 249 142 
rect 248 142 249 143 
rect 248 143 249 144 
rect 248 144 249 145 
rect 248 145 249 146 
rect 248 146 249 147 
rect 248 147 249 148 
rect 248 148 249 149 
rect 248 149 249 150 
rect 248 150 249 151 
rect 248 151 249 152 
rect 248 152 249 153 
rect 248 153 249 154 
rect 248 154 249 155 
rect 248 155 249 156 
rect 248 156 249 157 
rect 248 157 249 158 
rect 248 158 249 159 
rect 248 159 249 160 
rect 248 160 249 161 
rect 248 168 249 169 
rect 248 169 249 170 
rect 248 170 249 171 
rect 248 171 249 172 
rect 248 172 249 173 
rect 248 173 249 174 
rect 248 174 249 175 
rect 248 175 249 176 
rect 248 176 249 177 
rect 248 184 249 185 
rect 248 186 249 187 
rect 248 187 249 188 
rect 248 194 249 195 
rect 248 198 249 199 
rect 248 203 249 204 
rect 248 204 249 205 
rect 248 205 249 206 
rect 248 206 249 207 
rect 248 210 249 211 
rect 248 227 249 228 
rect 248 230 249 231 
rect 248 232 249 233 
rect 248 234 249 235 
rect 248 235 249 236 
rect 248 236 249 237 
rect 248 237 249 238 
rect 248 238 249 239 
rect 248 239 249 240 
rect 248 240 249 241 
rect 248 241 249 242 
rect 248 242 249 243 
rect 248 243 249 244 
rect 248 244 249 245 
rect 248 245 249 246 
rect 248 246 249 247 
rect 248 247 249 248 
rect 248 248 249 249 
rect 248 249 249 250 
rect 248 250 249 251 
rect 248 251 249 252 
rect 248 252 249 253 
rect 248 253 249 254 
rect 248 254 249 255 
rect 248 255 249 256 
rect 248 258 249 259 
rect 248 262 249 263 
rect 248 268 249 269 
rect 248 269 249 270 
rect 248 270 249 271 
rect 248 273 249 274 
rect 248 276 249 277 
rect 248 278 249 279 
rect 248 280 249 281 
rect 248 282 249 283 
rect 248 305 249 306 
rect 249 3 250 4 
rect 249 8 250 9 
rect 249 14 250 15 
rect 249 40 250 41 
rect 249 41 250 42 
rect 249 49 250 50 
rect 249 50 250 51 
rect 249 51 250 52 
rect 249 52 250 53 
rect 249 53 250 54 
rect 249 54 250 55 
rect 249 55 250 56 
rect 249 56 250 57 
rect 249 57 250 58 
rect 249 88 250 89 
rect 249 91 250 92 
rect 249 160 250 161 
rect 249 161 250 162 
rect 249 162 250 163 
rect 249 163 250 164 
rect 249 164 250 165 
rect 249 165 250 166 
rect 249 166 250 167 
rect 249 167 250 168 
rect 249 168 250 169 
rect 249 176 250 177 
rect 249 177 250 178 
rect 249 178 250 179 
rect 249 179 250 180 
rect 249 180 250 181 
rect 249 181 250 182 
rect 249 182 250 183 
rect 249 184 250 185 
rect 249 187 250 188 
rect 249 194 250 195 
rect 249 198 250 199 
rect 249 203 250 204 
rect 249 210 250 211 
rect 249 226 250 227 
rect 249 227 250 228 
rect 249 230 250 231 
rect 249 232 250 233 
rect 249 258 250 259 
rect 249 262 250 263 
rect 249 270 250 271 
rect 249 273 250 274 
rect 249 276 250 277 
rect 249 278 250 279 
rect 249 280 250 281 
rect 249 305 250 306 
rect 250 3 251 4 
rect 250 8 251 9 
rect 250 14 251 15 
rect 250 34 251 35 
rect 250 35 251 36 
rect 250 38 251 39 
rect 250 40 251 41 
rect 250 83 251 84 
rect 250 84 251 85 
rect 250 85 251 86 
rect 250 88 251 89 
rect 250 91 251 92 
rect 250 145 251 146 
rect 250 146 251 147 
rect 250 147 251 148 
rect 250 184 251 185 
rect 250 187 251 188 
rect 250 194 251 195 
rect 250 198 251 199 
rect 250 203 251 204 
rect 250 210 251 211 
rect 250 226 251 227 
rect 250 230 251 231 
rect 250 232 251 233 
rect 250 258 251 259 
rect 250 262 251 263 
rect 250 270 251 271 
rect 250 273 251 274 
rect 250 276 251 277 
rect 250 278 251 279 
rect 250 280 251 281 
rect 250 305 251 306 
rect 251 3 252 4 
rect 251 8 252 9 
rect 251 35 252 36 
rect 251 36 252 37 
rect 251 38 252 39 
rect 251 40 252 41 
rect 251 49 252 50 
rect 251 50 252 51 
rect 251 51 252 52 
rect 251 52 252 53 
rect 251 53 252 54 
rect 251 56 252 57 
rect 251 85 252 86 
rect 251 88 252 89 
rect 251 145 252 146 
rect 251 184 252 185 
rect 251 194 252 195 
rect 251 198 252 199 
rect 251 210 252 211 
rect 251 226 252 227 
rect 251 230 252 231 
rect 251 232 252 233 
rect 251 258 252 259 
rect 251 262 252 263 
rect 251 273 252 274 
rect 251 276 252 277 
rect 251 278 252 279 
rect 251 280 252 281 
rect 251 305 252 306 
rect 252 3 253 4 
rect 252 8 253 9 
rect 252 36 253 37 
rect 252 38 253 39 
rect 252 40 253 41 
rect 252 49 253 50 
rect 252 56 253 57 
rect 252 85 253 86 
rect 252 88 253 89 
rect 252 145 253 146 
rect 252 165 253 166 
rect 252 184 253 185 
rect 252 194 253 195 
rect 252 198 253 199 
rect 252 210 253 211 
rect 252 226 253 227 
rect 252 230 253 231 
rect 252 232 253 233 
rect 252 258 253 259 
rect 252 262 253 263 
rect 252 273 253 274 
rect 252 276 253 277 
rect 252 278 253 279 
rect 252 280 253 281 
rect 252 305 253 306 
rect 253 3 254 4 
rect 253 8 254 9 
rect 253 36 254 37 
rect 253 38 254 39 
rect 253 40 254 41 
rect 253 49 254 50 
rect 253 56 254 57 
rect 253 85 254 86 
rect 253 88 254 89 
rect 253 145 254 146 
rect 253 165 254 166 
rect 253 184 254 185 
rect 253 194 254 195 
rect 253 198 254 199 
rect 253 210 254 211 
rect 253 226 254 227 
rect 253 230 254 231 
rect 253 232 254 233 
rect 253 258 254 259 
rect 253 262 254 263 
rect 253 273 254 274 
rect 253 276 254 277 
rect 253 278 254 279 
rect 253 280 254 281 
rect 253 305 254 306 
rect 254 3 255 4 
rect 254 8 255 9 
rect 254 36 255 37 
rect 254 38 255 39 
rect 254 40 255 41 
rect 254 49 255 50 
rect 254 56 255 57 
rect 254 85 255 86 
rect 254 88 255 89 
rect 254 145 255 146 
rect 254 165 255 166 
rect 254 184 255 185 
rect 254 194 255 195 
rect 254 198 255 199 
rect 254 210 255 211 
rect 254 230 255 231 
rect 254 232 255 233 
rect 254 258 255 259 
rect 254 262 255 263 
rect 254 273 255 274 
rect 254 276 255 277 
rect 254 278 255 279 
rect 254 280 255 281 
rect 254 305 255 306 
rect 255 3 256 4 
rect 255 8 256 9 
rect 255 36 256 37 
rect 255 38 256 39 
rect 255 40 256 41 
rect 255 49 256 50 
rect 255 56 256 57 
rect 255 85 256 86 
rect 255 88 256 89 
rect 255 145 256 146 
rect 255 165 256 166 
rect 255 171 256 172 
rect 255 184 256 185 
rect 255 194 256 195 
rect 255 198 256 199 
rect 255 209 256 210 
rect 255 210 256 211 
rect 255 230 256 231 
rect 255 232 256 233 
rect 255 258 256 259 
rect 255 262 256 263 
rect 255 267 256 268 
rect 255 273 256 274 
rect 255 276 256 277 
rect 255 278 256 279 
rect 255 280 256 281 
rect 255 305 256 306 
rect 256 3 257 4 
rect 256 8 257 9 
rect 256 36 257 37 
rect 256 38 257 39 
rect 256 40 257 41 
rect 256 48 257 49 
rect 256 49 257 50 
rect 256 56 257 57 
rect 256 57 257 58 
rect 256 85 257 86 
rect 256 88 257 89 
rect 256 89 257 90 
rect 256 115 257 116 
rect 256 116 257 117 
rect 256 117 257 118 
rect 256 118 257 119 
rect 256 119 257 120 
rect 256 120 257 121 
rect 256 145 257 146 
rect 256 165 257 166 
rect 256 171 257 172 
rect 256 184 257 185 
rect 256 185 257 186 
rect 256 194 257 195 
rect 256 230 257 231 
rect 256 232 257 233 
rect 256 233 257 234 
rect 256 241 257 242 
rect 256 242 257 243 
rect 256 243 257 244 
rect 256 244 257 245 
rect 256 245 257 246 
rect 256 246 257 247 
rect 256 247 257 248 
rect 256 248 257 249 
rect 256 249 257 250 
rect 256 258 257 259 
rect 256 262 257 263 
rect 256 267 257 268 
rect 256 273 257 274 
rect 256 276 257 277 
rect 256 278 257 279 
rect 256 280 257 281 
rect 256 305 257 306 
rect 257 3 258 4 
rect 257 4 258 5 
rect 257 5 258 6 
rect 257 6 258 7 
rect 257 8 258 9 
rect 257 36 258 37 
rect 257 38 258 39 
rect 257 40 258 41 
rect 257 43 258 44 
rect 257 44 258 45 
rect 257 45 258 46 
rect 257 46 258 47 
rect 257 47 258 48 
rect 257 48 258 49 
rect 257 57 258 58 
rect 257 58 258 59 
rect 257 59 258 60 
rect 257 60 258 61 
rect 257 61 258 62 
rect 257 62 258 63 
rect 257 63 258 64 
rect 257 64 258 65 
rect 257 65 258 66 
rect 257 66 258 67 
rect 257 67 258 68 
rect 257 68 258 69 
rect 257 69 258 70 
rect 257 70 258 71 
rect 257 71 258 72 
rect 257 72 258 73 
rect 257 73 258 74 
rect 257 74 258 75 
rect 257 75 258 76 
rect 257 76 258 77 
rect 257 77 258 78 
rect 257 78 258 79 
rect 257 79 258 80 
rect 257 80 258 81 
rect 257 81 258 82 
rect 257 82 258 83 
rect 257 85 258 86 
rect 257 87 258 88 
rect 257 89 258 90 
rect 257 90 258 91 
rect 257 91 258 92 
rect 257 92 258 93 
rect 257 93 258 94 
rect 257 94 258 95 
rect 257 95 258 96 
rect 257 96 258 97 
rect 257 97 258 98 
rect 257 98 258 99 
rect 257 124 258 125 
rect 257 125 258 126 
rect 257 126 258 127 
rect 257 127 258 128 
rect 257 128 258 129 
rect 257 129 258 130 
rect 257 130 258 131 
rect 257 131 258 132 
rect 257 132 258 133 
rect 257 133 258 134 
rect 257 134 258 135 
rect 257 135 258 136 
rect 257 136 258 137 
rect 257 145 258 146 
rect 257 165 258 166 
rect 257 171 258 172 
rect 257 172 258 173 
rect 257 173 258 174 
rect 257 174 258 175 
rect 257 175 258 176 
rect 257 176 258 177 
rect 257 185 258 186 
rect 257 186 258 187 
rect 257 187 258 188 
rect 257 190 258 191 
rect 257 191 258 192 
rect 257 192 258 193 
rect 257 194 258 195 
rect 257 197 258 198 
rect 257 198 258 199 
rect 257 199 258 200 
rect 257 200 258 201 
rect 257 201 258 202 
rect 257 202 258 203 
rect 257 203 258 204 
rect 257 204 258 205 
rect 257 205 258 206 
rect 257 206 258 207 
rect 257 207 258 208 
rect 257 208 258 209 
rect 257 209 258 210 
rect 257 210 258 211 
rect 257 211 258 212 
rect 257 212 258 213 
rect 257 213 258 214 
rect 257 214 258 215 
rect 257 215 258 216 
rect 257 216 258 217 
rect 257 217 258 218 
rect 257 218 258 219 
rect 257 219 258 220 
rect 257 220 258 221 
rect 257 221 258 222 
rect 257 222 258 223 
rect 257 223 258 224 
rect 257 224 258 225 
rect 257 225 258 226 
rect 257 226 258 227 
rect 257 227 258 228 
rect 257 228 258 229 
rect 257 230 258 231 
rect 257 231 258 232 
rect 257 233 258 234 
rect 257 234 258 235 
rect 257 235 258 236 
rect 257 238 258 239 
rect 257 239 258 240 
rect 257 240 258 241 
rect 257 241 258 242 
rect 257 249 258 250 
rect 257 250 258 251 
rect 257 251 258 252 
rect 257 252 258 253 
rect 257 253 258 254 
rect 257 254 258 255 
rect 257 258 258 259 
rect 257 262 258 263 
rect 257 265 258 266 
rect 257 266 258 267 
rect 257 267 258 268 
rect 257 273 258 274 
rect 257 276 258 277 
rect 257 278 258 279 
rect 257 280 258 281 
rect 257 305 258 306 
rect 258 8 259 9 
rect 258 10 259 11 
rect 258 36 259 37 
rect 258 38 259 39 
rect 258 40 259 41 
rect 258 43 259 44 
rect 258 85 259 86 
rect 258 87 259 88 
rect 258 88 259 89 
rect 258 98 259 99 
rect 258 99 259 100 
rect 258 100 259 101 
rect 258 101 259 102 
rect 258 102 259 103 
rect 258 103 259 104 
rect 258 104 259 105 
rect 258 105 259 106 
rect 258 106 259 107 
rect 258 107 259 108 
rect 258 108 259 109 
rect 258 109 259 110 
rect 258 110 259 111 
rect 258 111 259 112 
rect 258 112 259 113 
rect 258 113 259 114 
rect 258 114 259 115 
rect 258 115 259 116 
rect 258 116 259 117 
rect 258 117 259 118 
rect 258 118 259 119 
rect 258 119 259 120 
rect 258 120 259 121 
rect 258 121 259 122 
rect 258 122 259 123 
rect 258 123 259 124 
rect 258 136 259 137 
rect 258 145 259 146 
rect 258 165 259 166 
rect 258 176 259 177 
rect 258 187 259 188 
rect 258 190 259 191 
rect 258 194 259 195 
rect 258 197 259 198 
rect 258 231 259 232 
rect 258 232 259 233 
rect 258 235 259 236 
rect 258 243 259 244 
rect 258 254 259 255 
rect 258 258 259 259 
rect 258 262 259 263 
rect 258 273 259 274 
rect 258 276 259 277 
rect 258 278 259 279 
rect 258 280 259 281 
rect 258 305 259 306 
rect 259 8 260 9 
rect 259 10 260 11 
rect 259 36 260 37 
rect 259 38 260 39 
rect 259 40 260 41 
rect 259 43 260 44 
rect 259 85 260 86 
rect 259 88 260 89 
rect 259 89 260 90 
rect 259 95 260 96 
rect 259 96 260 97 
rect 259 97 260 98 
rect 259 123 260 124 
rect 259 136 260 137 
rect 259 142 260 143 
rect 259 145 260 146 
rect 259 147 260 148 
rect 259 148 260 149 
rect 259 149 260 150 
rect 259 150 260 151 
rect 259 151 260 152 
rect 259 152 260 153 
rect 259 153 260 154 
rect 259 154 260 155 
rect 259 155 260 156 
rect 259 156 260 157 
rect 259 157 260 158 
rect 259 158 260 159 
rect 259 159 260 160 
rect 259 160 260 161 
rect 259 161 260 162 
rect 259 162 260 163 
rect 259 165 260 166 
rect 259 167 260 168 
rect 259 168 260 169 
rect 259 169 260 170 
rect 259 170 260 171 
rect 259 171 260 172 
rect 259 172 260 173 
rect 259 173 260 174 
rect 259 174 260 175 
rect 259 176 260 177 
rect 259 187 260 188 
rect 259 190 260 191 
rect 259 194 260 195 
rect 259 198 260 199 
rect 259 199 260 200 
rect 259 200 260 201 
rect 259 201 260 202 
rect 259 202 260 203 
rect 259 203 260 204 
rect 259 204 260 205 
rect 259 205 260 206 
rect 259 206 260 207 
rect 259 207 260 208 
rect 259 208 260 209 
rect 259 209 260 210 
rect 259 210 260 211 
rect 259 223 260 224 
rect 259 224 260 225 
rect 259 225 260 226 
rect 259 232 260 233 
rect 259 235 260 236 
rect 259 243 260 244 
rect 259 254 260 255 
rect 259 258 260 259 
rect 259 262 260 263 
rect 259 273 260 274 
rect 259 276 260 277 
rect 259 278 260 279 
rect 259 280 260 281 
rect 259 305 260 306 
rect 260 8 261 9 
rect 260 10 261 11 
rect 260 38 261 39 
rect 260 40 261 41 
rect 260 43 261 44 
rect 260 45 261 46 
rect 260 47 261 48 
rect 260 48 261 49 
rect 260 49 261 50 
rect 260 50 261 51 
rect 260 51 261 52 
rect 260 52 261 53 
rect 260 53 261 54 
rect 260 54 261 55 
rect 260 55 261 56 
rect 260 56 261 57 
rect 260 57 261 58 
rect 260 58 261 59 
rect 260 59 261 60 
rect 260 60 261 61 
rect 260 61 261 62 
rect 260 62 261 63 
rect 260 63 261 64 
rect 260 64 261 65 
rect 260 65 261 66 
rect 260 66 261 67 
rect 260 67 261 68 
rect 260 68 261 69 
rect 260 69 261 70 
rect 260 70 261 71 
rect 260 71 261 72 
rect 260 72 261 73 
rect 260 73 261 74 
rect 260 74 261 75 
rect 260 75 261 76 
rect 260 76 261 77 
rect 260 77 261 78 
rect 260 78 261 79 
rect 260 79 261 80 
rect 260 80 261 81 
rect 260 81 261 82 
rect 260 82 261 83 
rect 260 85 261 86 
rect 260 89 261 90 
rect 260 97 261 98 
rect 260 114 261 115 
rect 260 123 261 124 
rect 260 129 261 130 
rect 260 130 261 131 
rect 260 131 261 132 
rect 260 132 261 133 
rect 260 133 261 134 
rect 260 134 261 135 
rect 260 136 261 137 
rect 260 137 261 138 
rect 260 138 261 139 
rect 260 139 261 140 
rect 260 140 261 141 
rect 260 141 261 142 
rect 260 142 261 143 
rect 260 145 261 146 
rect 260 165 261 166 
rect 260 174 261 175 
rect 260 176 261 177 
rect 260 184 261 185 
rect 260 187 261 188 
rect 260 190 261 191 
rect 260 194 261 195 
rect 260 196 261 197 
rect 260 197 261 198 
rect 260 198 261 199 
rect 260 217 261 218 
rect 260 218 261 219 
rect 260 219 261 220 
rect 260 220 261 221 
rect 260 221 261 222 
rect 260 222 261 223 
rect 260 223 261 224 
rect 260 230 261 231 
rect 260 232 261 233 
rect 260 235 261 236 
rect 260 243 261 244 
rect 260 254 261 255 
rect 260 258 261 259 
rect 260 262 261 263 
rect 260 273 261 274 
rect 260 276 261 277 
rect 260 278 261 279 
rect 260 280 261 281 
rect 260 305 261 306 
rect 261 8 262 9 
rect 261 10 262 11 
rect 261 38 262 39 
rect 261 40 262 41 
rect 261 43 262 44 
rect 261 45 262 46 
rect 261 47 262 48 
rect 261 82 262 83 
rect 261 85 262 86 
rect 261 89 262 90 
rect 261 90 262 91 
rect 261 91 262 92 
rect 261 92 262 93 
rect 261 93 262 94 
rect 261 94 262 95 
rect 261 95 262 96 
rect 261 97 262 98 
rect 261 114 262 115 
rect 261 116 262 117 
rect 261 117 262 118 
rect 261 118 262 119 
rect 261 119 262 120 
rect 261 120 262 121 
rect 261 123 262 124 
rect 261 134 262 135 
rect 261 135 262 136 
rect 261 145 262 146 
rect 261 147 262 148 
rect 261 148 262 149 
rect 261 149 262 150 
rect 261 150 262 151 
rect 261 151 262 152 
rect 261 152 262 153 
rect 261 153 262 154 
rect 261 154 262 155 
rect 261 155 262 156 
rect 261 156 262 157 
rect 261 157 262 158 
rect 261 158 262 159 
rect 261 159 262 160 
rect 261 160 262 161 
rect 261 161 262 162 
rect 261 162 262 163 
rect 261 163 262 164 
rect 261 165 262 166 
rect 261 174 262 175 
rect 261 176 262 177 
rect 261 177 262 178 
rect 261 178 262 179 
rect 261 179 262 180 
rect 261 180 262 181 
rect 261 181 262 182 
rect 261 182 262 183 
rect 261 183 262 184 
rect 261 184 262 185 
rect 261 187 262 188 
rect 261 190 262 191 
rect 261 194 262 195 
rect 261 196 262 197 
rect 261 199 262 200 
rect 261 200 262 201 
rect 261 201 262 202 
rect 261 202 262 203 
rect 261 203 262 204 
rect 261 204 262 205 
rect 261 205 262 206 
rect 261 206 262 207 
rect 261 207 262 208 
rect 261 208 262 209 
rect 261 209 262 210 
rect 261 210 262 211 
rect 261 211 262 212 
rect 261 212 262 213 
rect 261 213 262 214 
rect 261 214 262 215 
rect 261 215 262 216 
rect 261 216 262 217 
rect 261 217 262 218 
rect 261 230 262 231 
rect 261 232 262 233 
rect 261 235 262 236 
rect 261 243 262 244 
rect 261 254 262 255 
rect 261 258 262 259 
rect 261 262 262 263 
rect 261 273 262 274 
rect 261 276 262 277 
rect 261 278 262 279 
rect 261 280 262 281 
rect 261 305 262 306 
rect 262 8 263 9 
rect 262 10 263 11 
rect 262 36 263 37 
rect 262 38 263 39 
rect 262 40 263 41 
rect 262 43 263 44 
rect 262 45 263 46 
rect 262 66 263 67 
rect 262 67 263 68 
rect 262 68 263 69 
rect 262 69 263 70 
rect 262 85 263 86 
rect 262 95 263 96 
rect 262 97 263 98 
rect 262 111 263 112 
rect 262 114 263 115 
rect 262 116 263 117 
rect 262 123 263 124 
rect 262 135 263 136 
rect 262 136 263 137 
rect 262 137 263 138 
rect 262 138 263 139 
rect 262 139 263 140 
rect 262 140 263 141 
rect 262 141 263 142 
rect 262 142 263 143 
rect 262 143 263 144 
rect 262 145 263 146 
rect 262 165 263 166 
rect 262 174 263 175 
rect 262 175 263 176 
rect 262 187 263 188 
rect 262 190 263 191 
rect 262 194 263 195 
rect 262 196 263 197 
rect 262 198 263 199 
rect 262 199 263 200 
rect 262 230 263 231 
rect 262 232 263 233 
rect 262 235 263 236 
rect 262 243 263 244 
rect 262 254 263 255 
rect 262 258 263 259 
rect 262 262 263 263 
rect 262 273 263 274 
rect 262 276 263 277 
rect 262 278 263 279 
rect 262 280 263 281 
rect 262 305 263 306 
rect 263 8 264 9 
rect 263 10 264 11 
rect 263 36 264 37 
rect 263 38 264 39 
rect 263 40 264 41 
rect 263 43 264 44 
rect 263 45 264 46 
rect 263 69 264 70 
rect 263 85 264 86 
rect 263 97 264 98 
rect 263 99 264 100 
rect 263 100 264 101 
rect 263 101 264 102 
rect 263 102 264 103 
rect 263 103 264 104 
rect 263 104 264 105 
rect 263 105 264 106 
rect 263 106 264 107 
rect 263 107 264 108 
rect 263 108 264 109 
rect 263 109 264 110 
rect 263 110 264 111 
rect 263 111 264 112 
rect 263 114 264 115 
rect 263 116 264 117 
rect 263 123 264 124 
rect 263 143 264 144 
rect 263 145 264 146 
rect 263 165 264 166 
rect 263 175 264 176 
rect 263 176 264 177 
rect 263 177 264 178 
rect 263 178 264 179 
rect 263 179 264 180 
rect 263 180 264 181 
rect 263 181 264 182 
rect 263 182 264 183 
rect 263 183 264 184 
rect 263 184 264 185 
rect 263 185 264 186 
rect 263 187 264 188 
rect 263 190 264 191 
rect 263 194 264 195 
rect 263 197 264 198 
rect 263 198 264 199 
rect 263 230 264 231 
rect 263 232 264 233 
rect 263 235 264 236 
rect 263 243 264 244 
rect 263 254 264 255 
rect 263 258 264 259 
rect 263 262 264 263 
rect 263 273 264 274 
rect 263 276 264 277 
rect 263 278 264 279 
rect 263 280 264 281 
rect 263 305 264 306 
rect 264 8 265 9 
rect 264 10 265 11 
rect 264 11 265 12 
rect 264 36 265 37 
rect 264 38 265 39 
rect 264 40 265 41 
rect 264 43 265 44 
rect 264 45 265 46 
rect 264 46 265 47 
rect 264 69 265 70 
rect 264 70 265 71 
rect 264 71 265 72 
rect 264 72 265 73 
rect 264 73 265 74 
rect 264 74 265 75 
rect 264 75 265 76 
rect 264 76 265 77 
rect 264 77 265 78 
rect 264 78 265 79 
rect 264 79 265 80 
rect 264 80 265 81 
rect 264 81 265 82 
rect 264 82 265 83 
rect 264 83 265 84 
rect 264 85 265 86 
rect 264 88 265 89 
rect 264 89 265 90 
rect 264 90 265 91 
rect 264 91 265 92 
rect 264 97 265 98 
rect 264 114 265 115 
rect 264 116 265 117 
rect 264 123 265 124 
rect 264 145 265 146 
rect 264 147 265 148 
rect 264 165 265 166 
rect 264 166 265 167 
rect 264 167 265 168 
rect 264 187 265 188 
rect 264 190 265 191 
rect 264 194 265 195 
rect 264 196 265 197 
rect 264 197 265 198 
rect 264 199 265 200 
rect 264 200 265 201 
rect 264 203 265 204 
rect 264 204 265 205 
rect 264 205 265 206 
rect 264 206 265 207 
rect 264 207 265 208 
rect 264 208 265 209 
rect 264 209 265 210 
rect 264 210 265 211 
rect 264 211 265 212 
rect 264 212 265 213 
rect 264 213 265 214 
rect 264 214 265 215 
rect 264 215 265 216 
rect 264 216 265 217 
rect 264 217 265 218 
rect 264 218 265 219 
rect 264 219 265 220 
rect 264 220 265 221 
rect 264 221 265 222 
rect 264 222 265 223 
rect 264 223 265 224 
rect 264 224 265 225 
rect 264 225 265 226 
rect 264 226 265 227 
rect 264 227 265 228 
rect 264 228 265 229 
rect 264 230 265 231 
rect 264 232 265 233 
rect 264 235 265 236 
rect 264 238 265 239 
rect 264 239 265 240 
rect 264 240 265 241 
rect 264 243 265 244 
rect 264 254 265 255 
rect 264 258 265 259 
rect 264 262 265 263 
rect 264 273 265 274 
rect 264 276 265 277 
rect 264 278 265 279 
rect 264 280 265 281 
rect 264 283 265 284 
rect 264 284 265 285 
rect 264 285 265 286 
rect 264 286 265 287 
rect 264 287 265 288 
rect 264 288 265 289 
rect 264 289 265 290 
rect 264 290 265 291 
rect 264 291 265 292 
rect 264 292 265 293 
rect 264 293 265 294 
rect 264 294 265 295 
rect 264 295 265 296 
rect 264 296 265 297 
rect 264 297 265 298 
rect 264 298 265 299 
rect 264 299 265 300 
rect 264 305 265 306 
rect 265 8 266 9 
rect 265 11 266 12 
rect 265 36 266 37 
rect 265 38 266 39 
rect 265 40 266 41 
rect 265 43 266 44 
rect 265 46 266 47 
rect 265 85 266 86 
rect 265 91 266 92 
rect 265 97 266 98 
rect 265 114 266 115 
rect 265 116 266 117 
rect 265 123 266 124 
rect 265 145 266 146 
rect 265 147 266 148 
rect 265 167 266 168 
rect 265 187 266 188 
rect 265 190 266 191 
rect 265 194 266 195 
rect 265 199 266 200 
rect 265 203 266 204 
rect 265 230 266 231 
rect 265 232 266 233 
rect 265 235 266 236 
rect 265 238 266 239 
rect 265 240 266 241 
rect 265 241 266 242 
rect 265 243 266 244 
rect 265 245 266 246 
rect 265 254 266 255 
rect 265 258 266 259 
rect 265 262 266 263 
rect 265 273 266 274 
rect 265 276 266 277 
rect 265 278 266 279 
rect 265 280 266 281 
rect 265 283 266 284 
rect 265 299 266 300 
rect 265 305 266 306 
rect 266 8 267 9 
rect 266 11 267 12 
rect 266 36 267 37 
rect 266 38 267 39 
rect 266 40 267 41 
rect 266 43 267 44 
rect 266 46 267 47 
rect 266 85 267 86 
rect 266 91 267 92 
rect 266 97 267 98 
rect 266 114 267 115 
rect 266 116 267 117 
rect 266 123 267 124 
rect 266 145 267 146 
rect 266 147 267 148 
rect 266 167 267 168 
rect 266 187 267 188 
rect 266 190 267 191 
rect 266 194 267 195 
rect 266 199 267 200 
rect 266 203 267 204 
rect 266 230 267 231 
rect 266 232 267 233 
rect 266 235 267 236 
rect 266 238 267 239 
rect 266 241 267 242 
rect 266 243 267 244 
rect 266 245 267 246 
rect 266 254 267 255 
rect 266 258 267 259 
rect 266 262 267 263 
rect 266 273 267 274 
rect 266 276 267 277 
rect 266 278 267 279 
rect 266 280 267 281 
rect 266 283 267 284 
rect 266 299 267 300 
rect 266 305 267 306 
rect 267 8 268 9 
rect 267 36 268 37 
rect 267 38 268 39 
rect 267 40 268 41 
rect 267 85 268 86 
rect 267 97 268 98 
rect 267 114 268 115 
rect 267 145 268 146 
rect 267 147 268 148 
rect 267 167 268 168 
rect 267 194 268 195 
rect 267 199 268 200 
rect 267 230 268 231 
rect 267 232 268 233 
rect 267 241 268 242 
rect 267 243 268 244 
rect 267 245 268 246 
rect 267 258 268 259 
rect 267 262 268 263 
rect 267 273 268 274 
rect 267 276 268 277 
rect 267 278 268 279 
rect 267 280 268 281 
rect 267 305 268 306 
rect 268 8 269 9 
rect 268 36 269 37 
rect 268 38 269 39 
rect 268 40 269 41 
rect 268 85 269 86 
rect 268 97 269 98 
rect 268 98 269 99 
rect 268 99 269 100 
rect 268 100 269 101 
rect 268 101 269 102 
rect 268 102 269 103 
rect 268 103 269 104 
rect 268 104 269 105 
rect 268 114 269 115 
rect 268 115 269 116 
rect 268 116 269 117 
rect 268 117 269 118 
rect 268 118 269 119 
rect 268 119 269 120 
rect 268 145 269 146 
rect 268 147 269 148 
rect 268 148 269 149 
rect 268 149 269 150 
rect 268 150 269 151 
rect 268 151 269 152 
rect 268 152 269 153 
rect 268 167 269 168 
rect 268 194 269 195 
rect 268 198 269 199 
rect 268 199 269 200 
rect 268 225 269 226 
rect 268 226 269 227 
rect 268 227 269 228 
rect 268 228 269 229 
rect 268 229 269 230 
rect 268 230 269 231 
rect 268 232 269 233 
rect 268 241 269 242 
rect 268 243 269 244 
rect 268 245 269 246 
rect 268 246 269 247 
rect 268 258 269 259 
rect 268 262 269 263 
rect 268 273 269 274 
rect 268 275 269 276 
rect 268 276 269 277 
rect 268 278 269 279 
rect 268 280 269 281 
rect 268 305 269 306 
rect 269 8 270 9 
rect 269 36 270 37 
rect 269 38 270 39 
rect 269 40 270 41 
rect 269 85 270 86 
rect 269 104 270 105 
rect 269 119 270 120 
rect 269 145 270 146 
rect 269 152 270 153 
rect 269 167 270 168 
rect 269 194 270 195 
rect 269 198 270 199 
rect 269 225 270 226 
rect 269 232 270 233 
rect 269 241 270 242 
rect 269 243 270 244 
rect 269 246 270 247 
rect 269 258 270 259 
rect 269 262 270 263 
rect 269 273 270 274 
rect 269 275 270 276 
rect 269 277 270 278 
rect 269 278 270 279 
rect 269 280 270 281 
rect 269 305 270 306 
rect 270 8 271 9 
rect 270 36 271 37 
rect 270 38 271 39 
rect 270 40 271 41 
rect 270 85 271 86 
rect 270 104 271 105 
rect 270 119 271 120 
rect 270 145 271 146 
rect 270 152 271 153 
rect 270 167 271 168 
rect 270 194 271 195 
rect 270 198 271 199 
rect 270 225 271 226 
rect 270 232 271 233 
rect 270 241 271 242 
rect 270 243 271 244 
rect 270 246 271 247 
rect 270 258 271 259 
rect 270 262 271 263 
rect 270 273 271 274 
rect 270 275 271 276 
rect 270 277 271 278 
rect 270 279 271 280 
rect 270 280 271 281 
rect 270 305 271 306 
rect 271 8 272 9 
rect 271 36 272 37 
rect 271 38 272 39 
rect 271 40 272 41 
rect 271 85 272 86 
rect 271 104 272 105 
rect 271 119 272 120 
rect 271 145 272 146 
rect 271 152 272 153 
rect 271 158 272 159 
rect 271 167 272 168 
rect 271 171 272 172 
rect 271 174 272 175 
rect 271 194 272 195 
rect 271 198 272 199 
rect 271 225 272 226 
rect 271 232 272 233 
rect 271 241 272 242 
rect 271 243 272 244 
rect 271 246 272 247 
rect 271 258 272 259 
rect 271 262 272 263 
rect 271 273 272 274 
rect 271 275 272 276 
rect 271 277 272 278 
rect 271 279 272 280 
rect 271 305 272 306 
rect 272 8 273 9 
rect 272 36 273 37 
rect 272 38 273 39 
rect 272 40 273 41 
rect 272 144 273 145 
rect 272 145 273 146 
rect 272 152 273 153 
rect 272 153 273 154 
rect 272 158 273 159 
rect 272 167 273 168 
rect 272 171 273 172 
rect 272 174 273 175 
rect 272 194 273 195 
rect 272 224 273 225 
rect 272 225 273 226 
rect 272 232 273 233 
rect 272 233 273 234 
rect 272 262 273 263 
rect 272 273 273 274 
rect 272 275 273 276 
rect 272 277 273 278 
rect 272 279 273 280 
rect 272 305 273 306 
rect 273 8 274 9 
rect 273 36 274 37 
rect 273 38 274 39 
rect 273 40 274 41 
rect 273 49 274 50 
rect 273 50 274 51 
rect 273 51 274 52 
rect 273 52 274 53 
rect 273 53 274 54 
rect 273 54 274 55 
rect 273 55 274 56 
rect 273 56 274 57 
rect 273 57 274 58 
rect 273 58 274 59 
rect 273 59 274 60 
rect 273 60 274 61 
rect 273 61 274 62 
rect 273 62 274 63 
rect 273 63 274 64 
rect 273 64 274 65 
rect 273 65 274 66 
rect 273 66 274 67 
rect 273 67 274 68 
rect 273 68 274 69 
rect 273 69 274 70 
rect 273 70 274 71 
rect 273 71 274 72 
rect 273 72 274 73 
rect 273 73 274 74 
rect 273 74 274 75 
rect 273 75 274 76 
rect 273 76 274 77 
rect 273 77 274 78 
rect 273 78 274 79 
rect 273 79 274 80 
rect 273 80 274 81 
rect 273 81 274 82 
rect 273 82 274 83 
rect 273 83 274 84 
rect 273 84 274 85 
rect 273 85 274 86 
rect 273 86 274 87 
rect 273 87 274 88 
rect 273 88 274 89 
rect 273 89 274 90 
rect 273 90 274 91 
rect 273 91 274 92 
rect 273 92 274 93 
rect 273 93 274 94 
rect 273 94 274 95 
rect 273 95 274 96 
rect 273 96 274 97 
rect 273 97 274 98 
rect 273 98 274 99 
rect 273 99 274 100 
rect 273 100 274 101 
rect 273 101 274 102 
rect 273 102 274 103 
rect 273 103 274 104 
rect 273 104 274 105 
rect 273 105 274 106 
rect 273 106 274 107 
rect 273 107 274 108 
rect 273 108 274 109 
rect 273 109 274 110 
rect 273 110 274 111 
rect 273 111 274 112 
rect 273 112 274 113 
rect 273 113 274 114 
rect 273 114 274 115 
rect 273 115 274 116 
rect 273 116 274 117 
rect 273 117 274 118 
rect 273 118 274 119 
rect 273 119 274 120 
rect 273 120 274 121 
rect 273 121 274 122 
rect 273 122 274 123 
rect 273 123 274 124 
rect 273 124 274 125 
rect 273 125 274 126 
rect 273 126 274 127 
rect 273 127 274 128 
rect 273 128 274 129 
rect 273 129 274 130 
rect 273 130 274 131 
rect 273 131 274 132 
rect 273 132 274 133 
rect 273 133 274 134 
rect 273 134 274 135 
rect 273 135 274 136 
rect 273 136 274 137 
rect 273 137 274 138 
rect 273 138 274 139 
rect 273 139 274 140 
rect 273 140 274 141 
rect 273 141 274 142 
rect 273 142 274 143 
rect 273 143 274 144 
rect 273 144 274 145 
rect 273 153 274 154 
rect 273 154 274 155 
rect 273 155 274 156 
rect 273 156 274 157 
rect 273 158 274 159 
rect 273 159 274 160 
rect 273 160 274 161 
rect 273 161 274 162 
rect 273 162 274 163 
rect 273 163 274 164 
rect 273 164 274 165 
rect 273 166 274 167 
rect 273 167 274 168 
rect 273 171 274 172 
rect 273 174 274 175 
rect 273 175 274 176 
rect 273 176 274 177 
rect 273 177 274 178 
rect 273 178 274 179 
rect 273 179 274 180 
rect 273 180 274 181 
rect 273 181 274 182 
rect 273 182 274 183 
rect 273 183 274 184 
rect 273 184 274 185 
rect 273 190 274 191 
rect 273 191 274 192 
rect 273 194 274 195 
rect 273 196 274 197 
rect 273 197 274 198 
rect 273 198 274 199 
rect 273 199 274 200 
rect 273 200 274 201 
rect 273 201 274 202 
rect 273 202 274 203 
rect 273 203 274 204 
rect 273 204 274 205 
rect 273 205 274 206 
rect 273 206 274 207 
rect 273 207 274 208 
rect 273 208 274 209 
rect 273 209 274 210 
rect 273 210 274 211 
rect 273 211 274 212 
rect 273 212 274 213 
rect 273 213 274 214 
rect 273 214 274 215 
rect 273 215 274 216 
rect 273 216 274 217 
rect 273 217 274 218 
rect 273 218 274 219 
rect 273 219 274 220 
rect 273 220 274 221 
rect 273 221 274 222 
rect 273 222 274 223 
rect 273 223 274 224 
rect 273 224 274 225 
rect 273 233 274 234 
rect 273 234 274 235 
rect 273 235 274 236 
rect 273 236 274 237 
rect 273 237 274 238 
rect 273 238 274 239 
rect 273 239 274 240 
rect 273 240 274 241 
rect 273 241 274 242 
rect 273 242 274 243 
rect 273 243 274 244 
rect 273 244 274 245 
rect 273 245 274 246 
rect 273 246 274 247 
rect 273 247 274 248 
rect 273 248 274 249 
rect 273 249 274 250 
rect 273 250 274 251 
rect 273 251 274 252 
rect 273 252 274 253 
rect 273 253 274 254 
rect 273 254 274 255 
rect 273 255 274 256 
rect 273 256 274 257 
rect 273 257 274 258 
rect 273 258 274 259 
rect 273 259 274 260 
rect 273 260 274 261 
rect 273 262 274 263 
rect 273 265 274 266 
rect 273 266 274 267 
rect 273 267 274 268 
rect 273 268 274 269 
rect 273 273 274 274 
rect 273 275 274 276 
rect 273 277 274 278 
rect 273 279 274 280 
rect 273 305 274 306 
rect 274 8 275 9 
rect 274 36 275 37 
rect 274 38 275 39 
rect 274 40 275 41 
rect 274 49 275 50 
rect 274 156 275 157 
rect 274 157 275 158 
rect 274 164 275 165 
rect 274 166 275 167 
rect 274 171 275 172 
rect 274 184 275 185 
rect 274 185 275 186 
rect 274 186 275 187 
rect 274 187 275 188 
rect 274 188 275 189 
rect 274 189 275 190 
rect 274 190 275 191 
rect 274 194 275 195 
rect 274 262 275 263 
rect 274 268 275 269 
rect 274 273 275 274 
rect 274 275 275 276 
rect 274 277 275 278 
rect 274 279 275 280 
rect 274 305 275 306 
rect 275 8 276 9 
rect 275 36 276 37 
rect 275 38 276 39 
rect 275 40 276 41 
rect 275 49 276 50 
rect 275 69 276 70 
rect 275 70 276 71 
rect 275 71 276 72 
rect 275 72 276 73 
rect 275 86 276 87 
rect 275 87 276 88 
rect 275 88 276 89 
rect 275 89 276 90 
rect 275 90 276 91 
rect 275 91 276 92 
rect 275 92 276 93 
rect 275 93 276 94 
rect 275 94 276 95 
rect 275 95 276 96 
rect 275 96 276 97 
rect 275 97 276 98 
rect 275 98 276 99 
rect 275 99 276 100 
rect 275 100 276 101 
rect 275 101 276 102 
rect 275 102 276 103 
rect 275 105 276 106 
rect 275 106 276 107 
rect 275 107 276 108 
rect 275 108 276 109 
rect 275 109 276 110 
rect 275 110 276 111 
rect 275 111 276 112 
rect 275 112 276 113 
rect 275 113 276 114 
rect 275 114 276 115 
rect 275 115 276 116 
rect 275 116 276 117 
rect 275 117 276 118 
rect 275 118 276 119 
rect 275 119 276 120 
rect 275 120 276 121 
rect 275 121 276 122 
rect 275 122 276 123 
rect 275 123 276 124 
rect 275 124 276 125 
rect 275 125 276 126 
rect 275 126 276 127 
rect 275 127 276 128 
rect 275 128 276 129 
rect 275 129 276 130 
rect 275 130 276 131 
rect 275 131 276 132 
rect 275 132 276 133 
rect 275 133 276 134 
rect 275 134 276 135 
rect 275 135 276 136 
rect 275 136 276 137 
rect 275 157 276 158 
rect 275 158 276 159 
rect 275 159 276 160 
rect 275 160 276 161 
rect 275 161 276 162 
rect 275 162 276 163 
rect 275 164 276 165 
rect 275 166 276 167 
rect 275 171 276 172 
rect 275 174 276 175 
rect 275 175 276 176 
rect 275 176 276 177 
rect 275 177 276 178 
rect 275 178 276 179 
rect 275 179 276 180 
rect 275 180 276 181 
rect 275 181 276 182 
rect 275 182 276 183 
rect 275 194 276 195 
rect 275 262 276 263 
rect 275 268 276 269 
rect 275 273 276 274 
rect 275 275 276 276 
rect 275 277 276 278 
rect 275 279 276 280 
rect 275 305 276 306 
rect 276 8 277 9 
rect 276 36 277 37 
rect 276 38 277 39 
rect 276 40 277 41 
rect 276 49 277 50 
rect 276 72 277 73 
rect 276 102 277 103 
rect 276 103 277 104 
rect 276 136 277 137 
rect 276 162 277 163 
rect 276 166 277 167 
rect 276 171 277 172 
rect 276 174 277 175 
rect 276 184 277 185 
rect 276 185 277 186 
rect 276 186 277 187 
rect 276 187 277 188 
rect 276 188 277 189 
rect 276 189 277 190 
rect 276 190 277 191 
rect 276 191 277 192 
rect 276 192 277 193 
rect 276 194 277 195 
rect 276 258 277 259 
rect 276 262 277 263 
rect 276 268 277 269 
rect 276 273 277 274 
rect 276 275 277 276 
rect 276 277 277 278 
rect 276 279 277 280 
rect 276 305 277 306 
rect 277 8 278 9 
rect 277 36 278 37 
rect 277 38 278 39 
rect 277 40 278 41 
rect 277 49 278 50 
rect 277 72 278 73 
rect 277 103 278 104 
rect 277 104 278 105 
rect 277 105 278 106 
rect 277 106 278 107 
rect 277 107 278 108 
rect 277 108 278 109 
rect 277 109 278 110 
rect 277 110 278 111 
rect 277 111 278 112 
rect 277 112 278 113 
rect 277 113 278 114 
rect 277 114 278 115 
rect 277 115 278 116 
rect 277 116 278 117 
rect 277 117 278 118 
rect 277 118 278 119 
rect 277 119 278 120 
rect 277 120 278 121 
rect 277 121 278 122 
rect 277 122 278 123 
rect 277 123 278 124 
rect 277 124 278 125 
rect 277 125 278 126 
rect 277 126 278 127 
rect 277 127 278 128 
rect 277 128 278 129 
rect 277 129 278 130 
rect 277 130 278 131 
rect 277 131 278 132 
rect 277 132 278 133 
rect 277 133 278 134 
rect 277 134 278 135 
rect 277 136 278 137 
rect 277 166 278 167 
rect 277 171 278 172 
rect 277 174 278 175 
rect 277 176 278 177 
rect 277 177 278 178 
rect 277 178 278 179 
rect 277 179 278 180 
rect 277 180 278 181 
rect 277 181 278 182 
rect 277 182 278 183 
rect 277 183 278 184 
rect 277 184 278 185 
rect 277 194 278 195 
rect 277 199 278 200 
rect 277 200 278 201 
rect 277 201 278 202 
rect 277 202 278 203 
rect 277 203 278 204 
rect 277 204 278 205 
rect 277 205 278 206 
rect 277 206 278 207 
rect 277 207 278 208 
rect 277 208 278 209 
rect 277 209 278 210 
rect 277 210 278 211 
rect 277 211 278 212 
rect 277 212 278 213 
rect 277 213 278 214 
rect 277 214 278 215 
rect 277 215 278 216 
rect 277 216 278 217 
rect 277 217 278 218 
rect 277 218 278 219 
rect 277 219 278 220 
rect 277 220 278 221 
rect 277 221 278 222 
rect 277 222 278 223 
rect 277 223 278 224 
rect 277 224 278 225 
rect 277 225 278 226 
rect 277 226 278 227 
rect 277 227 278 228 
rect 277 228 278 229 
rect 277 229 278 230 
rect 277 230 278 231 
rect 277 231 278 232 
rect 277 232 278 233 
rect 277 233 278 234 
rect 277 234 278 235 
rect 277 235 278 236 
rect 277 236 278 237 
rect 277 237 278 238 
rect 277 238 278 239 
rect 277 239 278 240 
rect 277 240 278 241 
rect 277 241 278 242 
rect 277 242 278 243 
rect 277 243 278 244 
rect 277 244 278 245 
rect 277 245 278 246 
rect 277 246 278 247 
rect 277 247 278 248 
rect 277 248 278 249 
rect 277 249 278 250 
rect 277 250 278 251 
rect 277 251 278 252 
rect 277 252 278 253 
rect 277 253 278 254 
rect 277 254 278 255 
rect 277 255 278 256 
rect 277 256 278 257 
rect 277 258 278 259 
rect 277 262 278 263 
rect 277 268 278 269 
rect 277 273 278 274 
rect 277 275 278 276 
rect 277 277 278 278 
rect 277 279 278 280 
rect 277 305 278 306 
rect 278 8 279 9 
rect 278 36 279 37 
rect 278 38 279 39 
rect 278 40 279 41 
rect 278 49 279 50 
rect 278 72 279 73 
rect 278 134 279 135 
rect 278 136 279 137 
rect 278 139 279 140 
rect 278 140 279 141 
rect 278 141 279 142 
rect 278 142 279 143 
rect 278 143 279 144 
rect 278 144 279 145 
rect 278 145 279 146 
rect 278 146 279 147 
rect 278 147 279 148 
rect 278 148 279 149 
rect 278 149 279 150 
rect 278 150 279 151 
rect 278 151 279 152 
rect 278 152 279 153 
rect 278 153 279 154 
rect 278 154 279 155 
rect 278 155 279 156 
rect 278 156 279 157 
rect 278 157 279 158 
rect 278 158 279 159 
rect 278 159 279 160 
rect 278 160 279 161 
rect 278 161 279 162 
rect 278 162 279 163 
rect 278 163 279 164 
rect 278 164 279 165 
rect 278 165 279 166 
rect 278 166 279 167 
rect 278 171 279 172 
rect 278 174 279 175 
rect 278 194 279 195 
rect 278 258 279 259 
rect 278 262 279 263 
rect 278 268 279 269 
rect 278 273 279 274 
rect 278 275 279 276 
rect 278 277 279 278 
rect 278 279 279 280 
rect 278 281 279 282 
rect 278 282 279 283 
rect 278 283 279 284 
rect 278 284 279 285 
rect 278 285 279 286 
rect 278 286 279 287 
rect 278 305 279 306 
rect 279 8 280 9 
rect 279 36 280 37 
rect 279 38 280 39 
rect 279 40 280 41 
rect 279 49 280 50 
rect 279 72 280 73 
rect 279 107 280 108 
rect 279 108 280 109 
rect 279 109 280 110 
rect 279 110 280 111 
rect 279 111 280 112 
rect 279 112 280 113 
rect 279 113 280 114 
rect 279 114 280 115 
rect 279 118 280 119 
rect 279 134 280 135 
rect 279 136 280 137 
rect 279 139 280 140 
rect 279 171 280 172 
rect 279 174 280 175 
rect 279 194 280 195 
rect 279 258 280 259 
rect 279 259 280 260 
rect 279 262 280 263 
rect 279 268 280 269 
rect 279 273 280 274 
rect 279 275 280 276 
rect 279 277 280 278 
rect 279 279 280 280 
rect 279 286 280 287 
rect 279 305 280 306 
rect 280 8 281 9 
rect 280 36 281 37 
rect 280 38 281 39 
rect 280 40 281 41 
rect 280 49 281 50 
rect 280 72 281 73 
rect 280 107 281 108 
rect 280 118 281 119 
rect 280 134 281 135 
rect 280 136 281 137 
rect 280 139 281 140 
rect 280 142 281 143 
rect 280 143 281 144 
rect 280 144 281 145 
rect 280 158 281 159 
rect 280 159 281 160 
rect 280 160 281 161 
rect 280 169 281 170 
rect 280 170 281 171 
rect 280 171 281 172 
rect 280 174 281 175 
rect 280 194 281 195 
rect 280 195 281 196 
rect 280 196 281 197 
rect 280 197 281 198 
rect 280 198 281 199 
rect 280 199 281 200 
rect 280 200 281 201 
rect 280 201 281 202 
rect 280 202 281 203 
rect 280 203 281 204 
rect 280 204 281 205 
rect 280 205 281 206 
rect 280 206 281 207 
rect 280 207 281 208 
rect 280 208 281 209 
rect 280 209 281 210 
rect 280 210 281 211 
rect 280 211 281 212 
rect 280 212 281 213 
rect 280 213 281 214 
rect 280 214 281 215 
rect 280 215 281 216 
rect 280 216 281 217 
rect 280 217 281 218 
rect 280 218 281 219 
rect 280 219 281 220 
rect 280 220 281 221 
rect 280 221 281 222 
rect 280 222 281 223 
rect 280 223 281 224 
rect 280 224 281 225 
rect 280 225 281 226 
rect 280 226 281 227 
rect 280 227 281 228 
rect 280 228 281 229 
rect 280 229 281 230 
rect 280 230 281 231 
rect 280 231 281 232 
rect 280 232 281 233 
rect 280 233 281 234 
rect 280 234 281 235 
rect 280 235 281 236 
rect 280 236 281 237 
rect 280 237 281 238 
rect 280 238 281 239 
rect 280 239 281 240 
rect 280 240 281 241 
rect 280 241 281 242 
rect 280 242 281 243 
rect 280 243 281 244 
rect 280 244 281 245 
rect 280 245 281 246 
rect 280 246 281 247 
rect 280 247 281 248 
rect 280 248 281 249 
rect 280 249 281 250 
rect 280 250 281 251 
rect 280 251 281 252 
rect 280 252 281 253 
rect 280 253 281 254 
rect 280 254 281 255 
rect 280 255 281 256 
rect 280 256 281 257 
rect 280 259 281 260 
rect 280 262 281 263 
rect 280 268 281 269 
rect 280 269 281 270 
rect 280 270 281 271 
rect 280 273 281 274 
rect 280 275 281 276 
rect 280 277 281 278 
rect 280 279 281 280 
rect 280 286 281 287 
rect 280 305 281 306 
rect 281 8 282 9 
rect 281 36 282 37 
rect 281 38 282 39 
rect 281 40 282 41 
rect 281 49 282 50 
rect 281 72 282 73 
rect 281 107 282 108 
rect 281 118 282 119 
rect 281 134 282 135 
rect 281 136 282 137 
rect 281 139 282 140 
rect 281 142 282 143 
rect 281 144 282 145 
rect 281 145 282 146 
rect 281 152 282 153 
rect 281 158 282 159 
rect 281 160 282 161 
rect 281 161 282 162 
rect 281 162 282 163 
rect 281 163 282 164 
rect 281 164 282 165 
rect 281 165 282 166 
rect 281 168 282 169 
rect 281 169 282 170 
rect 281 174 282 175 
rect 281 256 282 257 
rect 281 257 282 258 
rect 281 259 282 260 
rect 281 262 282 263 
rect 281 270 282 271 
rect 281 273 282 274 
rect 281 275 282 276 
rect 281 278 282 279 
rect 281 279 282 280 
rect 281 286 282 287 
rect 281 305 282 306 
rect 282 8 283 9 
rect 282 36 283 37 
rect 282 38 283 39 
rect 282 40 283 41 
rect 282 49 283 50 
rect 282 72 283 73 
rect 282 107 283 108 
rect 282 118 283 119 
rect 282 134 283 135 
rect 282 136 283 137 
rect 282 139 283 140 
rect 282 142 283 143 
rect 282 145 283 146 
rect 282 146 283 147 
rect 282 147 283 148 
rect 282 152 283 153 
rect 282 158 283 159 
rect 282 165 283 166 
rect 282 166 283 167 
rect 282 168 283 169 
rect 282 174 283 175 
rect 282 230 283 231 
rect 282 231 283 232 
rect 282 246 283 247 
rect 282 247 283 248 
rect 282 257 283 258 
rect 282 259 283 260 
rect 282 262 283 263 
rect 282 270 283 271 
rect 282 273 283 274 
rect 282 275 283 276 
rect 282 277 283 278 
rect 282 278 283 279 
rect 282 286 283 287 
rect 282 305 283 306 
rect 283 8 284 9 
rect 283 36 284 37 
rect 283 38 284 39 
rect 283 40 284 41 
rect 283 49 284 50 
rect 283 72 284 73 
rect 283 118 284 119 
rect 283 134 284 135 
rect 283 136 284 137 
rect 283 147 284 148 
rect 283 152 284 153 
rect 283 166 284 167 
rect 283 168 284 169 
rect 283 225 284 226 
rect 283 226 284 227 
rect 283 227 284 228 
rect 283 228 284 229 
rect 283 229 284 230 
rect 283 230 284 231 
rect 283 241 284 242 
rect 283 242 284 243 
rect 283 243 284 244 
rect 283 244 284 245 
rect 283 245 284 246 
rect 283 246 284 247 
rect 283 257 284 258 
rect 283 259 284 260 
rect 283 262 284 263 
rect 283 273 284 274 
rect 283 275 284 276 
rect 283 277 284 278 
rect 283 305 284 306 
rect 284 8 285 9 
rect 284 36 285 37 
rect 284 38 285 39 
rect 284 40 285 41 
rect 284 49 285 50 
rect 284 72 285 73 
rect 284 118 285 119 
rect 284 134 285 135 
rect 284 136 285 137 
rect 284 147 285 148 
rect 284 152 285 153 
rect 284 166 285 167 
rect 284 168 285 169 
rect 284 225 285 226 
rect 284 241 285 242 
rect 284 248 285 249 
rect 284 257 285 258 
rect 284 259 285 260 
rect 284 262 285 263 
rect 284 273 285 274 
rect 284 275 285 276 
rect 284 277 285 278 
rect 284 305 285 306 
rect 285 8 286 9 
rect 285 36 286 37 
rect 285 38 286 39 
rect 285 40 286 41 
rect 285 49 286 50 
rect 285 72 286 73 
rect 285 118 286 119 
rect 285 134 286 135 
rect 285 136 286 137 
rect 285 147 286 148 
rect 285 152 286 153 
rect 285 166 286 167 
rect 285 168 286 169 
rect 285 241 286 242 
rect 285 248 286 249 
rect 285 257 286 258 
rect 285 259 286 260 
rect 285 262 286 263 
rect 285 273 286 274 
rect 285 275 286 276 
rect 285 277 286 278 
rect 285 305 286 306 
rect 286 8 287 9 
rect 286 36 287 37 
rect 286 38 287 39 
rect 286 40 287 41 
rect 286 49 287 50 
rect 286 72 287 73 
rect 286 113 287 114 
rect 286 114 287 115 
rect 286 115 287 116 
rect 286 116 287 117 
rect 286 117 287 118 
rect 286 118 287 119 
rect 286 134 287 135 
rect 286 136 287 137 
rect 286 147 287 148 
rect 286 152 287 153 
rect 286 166 287 167 
rect 286 168 287 169 
rect 286 241 287 242 
rect 286 248 287 249 
rect 286 257 287 258 
rect 286 259 287 260 
rect 286 262 287 263 
rect 286 273 287 274 
rect 286 275 287 276 
rect 286 277 287 278 
rect 286 305 287 306 
rect 287 8 288 9 
rect 287 14 288 15 
rect 287 36 288 37 
rect 287 38 288 39 
rect 287 40 288 41 
rect 287 49 288 50 
rect 287 72 288 73 
rect 287 113 288 114 
rect 287 134 288 135 
rect 287 136 288 137 
rect 287 147 288 148 
rect 287 152 288 153 
rect 287 158 288 159 
rect 287 168 288 169 
rect 287 241 288 242 
rect 287 248 288 249 
rect 287 251 288 252 
rect 287 257 288 258 
rect 287 273 288 274 
rect 287 275 288 276 
rect 287 277 288 278 
rect 287 305 288 306 
rect 288 8 289 9 
rect 288 9 289 10 
rect 288 14 289 15 
rect 288 32 289 33 
rect 288 33 289 34 
rect 288 34 289 35 
rect 288 35 289 36 
rect 288 36 289 37 
rect 288 38 289 39 
rect 288 40 289 41 
rect 288 41 289 42 
rect 288 48 289 49 
rect 288 49 289 50 
rect 288 72 289 73 
rect 288 73 289 74 
rect 288 112 289 113 
rect 288 113 289 114 
rect 288 134 289 135 
rect 288 136 289 137 
rect 288 137 289 138 
rect 288 147 289 148 
rect 288 152 289 153 
rect 288 153 289 154 
rect 288 158 289 159 
rect 288 240 289 241 
rect 288 241 289 242 
rect 288 248 289 249 
rect 288 249 289 250 
rect 288 251 289 252 
rect 288 257 289 258 
rect 288 258 289 259 
rect 288 259 289 260 
rect 288 260 289 261 
rect 288 261 289 262 
rect 288 262 289 263 
rect 288 263 289 264 
rect 288 264 289 265 
rect 288 272 289 273 
rect 288 273 289 274 
rect 288 275 289 276 
rect 288 277 289 278 
rect 288 305 289 306 
rect 289 9 290 10 
rect 289 10 290 11 
rect 289 11 290 12 
rect 289 12 290 13 
rect 289 13 290 14 
rect 289 14 290 15 
rect 289 27 290 28 
rect 289 28 290 29 
rect 289 29 290 30 
rect 289 30 290 31 
rect 289 31 290 32 
rect 289 32 290 33 
rect 289 38 290 39 
rect 289 41 290 42 
rect 289 42 290 43 
rect 289 43 290 44 
rect 289 45 290 46 
rect 289 46 290 47 
rect 289 47 290 48 
rect 289 48 290 49 
rect 289 73 290 74 
rect 289 74 290 75 
rect 289 75 290 76 
rect 289 76 290 77 
rect 289 77 290 78 
rect 289 78 290 79 
rect 289 79 290 80 
rect 289 80 290 81 
rect 289 107 290 108 
rect 289 108 290 109 
rect 289 109 290 110 
rect 289 110 290 111 
rect 289 111 290 112 
rect 289 112 290 113 
rect 289 134 290 135 
rect 289 135 290 136 
rect 289 137 290 138 
rect 289 138 290 139 
rect 289 139 290 140 
rect 289 140 290 141 
rect 289 141 290 142 
rect 289 142 290 143 
rect 289 143 290 144 
rect 289 144 290 145 
rect 289 145 290 146 
rect 289 147 290 148 
rect 289 153 290 154 
rect 289 154 290 155 
rect 289 155 290 156 
rect 289 156 290 157 
rect 289 157 290 158 
rect 289 158 290 159 
rect 289 160 290 161 
rect 289 161 290 162 
rect 289 162 290 163 
rect 289 163 290 164 
rect 289 164 290 165 
rect 289 165 290 166 
rect 289 166 290 167 
rect 289 167 290 168 
rect 289 168 290 169 
rect 289 169 290 170 
rect 289 170 290 171 
rect 289 171 290 172 
rect 289 172 290 173 
rect 289 173 290 174 
rect 289 174 290 175 
rect 289 175 290 176 
rect 289 176 290 177 
rect 289 177 290 178 
rect 289 178 290 179 
rect 289 179 290 180 
rect 289 180 290 181 
rect 289 181 290 182 
rect 289 182 290 183 
rect 289 183 290 184 
rect 289 184 290 185 
rect 289 185 290 186 
rect 289 186 290 187 
rect 289 187 290 188 
rect 289 188 290 189 
rect 289 189 290 190 
rect 289 190 290 191 
rect 289 191 290 192 
rect 289 192 290 193 
rect 289 193 290 194 
rect 289 194 290 195 
rect 289 195 290 196 
rect 289 196 290 197 
rect 289 197 290 198 
rect 289 198 290 199 
rect 289 199 290 200 
rect 289 200 290 201 
rect 289 201 290 202 
rect 289 202 290 203 
rect 289 203 290 204 
rect 289 204 290 205 
rect 289 205 290 206 
rect 289 206 290 207 
rect 289 207 290 208 
rect 289 208 290 209 
rect 289 209 290 210 
rect 289 210 290 211 
rect 289 211 290 212 
rect 289 212 290 213 
rect 289 213 290 214 
rect 289 214 290 215 
rect 289 215 290 216 
rect 289 216 290 217 
rect 289 217 290 218 
rect 289 218 290 219 
rect 289 219 290 220 
rect 289 220 290 221 
rect 289 221 290 222 
rect 289 222 290 223 
rect 289 223 290 224 
rect 289 224 290 225 
rect 289 225 290 226 
rect 289 226 290 227 
rect 289 227 290 228 
rect 289 228 290 229 
rect 289 229 290 230 
rect 289 230 290 231 
rect 289 231 290 232 
rect 289 232 290 233 
rect 289 233 290 234 
rect 289 234 290 235 
rect 289 235 290 236 
rect 289 236 290 237 
rect 289 237 290 238 
rect 289 238 290 239 
rect 289 239 290 240 
rect 289 240 290 241 
rect 289 249 290 250 
rect 289 250 290 251 
rect 289 251 290 252 
rect 289 264 290 265 
rect 289 270 290 271 
rect 289 271 290 272 
rect 289 272 290 273 
rect 289 274 290 275 
rect 289 275 290 276 
rect 289 277 290 278 
rect 289 305 290 306 
rect 290 27 291 28 
rect 290 38 291 39 
rect 290 43 291 44 
rect 290 45 291 46 
rect 290 80 291 81 
rect 290 107 291 108 
rect 290 123 291 124 
rect 290 135 291 136 
rect 290 136 291 137 
rect 290 145 291 146 
rect 290 147 291 148 
rect 290 148 291 149 
rect 290 149 291 150 
rect 290 150 291 151 
rect 290 151 291 152 
rect 290 152 291 153 
rect 290 159 291 160 
rect 290 160 291 161 
rect 290 264 291 265 
rect 290 270 291 271 
rect 290 274 291 275 
rect 290 305 291 306 
rect 291 27 292 28 
rect 291 38 292 39 
rect 291 43 292 44 
rect 291 45 292 46 
rect 291 80 292 81 
rect 291 107 292 108 
rect 291 123 292 124 
rect 291 136 292 137 
rect 291 137 292 138 
rect 291 138 292 139 
rect 291 139 292 140 
rect 291 140 292 141 
rect 291 141 292 142 
rect 291 142 292 143 
rect 291 145 292 146 
rect 291 146 292 147 
rect 291 152 292 153 
rect 291 153 292 154 
rect 291 154 292 155 
rect 291 155 292 156 
rect 291 156 292 157 
rect 291 157 292 158 
rect 291 158 292 159 
rect 291 159 292 160 
rect 291 161 292 162 
rect 291 162 292 163 
rect 291 163 292 164 
rect 291 164 292 165 
rect 291 165 292 166 
rect 291 166 292 167 
rect 291 167 292 168 
rect 291 168 292 169 
rect 291 169 292 170 
rect 291 170 292 171 
rect 291 171 292 172 
rect 291 172 292 173 
rect 291 173 292 174 
rect 291 174 292 175 
rect 291 175 292 176 
rect 291 176 292 177 
rect 291 177 292 178 
rect 291 178 292 179 
rect 291 179 292 180 
rect 291 180 292 181 
rect 291 181 292 182 
rect 291 182 292 183 
rect 291 183 292 184 
rect 291 184 292 185 
rect 291 185 292 186 
rect 291 186 292 187 
rect 291 187 292 188 
rect 291 188 292 189 
rect 291 189 292 190 
rect 291 190 292 191 
rect 291 191 292 192 
rect 291 192 292 193 
rect 291 193 292 194 
rect 291 194 292 195 
rect 291 195 292 196 
rect 291 196 292 197 
rect 291 197 292 198 
rect 291 198 292 199 
rect 291 199 292 200 
rect 291 200 292 201 
rect 291 201 292 202 
rect 291 202 292 203 
rect 291 203 292 204 
rect 291 204 292 205 
rect 291 205 292 206 
rect 291 206 292 207 
rect 291 207 292 208 
rect 291 208 292 209 
rect 291 209 292 210 
rect 291 210 292 211 
rect 291 211 292 212 
rect 291 212 292 213 
rect 291 213 292 214 
rect 291 214 292 215 
rect 291 215 292 216 
rect 291 216 292 217 
rect 291 217 292 218 
rect 291 218 292 219 
rect 291 219 292 220 
rect 291 220 292 221 
rect 291 221 292 222 
rect 291 222 292 223 
rect 291 223 292 224 
rect 291 224 292 225 
rect 291 225 292 226 
rect 291 226 292 227 
rect 291 227 292 228 
rect 291 228 292 229 
rect 291 229 292 230 
rect 291 230 292 231 
rect 291 231 292 232 
rect 291 232 292 233 
rect 291 233 292 234 
rect 291 234 292 235 
rect 291 235 292 236 
rect 291 236 292 237 
rect 291 237 292 238 
rect 291 238 292 239 
rect 291 239 292 240 
rect 291 240 292 241 
rect 291 241 292 242 
rect 291 242 292 243 
rect 291 243 292 244 
rect 291 244 292 245 
rect 291 245 292 246 
rect 291 246 292 247 
rect 291 247 292 248 
rect 291 248 292 249 
rect 291 249 292 250 
rect 291 250 292 251 
rect 291 251 292 252 
rect 291 252 292 253 
rect 291 253 292 254 
rect 291 254 292 255 
rect 291 255 292 256 
rect 291 256 292 257 
rect 291 257 292 258 
rect 291 258 292 259 
rect 291 259 292 260 
rect 291 260 292 261 
rect 291 262 292 263 
rect 291 264 292 265 
rect 291 270 292 271 
rect 291 274 292 275 
rect 291 305 292 306 
rect 292 27 293 28 
rect 292 38 293 39 
rect 292 41 293 42 
rect 292 43 293 44 
rect 292 80 293 81 
rect 292 107 293 108 
rect 292 123 293 124 
rect 292 142 293 143 
rect 292 146 293 147 
rect 292 147 293 148 
rect 292 148 293 149 
rect 292 160 293 161 
rect 292 161 293 162 
rect 292 262 293 263 
rect 292 264 293 265 
rect 292 270 293 271 
rect 292 305 293 306 
rect 293 27 294 28 
rect 293 38 294 39 
rect 293 40 294 41 
rect 293 41 294 42 
rect 293 43 294 44 
rect 293 80 294 81 
rect 293 107 294 108 
rect 293 123 294 124 
rect 293 142 294 143 
rect 293 148 294 149 
rect 293 149 294 150 
rect 293 150 294 151 
rect 293 151 294 152 
rect 293 152 294 153 
rect 293 153 294 154 
rect 293 154 294 155 
rect 293 155 294 156 
rect 293 156 294 157 
rect 293 157 294 158 
rect 293 158 294 159 
rect 293 160 294 161 
rect 293 169 294 170 
rect 293 170 294 171 
rect 293 171 294 172 
rect 293 172 294 173 
rect 293 173 294 174 
rect 293 174 294 175 
rect 293 175 294 176 
rect 293 176 294 177 
rect 293 178 294 179 
rect 293 179 294 180 
rect 293 180 294 181 
rect 293 181 294 182 
rect 293 182 294 183 
rect 293 183 294 184 
rect 293 184 294 185 
rect 293 185 294 186 
rect 293 186 294 187 
rect 293 187 294 188 
rect 293 188 294 189 
rect 293 189 294 190 
rect 293 190 294 191 
rect 293 191 294 192 
rect 293 192 294 193 
rect 293 193 294 194 
rect 293 194 294 195 
rect 293 195 294 196 
rect 293 196 294 197 
rect 293 197 294 198 
rect 293 198 294 199 
rect 293 199 294 200 
rect 293 200 294 201 
rect 293 201 294 202 
rect 293 202 294 203 
rect 293 203 294 204 
rect 293 204 294 205 
rect 293 205 294 206 
rect 293 206 294 207 
rect 293 207 294 208 
rect 293 208 294 209 
rect 293 209 294 210 
rect 293 210 294 211 
rect 293 211 294 212 
rect 293 212 294 213 
rect 293 213 294 214 
rect 293 214 294 215 
rect 293 215 294 216 
rect 293 216 294 217 
rect 293 217 294 218 
rect 293 218 294 219 
rect 293 219 294 220 
rect 293 220 294 221 
rect 293 221 294 222 
rect 293 222 294 223 
rect 293 223 294 224 
rect 293 224 294 225 
rect 293 262 294 263 
rect 293 264 294 265 
rect 293 265 294 266 
rect 293 266 294 267 
rect 293 267 294 268 
rect 293 270 294 271 
rect 293 272 294 273 
rect 293 273 294 274 
rect 293 274 294 275 
rect 293 275 294 276 
rect 293 276 294 277 
rect 293 277 294 278 
rect 293 278 294 279 
rect 293 279 294 280 
rect 293 280 294 281 
rect 293 281 294 282 
rect 293 282 294 283 
rect 293 283 294 284 
rect 293 284 294 285 
rect 293 285 294 286 
rect 293 286 294 287 
rect 293 287 294 288 
rect 293 288 294 289 
rect 293 289 294 290 
rect 293 290 294 291 
rect 293 291 294 292 
rect 293 292 294 293 
rect 293 293 294 294 
rect 293 294 294 295 
rect 293 295 294 296 
rect 293 296 294 297 
rect 293 297 294 298 
rect 293 298 294 299 
rect 293 299 294 300 
rect 293 300 294 301 
rect 293 301 294 302 
rect 293 302 294 303 
rect 293 305 294 306 
rect 294 27 295 28 
rect 294 38 295 39 
rect 294 40 295 41 
rect 294 43 295 44 
rect 294 80 295 81 
rect 294 107 295 108 
rect 294 123 295 124 
rect 294 142 295 143 
rect 294 158 295 159 
rect 294 176 295 177 
rect 294 262 295 263 
rect 294 270 295 271 
rect 294 302 295 303 
rect 294 305 295 306 
rect 295 27 296 28 
rect 295 38 296 39 
rect 295 40 296 41 
rect 295 43 296 44 
rect 295 80 296 81 
rect 295 107 296 108 
rect 295 123 296 124 
rect 295 142 296 143 
rect 295 155 296 156 
rect 295 158 296 159 
rect 295 176 296 177 
rect 295 262 296 263 
rect 295 270 296 271 
rect 295 302 296 303 
rect 295 305 296 306 
rect 296 27 297 28 
rect 296 30 297 31 
rect 296 31 297 32 
rect 296 32 297 33 
rect 296 40 297 41 
rect 296 43 297 44 
rect 296 80 297 81 
rect 296 107 297 108 
rect 296 123 297 124 
rect 296 142 297 143 
rect 296 155 297 156 
rect 296 158 297 159 
rect 296 176 297 177 
rect 296 185 297 186 
rect 296 186 297 187 
rect 296 187 297 188 
rect 296 188 297 189 
rect 296 189 297 190 
rect 296 190 297 191 
rect 296 191 297 192 
rect 296 192 297 193 
rect 296 201 297 202 
rect 296 202 297 203 
rect 296 203 297 204 
rect 296 204 297 205 
rect 296 205 297 206 
rect 296 206 297 207 
rect 296 207 297 208 
rect 296 208 297 209 
rect 296 217 297 218 
rect 296 218 297 219 
rect 296 219 297 220 
rect 296 220 297 221 
rect 296 221 297 222 
rect 296 222 297 223 
rect 296 223 297 224 
rect 296 224 297 225 
rect 296 233 297 234 
rect 296 234 297 235 
rect 296 235 297 236 
rect 296 236 297 237 
rect 296 237 297 238 
rect 296 238 297 239 
rect 296 239 297 240 
rect 296 240 297 241 
rect 296 249 297 250 
rect 296 250 297 251 
rect 296 251 297 252 
rect 296 252 297 253 
rect 296 253 297 254 
rect 296 254 297 255 
rect 296 262 297 263 
rect 296 267 297 268 
rect 296 268 297 269 
rect 296 270 297 271 
rect 296 302 297 303 
rect 296 305 297 306 
rect 297 27 298 28 
rect 297 30 298 31 
rect 297 32 298 33 
rect 297 33 298 34 
rect 297 34 298 35 
rect 297 35 298 36 
rect 297 36 298 37 
rect 297 37 298 38 
rect 297 38 298 39 
rect 297 39 298 40 
rect 297 40 298 41 
rect 297 43 298 44 
rect 297 80 298 81 
rect 297 81 298 82 
rect 297 82 298 83 
rect 297 83 298 84 
rect 297 84 298 85 
rect 297 85 298 86 
rect 297 86 298 87 
rect 297 87 298 88 
rect 297 88 298 89 
rect 297 107 298 108 
rect 297 123 298 124 
rect 297 142 298 143 
rect 297 155 298 156 
rect 297 158 298 159 
rect 297 176 298 177 
rect 297 177 298 178 
rect 297 178 298 179 
rect 297 179 298 180 
rect 297 180 298 181 
rect 297 181 298 182 
rect 297 182 298 183 
rect 297 183 298 184 
rect 297 184 298 185 
rect 297 185 298 186 
rect 297 192 298 193 
rect 297 193 298 194 
rect 297 194 298 195 
rect 297 195 298 196 
rect 297 196 298 197 
rect 297 197 298 198 
rect 297 198 298 199 
rect 297 199 298 200 
rect 297 200 298 201 
rect 297 201 298 202 
rect 297 208 298 209 
rect 297 209 298 210 
rect 297 210 298 211 
rect 297 211 298 212 
rect 297 212 298 213 
rect 297 213 298 214 
rect 297 214 298 215 
rect 297 215 298 216 
rect 297 216 298 217 
rect 297 217 298 218 
rect 297 224 298 225 
rect 297 225 298 226 
rect 297 226 298 227 
rect 297 227 298 228 
rect 297 228 298 229 
rect 297 229 298 230 
rect 297 230 298 231 
rect 297 231 298 232 
rect 297 232 298 233 
rect 297 233 298 234 
rect 297 240 298 241 
rect 297 241 298 242 
rect 297 242 298 243 
rect 297 243 298 244 
rect 297 244 298 245 
rect 297 245 298 246 
rect 297 246 298 247 
rect 297 247 298 248 
rect 297 248 298 249 
rect 297 249 298 250 
rect 297 254 298 255 
rect 297 257 298 258 
rect 297 258 298 259 
rect 297 259 298 260 
rect 297 260 298 261 
rect 297 261 298 262 
rect 297 262 298 263 
rect 297 267 298 268 
rect 297 270 298 271 
rect 297 302 298 303 
rect 297 305 298 306 
rect 298 27 299 28 
rect 298 30 299 31 
rect 298 43 299 44 
rect 298 88 299 89 
rect 298 107 299 108 
rect 298 123 299 124 
rect 298 142 299 143 
rect 298 155 299 156 
rect 298 158 299 159 
rect 298 254 299 255 
rect 298 257 299 258 
rect 298 267 299 268 
rect 298 270 299 271 
rect 298 302 299 303 
rect 298 305 299 306 
rect 299 39 300 40 
rect 299 40 300 41 
rect 299 88 300 89 
rect 299 257 300 258 
rect 299 260 300 261 
rect 299 305 300 306 
rect 300 40 301 41 
rect 300 88 301 89 
rect 300 257 301 258 
rect 300 260 301 261 
rect 300 305 301 306 
rect 301 40 302 41 
rect 301 88 302 89 
rect 301 257 302 258 
rect 301 260 302 261 
rect 301 305 302 306 
rect 302 40 303 41 
rect 302 88 303 89 
rect 302 257 303 258 
rect 302 260 303 261 
rect 302 305 303 306 
rect 303 30 304 31 
rect 303 40 304 41 
rect 303 43 304 44 
rect 303 88 304 89 
rect 303 94 304 95 
rect 303 123 304 124 
rect 303 257 304 258 
rect 303 260 304 261 
rect 303 267 304 268 
rect 303 270 304 271 
rect 303 305 304 306 
rect 304 30 305 31 
rect 304 40 305 41 
rect 304 41 305 42 
rect 304 43 305 44 
rect 304 88 305 89 
rect 304 89 305 90 
rect 304 94 305 95 
rect 304 123 305 124 
rect 304 256 305 257 
rect 304 257 305 258 
rect 304 260 305 261 
rect 304 261 305 262 
rect 304 262 305 263 
rect 304 263 305 264 
rect 304 264 305 265 
rect 304 265 305 266 
rect 304 267 305 268 
rect 304 270 305 271 
rect 304 304 305 305 
rect 304 305 305 306 
rect 305 30 306 31 
rect 305 31 306 32 
rect 305 32 306 33 
rect 305 33 306 34 
rect 305 34 306 35 
rect 305 35 306 36 
rect 305 36 306 37 
rect 305 37 306 38 
rect 305 38 306 39 
rect 305 39 306 40 
rect 305 41 306 42 
rect 305 42 306 43 
rect 305 43 306 44 
rect 305 89 306 90 
rect 305 90 306 91 
rect 305 91 306 92 
rect 305 92 306 93 
rect 305 93 306 94 
rect 305 94 306 95 
rect 305 123 306 124 
rect 305 124 306 125 
rect 305 125 306 126 
rect 305 126 306 127 
rect 305 127 306 128 
rect 305 128 306 129 
rect 305 129 306 130 
rect 305 130 306 131 
rect 305 131 306 132 
rect 305 132 306 133 
rect 305 133 306 134 
rect 305 134 306 135 
rect 305 135 306 136 
rect 305 136 306 137 
rect 305 137 306 138 
rect 305 138 306 139 
rect 305 139 306 140 
rect 305 140 306 141 
rect 305 141 306 142 
rect 305 142 306 143 
rect 305 143 306 144 
rect 305 144 306 145 
rect 305 145 306 146 
rect 305 146 306 147 
rect 305 147 306 148 
rect 305 148 306 149 
rect 305 149 306 150 
rect 305 150 306 151 
rect 305 151 306 152 
rect 305 152 306 153 
rect 305 153 306 154 
rect 305 154 306 155 
rect 305 155 306 156 
rect 305 156 306 157 
rect 305 157 306 158 
rect 305 158 306 159 
rect 305 159 306 160 
rect 305 160 306 161 
rect 305 161 306 162 
rect 305 162 306 163 
rect 305 163 306 164 
rect 305 164 306 165 
rect 305 165 306 166 
rect 305 166 306 167 
rect 305 167 306 168 
rect 305 168 306 169 
rect 305 169 306 170 
rect 305 170 306 171 
rect 305 171 306 172 
rect 305 172 306 173 
rect 305 173 306 174 
rect 305 174 306 175 
rect 305 175 306 176 
rect 305 176 306 177 
rect 305 177 306 178 
rect 305 178 306 179 
rect 305 179 306 180 
rect 305 180 306 181 
rect 305 181 306 182 
rect 305 182 306 183 
rect 305 183 306 184 
rect 305 184 306 185 
rect 305 185 306 186 
rect 305 186 306 187 
rect 305 187 306 188 
rect 305 188 306 189 
rect 305 189 306 190 
rect 305 190 306 191 
rect 305 191 306 192 
rect 305 192 306 193 
rect 305 193 306 194 
rect 305 194 306 195 
rect 305 195 306 196 
rect 305 196 306 197 
rect 305 197 306 198 
rect 305 198 306 199 
rect 305 199 306 200 
rect 305 200 306 201 
rect 305 201 306 202 
rect 305 202 306 203 
rect 305 203 306 204 
rect 305 204 306 205 
rect 305 205 306 206 
rect 305 206 306 207 
rect 305 207 306 208 
rect 305 208 306 209 
rect 305 209 306 210 
rect 305 210 306 211 
rect 305 211 306 212 
rect 305 212 306 213 
rect 305 213 306 214 
rect 305 214 306 215 
rect 305 215 306 216 
rect 305 216 306 217 
rect 305 217 306 218 
rect 305 218 306 219 
rect 305 219 306 220 
rect 305 220 306 221 
rect 305 221 306 222 
rect 305 222 306 223 
rect 305 223 306 224 
rect 305 224 306 225 
rect 305 225 306 226 
rect 305 226 306 227 
rect 305 227 306 228 
rect 305 228 306 229 
rect 305 229 306 230 
rect 305 230 306 231 
rect 305 231 306 232 
rect 305 232 306 233 
rect 305 233 306 234 
rect 305 234 306 235 
rect 305 235 306 236 
rect 305 236 306 237 
rect 305 237 306 238 
rect 305 238 306 239 
rect 305 239 306 240 
rect 305 240 306 241 
rect 305 241 306 242 
rect 305 242 306 243 
rect 305 243 306 244 
rect 305 244 306 245 
rect 305 245 306 246 
rect 305 246 306 247 
rect 305 247 306 248 
rect 305 248 306 249 
rect 305 249 306 250 
rect 305 250 306 251 
rect 305 251 306 252 
rect 305 252 306 253 
rect 305 253 306 254 
rect 305 254 306 255 
rect 305 255 306 256 
rect 305 256 306 257 
rect 305 265 306 266 
rect 305 266 306 267 
rect 305 267 306 268 
rect 305 270 306 271 
rect 305 271 306 272 
rect 305 272 306 273 
rect 305 273 306 274 
rect 305 274 306 275 
rect 305 275 306 276 
rect 305 276 306 277 
rect 305 277 306 278 
rect 305 278 306 279 
rect 305 279 306 280 
rect 305 280 306 281 
rect 305 281 306 282 
rect 305 282 306 283 
rect 305 283 306 284 
rect 305 284 306 285 
rect 305 285 306 286 
rect 305 286 306 287 
rect 305 287 306 288 
rect 305 288 306 289 
rect 305 289 306 290 
rect 305 290 306 291 
rect 305 291 306 292 
rect 305 292 306 293 
rect 305 293 306 294 
rect 305 294 306 295 
rect 305 295 306 296 
rect 305 296 306 297 
rect 305 297 306 298 
rect 305 298 306 299 
rect 305 299 306 300 
rect 305 300 306 301 
rect 305 301 306 302 
rect 305 302 306 303 
rect 305 303 306 304 
rect 305 304 306 305 
rect 306 39 307 40 
rect 306 40 307 41 
rect 307 40 308 41 
rect 307 41 308 42 
rect 307 42 308 43 
rect 307 43 308 44 
rect 307 44 308 45 
rect 307 45 308 46 
rect 307 46 308 47 
rect 307 47 308 48 
rect 307 48 308 49 
rect 307 49 308 50 
rect 307 50 308 51 
rect 307 51 308 52 
rect 307 52 308 53 
rect 307 53 308 54 
rect 307 54 308 55 
rect 307 55 308 56 
rect 307 56 308 57 
rect 307 57 308 58 
rect 307 58 308 59 
rect 307 59 308 60 
rect 307 60 308 61 
rect 307 61 308 62 
rect 307 62 308 63 
rect 307 63 308 64 
rect 307 64 308 65 
rect 307 65 308 66 
rect 307 66 308 67 
rect 307 67 308 68 
rect 307 68 308 69 
rect 307 69 308 70 
rect 307 70 308 71 
rect 307 71 308 72 
rect 307 72 308 73 
rect 307 73 308 74 
rect 307 74 308 75 
rect 307 75 308 76 
rect 307 76 308 77 
rect 307 77 308 78 
rect 307 78 308 79 
rect 307 79 308 80 
rect 307 80 308 81 
rect 307 81 308 82 
rect 307 82 308 83 
rect 307 83 308 84 
rect 307 84 308 85 
rect 307 85 308 86 
rect 307 86 308 87 
rect 307 87 308 88 
rect 307 88 308 89 
rect 307 89 308 90 
rect 307 90 308 91 
rect 307 91 308 92 
rect 307 92 308 93 
rect 307 93 308 94 
rect 307 94 308 95 
rect 307 95 308 96 
rect 307 96 308 97 
rect 307 97 308 98 
rect 307 98 308 99 
rect 307 99 308 100 
rect 307 100 308 101 
rect 307 101 308 102 
rect 307 102 308 103 
rect 307 103 308 104 
rect 307 104 308 105 
rect 307 105 308 106 
rect 307 106 308 107 
rect 307 107 308 108 
rect 307 108 308 109 
rect 307 109 308 110 
rect 307 110 308 111 
rect 307 111 308 112 
rect 307 112 308 113 
rect 307 113 308 114 
rect 307 114 308 115 
rect 307 115 308 116 
rect 307 116 308 117 
rect 307 117 308 118 
rect 307 118 308 119 
rect 307 119 308 120 
rect 307 120 308 121 
rect 307 121 308 122 
rect 307 122 308 123 
rect 307 123 308 124 
rect 307 124 308 125 
rect 307 125 308 126 
rect 307 126 308 127 
rect 307 127 308 128 
rect 307 128 308 129 
rect 307 129 308 130 
rect 307 130 308 131 
rect 307 131 308 132 
rect 307 132 308 133 
rect 307 133 308 134 
rect 307 134 308 135 
rect 307 135 308 136 
rect 307 136 308 137 
rect 307 137 308 138 
rect 307 138 308 139 
rect 307 139 308 140 
rect 307 140 308 141 
rect 307 141 308 142 
rect 307 142 308 143 
rect 307 143 308 144 
rect 307 144 308 145 
rect 307 145 308 146 
rect 307 146 308 147 
rect 307 147 308 148 
rect 307 148 308 149 
rect 307 149 308 150 
rect 307 150 308 151 
rect 307 151 308 152 
rect 307 152 308 153 
rect 307 153 308 154 
rect 307 154 308 155 
rect 307 155 308 156 
rect 307 156 308 157 
rect 307 157 308 158 
rect 307 158 308 159 
rect 307 159 308 160 
rect 307 160 308 161 
rect 307 161 308 162 
rect 307 162 308 163 
rect 307 163 308 164 
rect 307 164 308 165 
rect 307 165 308 166 
rect 307 166 308 167 
rect 307 167 308 168 
rect 307 168 308 169 
rect 307 169 308 170 
rect 307 170 308 171 
rect 307 171 308 172 
rect 307 172 308 173 
rect 307 173 308 174 
rect 307 174 308 175 
rect 307 175 308 176 
rect 307 176 308 177 
rect 307 177 308 178 
rect 307 178 308 179 
rect 307 179 308 180 
rect 307 180 308 181 
rect 307 181 308 182 
rect 307 182 308 183 
rect 307 183 308 184 
rect 307 184 308 185 
rect 307 185 308 186 
rect 307 186 308 187 
rect 307 187 308 188 
rect 307 188 308 189 
rect 307 189 308 190 
rect 307 190 308 191 
rect 307 191 308 192 
rect 307 192 308 193 
rect 307 193 308 194 
rect 307 194 308 195 
rect 307 195 308 196 
rect 307 196 308 197 
rect 307 197 308 198 
rect 307 198 308 199 
rect 307 199 308 200 
rect 307 200 308 201 
rect 307 201 308 202 
rect 307 202 308 203 
rect 307 203 308 204 
rect 307 204 308 205 
rect 307 205 308 206 
rect 307 206 308 207 
rect 307 207 308 208 
rect 307 208 308 209 
rect 307 209 308 210 
rect 307 210 308 211 
rect 307 211 308 212 
rect 307 212 308 213 
rect 307 213 308 214 
rect 307 214 308 215 
rect 307 215 308 216 
rect 307 216 308 217 
rect 307 217 308 218 
rect 307 218 308 219 
rect 307 219 308 220 
rect 307 220 308 221 
rect 307 239 308 240 
rect 307 240 308 241 
rect 307 241 308 242 
rect 307 242 308 243 
rect 308 220 309 221 
rect 308 221 309 222 
rect 308 222 309 223 
rect 308 223 309 224 
rect 308 224 309 225 
rect 308 225 309 226 
rect 308 226 309 227 
rect 308 227 309 228 
rect 308 228 309 229 
rect 308 229 309 230 
rect 308 230 309 231 
rect 308 231 309 232 
rect 308 232 309 233 
rect 308 233 309 234 
rect 308 234 309 235 
rect 308 235 309 236 
rect 308 236 309 237 
rect 308 237 309 238 
rect 308 238 309 239 
rect 308 239 309 240 
<< metal2 >>
rect 2 134 3 135 
rect 2 135 3 136 
rect 2 136 3 137 
rect 3 136 4 137 
rect 4 136 5 137 
rect 5 136 6 137 
rect 6 136 7 137 
rect 7 136 8 137 
rect 8 136 9 137 
rect 8 137 9 138 
rect 8 138 9 139 
rect 8 139 9 140 
rect 8 140 9 141 
rect 8 141 9 142 
rect 8 142 9 143 
rect 8 143 9 144 
rect 8 144 9 145 
rect 8 145 9 146 
rect 8 146 9 147 
rect 8 147 9 148 
rect 8 148 9 149 
rect 8 149 9 150 
rect 8 150 9 151 
rect 8 151 9 152 
rect 8 152 9 153 
rect 8 153 9 154 
rect 8 154 9 155 
rect 8 155 9 156 
rect 8 156 9 157 
rect 8 157 9 158 
rect 8 158 9 159 
rect 8 159 9 160 
rect 8 160 9 161 
rect 8 161 9 162 
rect 8 162 9 163 
rect 8 163 9 164 
rect 8 164 9 165 
rect 8 165 9 166 
rect 8 166 9 167 
rect 8 167 9 168 
rect 8 168 9 169 
rect 8 169 9 170 
rect 8 170 9 171 
rect 8 171 9 172 
rect 8 172 9 173 
rect 8 173 9 174 
rect 8 174 9 175 
rect 8 175 9 176 
rect 8 176 9 177 
rect 8 177 9 178 
rect 8 178 9 179 
rect 8 179 9 180 
rect 8 180 9 181 
rect 8 181 9 182 
rect 8 182 9 183 
rect 8 183 9 184 
rect 8 184 9 185 
rect 8 185 9 186 
rect 8 186 9 187 
rect 8 187 9 188 
rect 8 188 9 189 
rect 8 189 9 190 
rect 8 190 9 191 
rect 8 191 9 192 
rect 8 192 9 193 
rect 8 193 9 194 
rect 8 194 9 195 
rect 8 195 9 196 
rect 8 196 9 197 
rect 8 197 9 198 
rect 8 198 9 199 
rect 8 199 9 200 
rect 8 200 9 201 
rect 8 201 9 202 
rect 8 202 9 203 
rect 8 203 9 204 
rect 8 204 9 205 
rect 17 160 18 161 
rect 17 161 18 162 
rect 17 162 18 163 
rect 17 163 18 164 
rect 17 164 18 165 
rect 17 165 18 166 
rect 17 166 18 167 
rect 17 215 18 216 
rect 17 216 18 217 
rect 17 217 18 218 
rect 17 218 18 219 
rect 17 285 18 286 
rect 17 286 18 287 
rect 17 287 18 288 
rect 17 288 18 289 
rect 18 159 19 160 
rect 18 160 19 161 
rect 18 166 19 167 
rect 18 167 19 168 
rect 18 168 19 169 
rect 18 169 19 170 
rect 19 159 20 160 
rect 19 162 20 163 
rect 19 163 20 164 
rect 19 164 20 165 
rect 19 165 20 166 
rect 19 169 20 170 
rect 19 170 20 171 
rect 19 172 20 173 
rect 20 159 21 160 
rect 20 168 21 169 
rect 20 170 21 171 
rect 20 172 21 173 
rect 20 219 21 220 
rect 21 159 22 160 
rect 21 168 22 169 
rect 21 170 22 171 
rect 21 172 22 173 
rect 21 219 22 220 
rect 22 98 23 99 
rect 22 99 23 100 
rect 22 100 23 101 
rect 22 101 23 102 
rect 22 102 23 103 
rect 22 103 23 104 
rect 22 104 23 105 
rect 22 105 23 106 
rect 22 106 23 107 
rect 22 107 23 108 
rect 22 108 23 109 
rect 22 109 23 110 
rect 22 110 23 111 
rect 22 111 23 112 
rect 22 112 23 113 
rect 22 113 23 114 
rect 22 114 23 115 
rect 22 115 23 116 
rect 22 116 23 117 
rect 22 117 23 118 
rect 22 118 23 119 
rect 22 119 23 120 
rect 22 120 23 121 
rect 22 121 23 122 
rect 22 122 23 123 
rect 22 123 23 124 
rect 22 124 23 125 
rect 22 125 23 126 
rect 22 126 23 127 
rect 22 127 23 128 
rect 22 128 23 129 
rect 22 129 23 130 
rect 22 130 23 131 
rect 22 131 23 132 
rect 22 132 23 133 
rect 22 133 23 134 
rect 22 134 23 135 
rect 22 135 23 136 
rect 22 136 23 137 
rect 22 137 23 138 
rect 22 138 23 139 
rect 22 139 23 140 
rect 22 140 23 141 
rect 22 141 23 142 
rect 22 142 23 143 
rect 22 143 23 144 
rect 22 144 23 145 
rect 22 145 23 146 
rect 22 146 23 147 
rect 22 147 23 148 
rect 22 148 23 149 
rect 22 149 23 150 
rect 22 150 23 151 
rect 22 151 23 152 
rect 22 152 23 153 
rect 22 153 23 154 
rect 22 154 23 155 
rect 22 155 23 156 
rect 22 156 23 157 
rect 22 157 23 158 
rect 22 158 23 159 
rect 22 159 23 160 
rect 22 161 23 162 
rect 22 162 23 163 
rect 22 163 23 164 
rect 22 164 23 165 
rect 22 168 23 169 
rect 22 170 23 171 
rect 22 172 23 173 
rect 22 219 23 220 
rect 23 168 24 169 
rect 23 170 24 171 
rect 23 172 24 173 
rect 23 219 24 220 
rect 24 137 25 138 
rect 24 138 25 139 
rect 24 170 25 171 
rect 24 172 25 173 
rect 24 173 25 174 
rect 24 174 25 175 
rect 24 175 25 176 
rect 24 176 25 177 
rect 24 200 25 201 
rect 24 201 25 202 
rect 24 202 25 203 
rect 24 203 25 204 
rect 24 204 25 205 
rect 24 205 25 206 
rect 25 133 26 134 
rect 25 134 26 135 
rect 25 135 26 136 
rect 25 136 26 137 
rect 25 137 26 138 
rect 25 176 26 177 
rect 25 177 26 178 
rect 26 98 27 99 
rect 26 99 27 100 
rect 26 100 27 101 
rect 26 101 27 102 
rect 26 177 27 178 
rect 27 177 28 178 
rect 28 177 29 178 
rect 29 177 30 178 
rect 30 123 31 124 
rect 30 177 31 178 
rect 31 123 32 124 
rect 31 162 32 163 
rect 31 163 32 164 
rect 31 164 32 165 
rect 31 165 32 166 
rect 31 166 32 167 
rect 31 167 32 168 
rect 31 168 32 169 
rect 31 177 32 178 
rect 32 123 33 124 
rect 32 132 33 133 
rect 32 133 33 134 
rect 32 134 33 135 
rect 32 135 33 136 
rect 32 136 33 137 
rect 32 137 33 138 
rect 32 144 33 145 
rect 32 145 33 146 
rect 32 146 33 147 
rect 32 147 33 148 
rect 32 148 33 149 
rect 32 149 33 150 
rect 32 150 33 151 
rect 32 151 33 152 
rect 32 152 33 153 
rect 32 153 33 154 
rect 32 168 33 169 
rect 32 169 33 170 
rect 32 177 33 178 
rect 33 123 34 124 
rect 33 132 34 133 
rect 33 137 34 138 
rect 33 138 34 139 
rect 33 139 34 140 
rect 33 140 34 141 
rect 33 141 34 142 
rect 33 142 34 143 
rect 33 143 34 144 
rect 33 144 34 145 
rect 33 153 34 154 
rect 33 154 34 155 
rect 33 155 34 156 
rect 33 156 34 157 
rect 33 157 34 158 
rect 33 158 34 159 
rect 33 159 34 160 
rect 33 160 34 161 
rect 33 161 34 162 
rect 33 162 34 163 
rect 33 163 34 164 
rect 33 164 34 165 
rect 33 165 34 166 
rect 33 166 34 167 
rect 33 167 34 168 
rect 33 169 34 170 
rect 33 177 34 178 
rect 34 123 35 124 
rect 34 132 35 133 
rect 34 167 35 168 
rect 34 169 35 170 
rect 34 177 35 178 
rect 35 67 36 68 
rect 35 99 36 100 
rect 35 123 36 124 
rect 35 130 36 131 
rect 35 132 36 133 
rect 35 134 36 135 
rect 35 136 36 137 
rect 35 145 36 146 
rect 35 167 36 168 
rect 35 169 36 170 
rect 35 170 36 171 
rect 35 177 36 178 
rect 36 67 37 68 
rect 36 99 37 100 
rect 36 123 37 124 
rect 36 130 37 131 
rect 36 132 37 133 
rect 36 134 37 135 
rect 36 136 37 137 
rect 36 145 37 146 
rect 36 157 37 158 
rect 36 160 37 161 
rect 36 161 37 162 
rect 36 162 37 163 
rect 36 163 37 164 
rect 36 164 37 165 
rect 36 165 37 166 
rect 36 167 37 168 
rect 36 168 37 169 
rect 36 170 37 171 
rect 36 177 37 178 
rect 36 200 37 201 
rect 37 67 38 68 
rect 37 99 38 100 
rect 37 123 38 124 
rect 37 130 38 131 
rect 37 132 38 133 
rect 37 134 38 135 
rect 37 136 38 137 
rect 37 145 38 146 
rect 37 157 38 158 
rect 37 159 38 160 
rect 37 160 38 161 
rect 37 168 38 169 
rect 37 170 38 171 
rect 37 177 38 178 
rect 37 200 38 201 
rect 38 67 39 68 
rect 38 81 39 82 
rect 38 82 39 83 
rect 38 83 39 84 
rect 38 84 39 85 
rect 38 99 39 100 
rect 38 123 39 124 
rect 38 130 39 131 
rect 38 134 39 135 
rect 38 136 39 137 
rect 38 145 39 146 
rect 38 152 39 153 
rect 38 153 39 154 
rect 38 154 39 155 
rect 38 155 39 156 
rect 38 156 39 157 
rect 38 157 39 158 
rect 38 159 39 160 
rect 38 162 39 163 
rect 38 163 39 164 
rect 38 164 39 165 
rect 38 165 39 166 
rect 38 168 39 169 
rect 38 170 39 171 
rect 38 177 39 178 
rect 38 178 39 179 
rect 38 179 39 180 
rect 38 180 39 181 
rect 38 181 39 182 
rect 38 182 39 183 
rect 38 183 39 184 
rect 38 184 39 185 
rect 38 185 39 186 
rect 38 186 39 187 
rect 38 187 39 188 
rect 38 188 39 189 
rect 38 189 39 190 
rect 38 190 39 191 
rect 38 191 39 192 
rect 38 192 39 193 
rect 38 193 39 194 
rect 38 200 39 201 
rect 39 67 40 68 
rect 39 99 40 100 
rect 39 123 40 124 
rect 39 130 40 131 
rect 39 131 40 132 
rect 39 136 40 137 
rect 39 145 40 146 
rect 39 151 40 152 
rect 39 152 40 153 
rect 39 159 40 160 
rect 39 168 40 169 
rect 39 170 40 171 
rect 39 193 40 194 
rect 39 200 40 201 
rect 40 67 41 68 
rect 40 89 41 90 
rect 40 90 41 91 
rect 40 91 41 92 
rect 40 92 41 93 
rect 40 93 41 94 
rect 40 94 41 95 
rect 40 95 41 96 
rect 40 96 41 97 
rect 40 99 41 100 
rect 40 105 41 106 
rect 40 106 41 107 
rect 40 107 41 108 
rect 40 108 41 109 
rect 40 109 41 110 
rect 40 110 41 111 
rect 40 111 41 112 
rect 40 112 41 113 
rect 40 121 41 122 
rect 40 122 41 123 
rect 40 123 41 124 
rect 40 131 41 132 
rect 40 132 41 133 
rect 40 133 41 134 
rect 40 136 41 137 
rect 40 145 41 146 
rect 40 150 41 151 
rect 40 151 41 152 
rect 40 153 41 154 
rect 40 154 41 155 
rect 40 155 41 156 
rect 40 156 41 157 
rect 40 157 41 158 
rect 40 158 41 159 
rect 40 159 41 160 
rect 40 161 41 162 
rect 40 162 41 163 
rect 40 163 41 164 
rect 40 164 41 165 
rect 40 168 41 169 
rect 40 170 41 171 
rect 40 171 41 172 
rect 40 172 41 173 
rect 40 173 41 174 
rect 40 174 41 175 
rect 40 175 41 176 
rect 40 176 41 177 
rect 40 177 41 178 
rect 40 178 41 179 
rect 40 179 41 180 
rect 40 180 41 181 
rect 40 181 41 182 
rect 40 182 41 183 
rect 40 183 41 184 
rect 40 184 41 185 
rect 40 185 41 186 
rect 40 186 41 187 
rect 40 187 41 188 
rect 40 188 41 189 
rect 40 189 41 190 
rect 40 190 41 191 
rect 40 191 41 192 
rect 40 192 41 193 
rect 40 200 41 201 
rect 41 67 42 68 
rect 41 88 42 89 
rect 41 89 42 90 
rect 41 96 42 97 
rect 41 97 42 98 
rect 41 99 42 100 
rect 41 104 42 105 
rect 41 105 42 106 
rect 41 112 42 113 
rect 41 113 42 114 
rect 41 120 42 121 
rect 41 121 42 122 
rect 41 133 42 134 
rect 41 136 42 137 
rect 41 150 42 151 
rect 41 152 42 153 
rect 41 153 42 154 
rect 41 168 42 169 
rect 41 192 42 193 
rect 41 193 42 194 
rect 41 200 42 201 
rect 42 67 43 68 
rect 42 88 43 89 
rect 42 99 43 100 
rect 42 104 43 105 
rect 42 120 43 121 
rect 42 133 43 134 
rect 42 136 43 137 
rect 42 150 43 151 
rect 42 152 43 153 
rect 42 168 43 169 
rect 42 193 43 194 
rect 42 200 43 201 
rect 43 67 44 68 
rect 43 88 44 89 
rect 43 99 44 100 
rect 43 120 44 121 
rect 43 133 44 134 
rect 43 136 44 137 
rect 43 150 44 151 
rect 43 152 44 153 
rect 43 168 44 169 
rect 43 193 44 194 
rect 43 200 44 201 
rect 44 67 45 68 
rect 44 88 45 89 
rect 44 99 45 100 
rect 44 120 45 121 
rect 44 133 45 134 
rect 44 136 45 137 
rect 44 150 45 151 
rect 44 152 45 153 
rect 44 168 45 169 
rect 44 193 45 194 
rect 44 200 45 201 
rect 45 53 46 54 
rect 45 54 46 55 
rect 45 55 46 56 
rect 45 56 46 57 
rect 45 67 46 68 
rect 45 88 46 89 
rect 45 99 46 100 
rect 45 120 46 121 
rect 45 133 46 134 
rect 45 136 46 137 
rect 45 150 46 151 
rect 45 152 46 153 
rect 45 168 46 169 
rect 45 193 46 194 
rect 45 194 46 195 
rect 45 200 46 201 
rect 46 52 47 53 
rect 46 53 47 54 
rect 46 67 47 68 
rect 46 88 47 89 
rect 46 99 47 100 
rect 46 120 47 121 
rect 46 133 47 134 
rect 46 136 47 137 
rect 46 150 47 151 
rect 46 152 47 153 
rect 46 168 47 169 
rect 46 194 47 195 
rect 46 195 47 196 
rect 46 200 47 201 
rect 47 52 48 53 
rect 47 67 48 68 
rect 47 88 48 89 
rect 47 99 48 100 
rect 47 116 48 117 
rect 47 120 48 121 
rect 47 133 48 134 
rect 47 136 48 137 
rect 47 145 48 146 
rect 47 150 48 151 
rect 47 152 48 153 
rect 47 168 48 169 
rect 47 195 48 196 
rect 47 200 48 201 
rect 47 212 48 213 
rect 47 215 48 216 
rect 47 228 48 229 
rect 48 49 49 50 
rect 48 52 49 53 
rect 48 54 49 55 
rect 48 67 49 68 
rect 48 88 49 89 
rect 48 99 49 100 
rect 48 116 49 117 
rect 48 120 49 121 
rect 48 133 49 134 
rect 48 136 49 137 
rect 48 145 49 146 
rect 48 150 49 151 
rect 48 152 49 153 
rect 48 168 49 169 
rect 48 193 49 194 
rect 48 195 49 196 
rect 48 197 49 198 
rect 48 200 49 201 
rect 48 212 49 213 
rect 48 215 49 216 
rect 48 228 49 229 
rect 49 49 50 50 
rect 49 52 50 53 
rect 49 54 50 55 
rect 49 67 50 68 
rect 49 88 50 89 
rect 49 97 50 98 
rect 49 99 50 100 
rect 49 101 50 102 
rect 49 102 50 103 
rect 49 103 50 104 
rect 49 104 50 105 
rect 49 105 50 106 
rect 49 106 50 107 
rect 49 116 50 117 
rect 49 120 50 121 
rect 49 133 50 134 
rect 49 136 50 137 
rect 49 145 50 146 
rect 49 150 50 151 
rect 49 152 50 153 
rect 49 161 50 162 
rect 49 162 50 163 
rect 49 163 50 164 
rect 49 164 50 165 
rect 49 168 50 169 
rect 49 193 50 194 
rect 49 195 50 196 
rect 49 197 50 198 
rect 49 200 50 201 
rect 49 212 50 213 
rect 49 215 50 216 
rect 49 228 50 229 
rect 49 230 50 231 
rect 49 231 50 232 
rect 49 232 50 233 
rect 49 233 50 234 
rect 49 234 50 235 
rect 49 235 50 236 
rect 49 236 50 237 
rect 49 237 50 238 
rect 49 238 50 239 
rect 49 239 50 240 
rect 49 240 50 241 
rect 49 241 50 242 
rect 49 242 50 243 
rect 49 243 50 244 
rect 49 244 50 245 
rect 49 245 50 246 
rect 50 49 51 50 
rect 50 52 51 53 
rect 50 54 51 55 
rect 50 67 51 68 
rect 50 80 51 81 
rect 50 81 51 82 
rect 50 82 51 83 
rect 50 83 51 84 
rect 50 88 51 89 
rect 50 97 51 98 
rect 50 99 51 100 
rect 50 106 51 107 
rect 50 107 51 108 
rect 50 116 51 117 
rect 50 120 51 121 
rect 50 133 51 134 
rect 50 136 51 137 
rect 50 145 51 146 
rect 50 150 51 151 
rect 50 152 51 153 
rect 50 168 51 169 
rect 50 193 51 194 
rect 50 195 51 196 
rect 50 197 51 198 
rect 50 200 51 201 
rect 50 212 51 213 
rect 50 215 51 216 
rect 50 228 51 229 
rect 50 229 51 230 
rect 51 49 52 50 
rect 51 52 52 53 
rect 51 54 52 55 
rect 51 67 52 68 
rect 51 88 52 89 
rect 51 97 52 98 
rect 51 99 52 100 
rect 51 101 52 102 
rect 51 102 52 103 
rect 51 103 52 104 
rect 51 104 52 105 
rect 51 107 52 108 
rect 51 116 52 117 
rect 51 120 52 121 
rect 51 133 52 134 
rect 51 136 52 137 
rect 51 145 52 146 
rect 51 150 52 151 
rect 51 152 52 153 
rect 51 161 52 162 
rect 51 162 52 163 
rect 51 163 52 164 
rect 51 164 52 165 
rect 51 168 52 169 
rect 51 193 52 194 
rect 51 195 52 196 
rect 51 197 52 198 
rect 51 200 52 201 
rect 51 212 52 213 
rect 51 229 52 230 
rect 51 230 52 231 
rect 51 231 52 232 
rect 51 232 52 233 
rect 51 233 52 234 
rect 51 234 52 235 
rect 52 51 53 52 
rect 52 52 53 53 
rect 52 54 53 55 
rect 52 67 53 68 
rect 52 80 53 81 
rect 52 81 53 82 
rect 52 82 53 83 
rect 52 83 53 84 
rect 52 84 53 85 
rect 52 85 53 86 
rect 52 86 53 87 
rect 52 87 53 88 
rect 52 88 53 89 
rect 52 97 53 98 
rect 52 99 53 100 
rect 52 100 53 101 
rect 52 107 53 108 
rect 52 116 53 117 
rect 52 120 53 121 
rect 52 133 53 134 
rect 52 136 53 137 
rect 52 145 53 146 
rect 52 150 53 151 
rect 52 152 53 153 
rect 52 168 53 169 
rect 52 193 53 194 
rect 52 195 53 196 
rect 52 197 53 198 
rect 52 200 53 201 
rect 52 212 53 213 
rect 53 51 54 52 
rect 53 54 54 55 
rect 53 67 54 68 
rect 53 97 54 98 
rect 53 100 54 101 
rect 53 107 54 108 
rect 53 116 54 117 
rect 53 120 54 121 
rect 53 133 54 134 
rect 53 136 54 137 
rect 53 145 54 146 
rect 53 150 54 151 
rect 53 168 54 169 
rect 53 193 54 194 
rect 53 195 54 196 
rect 53 197 54 198 
rect 53 200 54 201 
rect 53 212 54 213 
rect 54 51 55 52 
rect 54 54 55 55 
rect 54 67 55 68 
rect 54 97 55 98 
rect 54 100 55 101 
rect 54 107 55 108 
rect 54 116 55 117 
rect 54 120 55 121 
rect 54 129 55 130 
rect 54 133 55 134 
rect 54 136 55 137 
rect 54 145 55 146 
rect 54 150 55 151 
rect 54 160 55 161 
rect 54 161 55 162 
rect 54 162 55 163 
rect 54 163 55 164 
rect 54 164 55 165 
rect 54 168 55 169 
rect 54 193 55 194 
rect 54 197 55 198 
rect 54 200 55 201 
rect 54 212 55 213 
rect 54 231 55 232 
rect 54 232 55 233 
rect 54 233 55 234 
rect 54 234 55 235 
rect 54 235 55 236 
rect 54 236 55 237 
rect 54 237 55 238 
rect 54 238 55 239 
rect 54 239 55 240 
rect 54 240 55 241 
rect 54 241 55 242 
rect 54 242 55 243 
rect 54 243 55 244 
rect 54 244 55 245 
rect 54 245 55 246 
rect 54 246 55 247 
rect 55 51 56 52 
rect 55 54 56 55 
rect 55 67 56 68 
rect 55 79 56 80 
rect 55 80 56 81 
rect 55 81 56 82 
rect 55 82 56 83 
rect 55 83 56 84 
rect 55 84 56 85 
rect 55 85 56 86 
rect 55 86 56 87 
rect 55 87 56 88 
rect 55 88 56 89 
rect 55 89 56 90 
rect 55 90 56 91 
rect 55 91 56 92 
rect 55 92 56 93 
rect 55 93 56 94 
rect 55 94 56 95 
rect 55 95 56 96 
rect 55 96 56 97 
rect 55 97 56 98 
rect 55 100 56 101 
rect 55 107 56 108 
rect 55 116 56 117 
rect 55 120 56 121 
rect 55 129 56 130 
rect 55 133 56 134 
rect 55 136 56 137 
rect 55 145 56 146 
rect 55 150 56 151 
rect 55 159 56 160 
rect 55 160 56 161 
rect 55 168 56 169 
rect 55 193 56 194 
rect 55 197 56 198 
rect 55 200 56 201 
rect 55 212 56 213 
rect 56 51 57 52 
rect 56 54 57 55 
rect 56 67 57 68 
rect 56 73 57 74 
rect 56 74 57 75 
rect 56 75 57 76 
rect 56 76 57 77 
rect 56 77 57 78 
rect 56 78 57 79 
rect 56 79 57 80 
rect 56 100 57 101 
rect 56 107 57 108 
rect 56 108 57 109 
rect 56 109 57 110 
rect 56 110 57 111 
rect 56 111 57 112 
rect 56 112 57 113 
rect 56 116 57 117 
rect 56 120 57 121 
rect 56 129 57 130 
rect 56 133 57 134 
rect 56 136 57 137 
rect 56 145 57 146 
rect 56 150 57 151 
rect 56 153 57 154 
rect 56 154 57 155 
rect 56 155 57 156 
rect 56 156 57 157 
rect 56 157 57 158 
rect 56 158 57 159 
rect 56 159 57 160 
rect 56 161 57 162 
rect 56 162 57 163 
rect 56 163 57 164 
rect 56 164 57 165 
rect 56 168 57 169 
rect 56 193 57 194 
rect 56 197 57 198 
rect 56 200 57 201 
rect 56 212 57 213 
rect 56 233 57 234 
rect 56 234 57 235 
rect 56 271 57 272 
rect 56 272 57 273 
rect 56 273 57 274 
rect 56 274 57 275 
rect 56 303 57 304 
rect 56 304 57 305 
rect 56 305 57 306 
rect 56 306 57 307 
rect 56 307 57 308 
rect 56 308 57 309 
rect 56 309 57 310 
rect 57 51 58 52 
rect 57 54 58 55 
rect 57 56 58 57 
rect 57 67 58 68 
rect 57 72 58 73 
rect 57 73 58 74 
rect 57 81 58 82 
rect 57 100 58 101 
rect 57 103 58 104 
rect 57 112 58 113 
rect 57 113 58 114 
rect 57 116 58 117 
rect 57 120 58 121 
rect 57 129 58 130 
rect 57 133 58 134 
rect 57 136 58 137 
rect 57 145 58 146 
rect 57 150 58 151 
rect 57 152 58 153 
rect 57 153 58 154 
rect 57 168 58 169 
rect 57 193 58 194 
rect 57 197 58 198 
rect 57 200 58 201 
rect 57 212 58 213 
rect 57 232 58 233 
rect 57 233 58 234 
rect 57 261 58 262 
rect 58 51 59 52 
rect 58 54 59 55 
rect 58 56 59 57 
rect 58 67 59 68 
rect 58 72 59 73 
rect 58 81 59 82 
rect 58 82 59 83 
rect 58 83 59 84 
rect 58 84 59 85 
rect 58 85 59 86 
rect 58 86 59 87 
rect 58 100 59 101 
rect 58 103 59 104 
rect 58 113 59 114 
rect 58 116 59 117 
rect 58 120 59 121 
rect 58 129 59 130 
rect 58 133 59 134 
rect 58 136 59 137 
rect 58 145 59 146 
rect 58 148 59 149 
rect 58 149 59 150 
rect 58 150 59 151 
rect 58 152 59 153 
rect 58 168 59 169 
rect 58 193 59 194 
rect 58 197 59 198 
rect 58 200 59 201 
rect 58 212 59 213 
rect 58 232 59 233 
rect 58 261 59 262 
rect 59 51 60 52 
rect 59 54 60 55 
rect 59 56 60 57 
rect 59 67 60 68 
rect 59 72 60 73 
rect 59 86 60 87 
rect 59 100 60 101 
rect 59 103 60 104 
rect 59 113 60 114 
rect 59 116 60 117 
rect 59 120 60 121 
rect 59 129 60 130 
rect 59 133 60 134 
rect 59 136 60 137 
rect 59 145 60 146 
rect 59 148 60 149 
rect 59 152 60 153 
rect 59 168 60 169 
rect 59 193 60 194 
rect 59 197 60 198 
rect 59 200 60 201 
rect 59 212 60 213 
rect 59 232 60 233 
rect 59 261 60 262 
rect 60 51 61 52 
rect 60 54 61 55 
rect 60 56 61 57 
rect 60 67 61 68 
rect 60 72 61 73 
rect 60 86 61 87 
rect 60 100 61 101 
rect 60 103 61 104 
rect 60 113 61 114 
rect 60 116 61 117 
rect 60 120 61 121 
rect 60 129 61 130 
rect 60 133 61 134 
rect 60 136 61 137 
rect 60 145 61 146 
rect 60 148 61 149 
rect 60 152 61 153 
rect 60 168 61 169 
rect 60 193 61 194 
rect 60 197 61 198 
rect 60 200 61 201 
rect 60 212 61 213 
rect 60 232 61 233 
rect 60 261 61 262 
rect 61 54 62 55 
rect 61 56 62 57 
rect 61 67 62 68 
rect 61 72 62 73 
rect 61 86 62 87 
rect 61 100 62 101 
rect 61 103 62 104 
rect 61 113 62 114 
rect 61 116 62 117 
rect 61 119 62 120 
rect 61 120 62 121 
rect 61 129 62 130 
rect 61 133 62 134 
rect 61 136 62 137 
rect 61 145 62 146 
rect 61 148 62 149 
rect 61 152 62 153 
rect 61 162 62 163 
rect 61 163 62 164 
rect 61 164 62 165 
rect 61 165 62 166 
rect 61 166 62 167 
rect 61 168 62 169 
rect 61 193 62 194 
rect 61 197 62 198 
rect 61 200 62 201 
rect 61 212 62 213 
rect 61 231 62 232 
rect 61 232 62 233 
rect 61 261 62 262 
rect 62 54 63 55 
rect 62 56 63 57 
rect 62 67 63 68 
rect 62 72 63 73 
rect 62 86 63 87 
rect 62 100 63 101 
rect 62 103 63 104 
rect 62 113 63 114 
rect 62 116 63 117 
rect 62 119 63 120 
rect 62 129 63 130 
rect 62 133 63 134 
rect 62 136 63 137 
rect 62 145 63 146 
rect 62 148 63 149 
rect 62 152 63 153 
rect 62 161 63 162 
rect 62 162 63 163 
rect 62 166 63 167 
rect 62 168 63 169 
rect 62 193 63 194 
rect 62 197 63 198 
rect 62 200 63 201 
rect 62 212 63 213 
rect 62 231 63 232 
rect 62 261 63 262 
rect 63 54 64 55 
rect 63 56 64 57 
rect 63 67 64 68 
rect 63 72 64 73 
rect 63 86 64 87 
rect 63 100 64 101 
rect 63 103 64 104 
rect 63 113 64 114 
rect 63 116 64 117 
rect 63 119 64 120 
rect 63 129 64 130 
rect 63 133 64 134 
rect 63 136 64 137 
rect 63 145 64 146 
rect 63 148 64 149 
rect 63 152 64 153 
rect 63 161 64 162 
rect 63 166 64 167 
rect 63 168 64 169 
rect 63 193 64 194 
rect 63 197 64 198 
rect 63 200 64 201 
rect 63 212 64 213 
rect 63 225 64 226 
rect 63 231 64 232 
rect 63 261 64 262 
rect 64 54 65 55 
rect 64 56 65 57 
rect 64 67 65 68 
rect 64 71 65 72 
rect 64 72 65 73 
rect 64 86 65 87 
rect 64 98 65 99 
rect 64 100 65 101 
rect 64 103 65 104 
rect 64 113 65 114 
rect 64 116 65 117 
rect 64 119 65 120 
rect 64 129 65 130 
rect 64 133 65 134 
rect 64 136 65 137 
rect 64 145 65 146 
rect 64 148 65 149 
rect 64 152 65 153 
rect 64 161 65 162 
rect 64 163 65 164 
rect 64 166 65 167 
rect 64 168 65 169 
rect 64 193 65 194 
rect 64 197 65 198 
rect 64 200 65 201 
rect 64 212 65 213 
rect 64 225 65 226 
rect 64 231 65 232 
rect 64 261 65 262 
rect 65 54 66 55 
rect 65 56 66 57 
rect 65 67 66 68 
rect 65 71 66 72 
rect 65 74 66 75 
rect 65 75 66 76 
rect 65 76 66 77 
rect 65 77 66 78 
rect 65 78 66 79 
rect 65 79 66 80 
rect 65 80 66 81 
rect 65 81 66 82 
rect 65 82 66 83 
rect 65 83 66 84 
rect 65 84 66 85 
rect 65 86 66 87 
rect 65 98 66 99 
rect 65 100 66 101 
rect 65 103 66 104 
rect 65 113 66 114 
rect 65 116 66 117 
rect 65 119 66 120 
rect 65 129 66 130 
rect 65 133 66 134 
rect 65 136 66 137 
rect 65 145 66 146 
rect 65 148 66 149 
rect 65 152 66 153 
rect 65 161 66 162 
rect 65 163 66 164 
rect 65 166 66 167 
rect 65 168 66 169 
rect 65 193 66 194 
rect 65 197 66 198 
rect 65 200 66 201 
rect 65 212 66 213 
rect 65 225 66 226 
rect 65 231 66 232 
rect 65 261 66 262 
rect 66 54 67 55 
rect 66 56 67 57 
rect 66 67 67 68 
rect 66 71 67 72 
rect 66 86 67 87 
rect 66 98 67 99 
rect 66 100 67 101 
rect 66 103 67 104 
rect 66 113 67 114 
rect 66 116 67 117 
rect 66 119 67 120 
rect 66 129 67 130 
rect 66 133 67 134 
rect 66 136 67 137 
rect 66 145 67 146 
rect 66 148 67 149 
rect 66 152 67 153 
rect 66 161 67 162 
rect 66 163 67 164 
rect 66 166 67 167 
rect 66 168 67 169 
rect 66 193 67 194 
rect 66 197 67 198 
rect 66 200 67 201 
rect 66 212 67 213 
rect 66 225 67 226 
rect 66 231 67 232 
rect 66 240 67 241 
rect 66 241 67 242 
rect 66 242 67 243 
rect 66 243 67 244 
rect 66 244 67 245 
rect 66 245 67 246 
rect 66 261 67 262 
rect 67 54 68 55 
rect 67 56 68 57 
rect 67 67 68 68 
rect 67 70 68 71 
rect 67 71 68 72 
rect 67 86 68 87 
rect 67 98 68 99 
rect 67 100 68 101 
rect 67 103 68 104 
rect 67 113 68 114 
rect 67 116 68 117 
rect 67 119 68 120 
rect 67 129 68 130 
rect 67 133 68 134 
rect 67 136 68 137 
rect 67 145 68 146 
rect 67 148 68 149 
rect 67 152 68 153 
rect 67 161 68 162 
rect 67 163 68 164 
rect 67 166 68 167 
rect 67 168 68 169 
rect 67 193 68 194 
rect 67 197 68 198 
rect 67 200 68 201 
rect 67 212 68 213 
rect 67 225 68 226 
rect 67 231 68 232 
rect 67 261 68 262 
rect 68 54 69 55 
rect 68 56 69 57 
rect 68 67 69 68 
rect 68 70 69 71 
rect 68 72 69 73 
rect 68 73 69 74 
rect 68 74 69 75 
rect 68 86 69 87 
rect 68 88 69 89 
rect 68 98 69 99 
rect 68 100 69 101 
rect 68 103 69 104 
rect 68 113 69 114 
rect 68 116 69 117 
rect 68 119 69 120 
rect 68 129 69 130 
rect 68 133 69 134 
rect 68 136 69 137 
rect 68 145 69 146 
rect 68 148 69 149 
rect 68 152 69 153 
rect 68 161 69 162 
rect 68 163 69 164 
rect 68 166 69 167 
rect 68 193 69 194 
rect 68 200 69 201 
rect 68 210 69 211 
rect 68 215 69 216 
rect 68 216 69 217 
rect 68 217 69 218 
rect 68 225 69 226 
rect 68 231 69 232 
rect 68 239 69 240 
rect 68 240 69 241 
rect 68 241 69 242 
rect 68 242 69 243 
rect 68 243 69 244 
rect 68 244 69 245 
rect 68 245 69 246 
rect 68 246 69 247 
rect 68 247 69 248 
rect 68 248 69 249 
rect 68 249 69 250 
rect 68 250 69 251 
rect 68 251 69 252 
rect 68 252 69 253 
rect 68 253 69 254 
rect 68 254 69 255 
rect 68 255 69 256 
rect 68 256 69 257 
rect 68 257 69 258 
rect 68 258 69 259 
rect 68 261 69 262 
rect 69 54 70 55 
rect 69 56 70 57 
rect 69 65 70 66 
rect 69 67 70 68 
rect 69 70 70 71 
rect 69 72 70 73 
rect 69 86 70 87 
rect 69 88 70 89 
rect 69 98 70 99 
rect 69 100 70 101 
rect 69 103 70 104 
rect 69 113 70 114 
rect 69 116 70 117 
rect 69 119 70 120 
rect 69 129 70 130 
rect 69 131 70 132 
rect 69 133 70 134 
rect 69 136 70 137 
rect 69 145 70 146 
rect 69 148 70 149 
rect 69 152 70 153 
rect 69 161 70 162 
rect 69 163 70 164 
rect 69 166 70 167 
rect 69 167 70 168 
rect 69 193 70 194 
rect 69 200 70 201 
rect 69 210 70 211 
rect 69 214 70 215 
rect 69 215 70 216 
rect 69 217 70 218 
rect 69 218 70 219 
rect 69 225 70 226 
rect 69 231 70 232 
rect 69 239 70 240 
rect 69 261 70 262 
rect 70 54 71 55 
rect 70 56 71 57 
rect 70 65 71 66 
rect 70 67 71 68 
rect 70 70 71 71 
rect 70 72 71 73 
rect 70 86 71 87 
rect 70 88 71 89 
rect 70 98 71 99 
rect 70 100 71 101 
rect 70 103 71 104 
rect 70 113 71 114 
rect 70 116 71 117 
rect 70 119 71 120 
rect 70 129 71 130 
rect 70 131 71 132 
rect 70 133 71 134 
rect 70 136 71 137 
rect 70 145 71 146 
rect 70 148 71 149 
rect 70 152 71 153 
rect 70 161 71 162 
rect 70 163 71 164 
rect 70 167 71 168 
rect 70 193 71 194 
rect 70 200 71 201 
rect 70 210 71 211 
rect 70 214 71 215 
rect 70 225 71 226 
rect 70 231 71 232 
rect 70 239 71 240 
rect 70 257 71 258 
rect 70 261 71 262 
rect 70 276 71 277 
rect 71 54 72 55 
rect 71 56 72 57 
rect 71 65 72 66 
rect 71 67 72 68 
rect 71 70 72 71 
rect 71 72 72 73 
rect 71 86 72 87 
rect 71 88 72 89 
rect 71 98 72 99 
rect 71 100 72 101 
rect 71 103 72 104 
rect 71 113 72 114 
rect 71 116 72 117 
rect 71 119 72 120 
rect 71 129 72 130 
rect 71 131 72 132 
rect 71 133 72 134 
rect 71 136 72 137 
rect 71 145 72 146 
rect 71 148 72 149 
rect 71 152 72 153 
rect 71 161 72 162 
rect 71 163 72 164 
rect 71 165 72 166 
rect 71 167 72 168 
rect 71 193 72 194 
rect 71 200 72 201 
rect 71 210 72 211 
rect 71 214 72 215 
rect 71 216 72 217 
rect 71 225 72 226 
rect 71 227 72 228 
rect 71 231 72 232 
rect 71 239 72 240 
rect 71 241 72 242 
rect 71 243 72 244 
rect 71 245 72 246 
rect 71 257 72 258 
rect 71 261 72 262 
rect 71 276 72 277 
rect 72 19 73 20 
rect 72 20 73 21 
rect 72 21 73 22 
rect 72 22 73 23 
rect 72 23 73 24 
rect 72 24 73 25 
rect 72 25 73 26 
rect 72 26 73 27 
rect 72 38 73 39 
rect 72 54 73 55 
rect 72 56 73 57 
rect 72 65 73 66 
rect 72 67 73 68 
rect 72 70 73 71 
rect 72 72 73 73 
rect 72 86 73 87 
rect 72 88 73 89 
rect 72 98 73 99 
rect 72 100 73 101 
rect 72 103 73 104 
rect 72 113 73 114 
rect 72 116 73 117 
rect 72 119 73 120 
rect 72 129 73 130 
rect 72 131 73 132 
rect 72 133 73 134 
rect 72 136 73 137 
rect 72 145 73 146 
rect 72 148 73 149 
rect 72 152 73 153 
rect 72 161 73 162 
rect 72 163 73 164 
rect 72 165 73 166 
rect 72 167 73 168 
rect 72 193 73 194 
rect 72 200 73 201 
rect 72 210 73 211 
rect 72 214 73 215 
rect 72 216 73 217 
rect 72 225 73 226 
rect 72 227 73 228 
rect 72 230 73 231 
rect 72 231 73 232 
rect 72 233 73 234 
rect 72 234 73 235 
rect 72 235 73 236 
rect 72 236 73 237 
rect 72 237 73 238 
rect 72 238 73 239 
rect 72 239 73 240 
rect 72 241 73 242 
rect 72 243 73 244 
rect 72 245 73 246 
rect 72 257 73 258 
rect 72 261 73 262 
rect 72 276 73 277 
rect 73 19 74 20 
rect 73 38 74 39 
rect 73 54 74 55 
rect 73 56 74 57 
rect 73 65 74 66 
rect 73 67 74 68 
rect 73 70 74 71 
rect 73 72 74 73 
rect 73 86 74 87 
rect 73 88 74 89 
rect 73 98 74 99 
rect 73 100 74 101 
rect 73 103 74 104 
rect 73 113 74 114 
rect 73 116 74 117 
rect 73 119 74 120 
rect 73 129 74 130 
rect 73 131 74 132 
rect 73 133 74 134 
rect 73 136 74 137 
rect 73 145 74 146 
rect 73 148 74 149 
rect 73 152 74 153 
rect 73 161 74 162 
rect 73 163 74 164 
rect 73 165 74 166 
rect 73 167 74 168 
rect 73 193 74 194 
rect 73 200 74 201 
rect 73 210 74 211 
rect 73 214 74 215 
rect 73 216 74 217 
rect 73 225 74 226 
rect 73 227 74 228 
rect 73 230 74 231 
rect 73 232 74 233 
rect 73 233 74 234 
rect 73 241 74 242 
rect 73 243 74 244 
rect 73 245 74 246 
rect 73 257 74 258 
rect 73 261 74 262 
rect 73 276 74 277 
rect 74 19 75 20 
rect 74 38 75 39 
rect 74 54 75 55 
rect 74 56 75 57 
rect 74 65 75 66 
rect 74 67 75 68 
rect 74 70 75 71 
rect 74 72 75 73 
rect 74 86 75 87 
rect 74 88 75 89 
rect 74 98 75 99 
rect 74 100 75 101 
rect 74 103 75 104 
rect 74 113 75 114 
rect 74 116 75 117 
rect 74 119 75 120 
rect 74 131 75 132 
rect 74 133 75 134 
rect 74 136 75 137 
rect 74 145 75 146 
rect 74 152 75 153 
rect 74 161 75 162 
rect 74 163 75 164 
rect 74 165 75 166 
rect 74 167 75 168 
rect 74 193 75 194 
rect 74 200 75 201 
rect 74 210 75 211 
rect 74 214 75 215 
rect 74 216 75 217 
rect 74 225 75 226 
rect 74 227 75 228 
rect 74 230 75 231 
rect 74 232 75 233 
rect 74 241 75 242 
rect 74 243 75 244 
rect 74 245 75 246 
rect 74 261 75 262 
rect 74 276 75 277 
rect 75 19 76 20 
rect 75 38 76 39 
rect 75 54 76 55 
rect 75 67 76 68 
rect 75 86 76 87 
rect 75 88 76 89 
rect 75 98 76 99 
rect 75 100 76 101 
rect 75 113 76 114 
rect 75 116 76 117 
rect 75 119 76 120 
rect 75 145 76 146 
rect 75 161 76 162 
rect 75 163 76 164 
rect 75 167 76 168 
rect 75 193 76 194 
rect 75 200 76 201 
rect 75 214 76 215 
rect 75 216 76 217 
rect 75 225 76 226 
rect 75 227 76 228 
rect 75 230 76 231 
rect 75 243 76 244 
rect 75 261 76 262 
rect 75 276 76 277 
rect 76 19 77 20 
rect 76 38 77 39 
rect 76 54 77 55 
rect 76 67 77 68 
rect 76 86 77 87 
rect 76 88 77 89 
rect 76 98 77 99 
rect 76 100 77 101 
rect 76 113 77 114 
rect 76 116 77 117 
rect 76 119 77 120 
rect 76 145 77 146 
rect 76 161 77 162 
rect 76 163 77 164 
rect 76 167 77 168 
rect 76 193 77 194 
rect 76 200 77 201 
rect 76 214 77 215 
rect 76 216 77 217 
rect 76 227 77 228 
rect 76 230 77 231 
rect 76 243 77 244 
rect 76 261 77 262 
rect 76 276 77 277 
rect 77 19 78 20 
rect 77 38 78 39 
rect 77 54 78 55 
rect 77 67 78 68 
rect 77 86 78 87 
rect 77 88 78 89 
rect 77 98 78 99 
rect 77 113 78 114 
rect 77 116 78 117 
rect 77 119 78 120 
rect 77 145 78 146 
rect 77 161 78 162 
rect 77 163 78 164 
rect 77 167 78 168 
rect 77 193 78 194 
rect 77 200 78 201 
rect 77 214 78 215 
rect 77 216 78 217 
rect 77 227 78 228 
rect 77 230 78 231 
rect 77 243 78 244 
rect 77 261 78 262 
rect 77 276 78 277 
rect 78 19 79 20 
rect 78 38 79 39 
rect 78 54 79 55 
rect 78 67 79 68 
rect 78 86 79 87 
rect 78 88 79 89 
rect 78 98 79 99 
rect 78 113 79 114 
rect 78 116 79 117 
rect 78 119 79 120 
rect 78 145 79 146 
rect 78 161 79 162 
rect 78 163 79 164 
rect 78 167 79 168 
rect 78 193 79 194 
rect 78 200 79 201 
rect 78 214 79 215 
rect 78 216 79 217 
rect 78 227 79 228 
rect 78 230 79 231 
rect 78 243 79 244 
rect 78 261 79 262 
rect 78 276 79 277 
rect 79 19 80 20 
rect 79 38 80 39 
rect 79 54 80 55 
rect 79 67 80 68 
rect 79 86 80 87 
rect 79 88 80 89 
rect 79 98 80 99 
rect 79 113 80 114 
rect 79 116 80 117 
rect 79 119 80 120 
rect 79 145 80 146 
rect 79 161 80 162 
rect 79 163 80 164 
rect 79 167 80 168 
rect 79 193 80 194 
rect 79 200 80 201 
rect 79 214 80 215 
rect 79 216 80 217 
rect 79 227 80 228 
rect 79 230 80 231 
rect 79 243 80 244 
rect 79 261 80 262 
rect 79 276 80 277 
rect 80 19 81 20 
rect 80 54 81 55 
rect 80 67 81 68 
rect 80 86 81 87 
rect 80 88 81 89 
rect 80 98 81 99 
rect 80 113 81 114 
rect 80 116 81 117 
rect 80 119 81 120 
rect 80 144 81 145 
rect 80 145 81 146 
rect 80 161 81 162 
rect 80 163 81 164 
rect 80 167 81 168 
rect 80 193 81 194 
rect 80 200 81 201 
rect 80 214 81 215 
rect 80 216 81 217 
rect 80 227 81 228 
rect 80 229 81 230 
rect 80 230 81 231 
rect 80 243 81 244 
rect 80 261 81 262 
rect 80 276 81 277 
rect 81 19 82 20 
rect 81 21 82 22 
rect 81 22 82 23 
rect 81 23 82 24 
rect 81 24 82 25 
rect 81 54 82 55 
rect 81 67 82 68 
rect 81 86 82 87 
rect 81 88 82 89 
rect 81 98 82 99 
rect 81 113 82 114 
rect 81 116 82 117 
rect 81 119 82 120 
rect 81 127 82 128 
rect 81 128 82 129 
rect 81 129 82 130 
rect 81 130 82 131 
rect 81 131 82 132 
rect 81 132 82 133 
rect 81 133 82 134 
rect 81 134 82 135 
rect 81 135 82 136 
rect 81 136 82 137 
rect 81 137 82 138 
rect 81 138 82 139 
rect 81 139 82 140 
rect 81 140 82 141 
rect 81 141 82 142 
rect 81 142 82 143 
rect 81 143 82 144 
rect 81 144 82 145 
rect 81 161 82 162 
rect 81 163 82 164 
rect 81 167 82 168 
rect 81 193 82 194 
rect 81 200 82 201 
rect 81 214 82 215 
rect 81 216 82 217 
rect 81 227 82 228 
rect 81 229 82 230 
rect 81 231 82 232 
rect 81 232 82 233 
rect 81 233 82 234 
rect 81 234 82 235 
rect 81 235 82 236 
rect 81 236 82 237 
rect 81 243 82 244 
rect 81 261 82 262 
rect 81 276 82 277 
rect 81 303 82 304 
rect 81 304 82 305 
rect 81 305 82 306 
rect 81 306 82 307 
rect 81 307 82 308 
rect 81 308 82 309 
rect 81 309 82 310 
rect 82 19 83 20 
rect 82 54 83 55 
rect 82 67 83 68 
rect 82 71 83 72 
rect 82 72 83 73 
rect 82 73 83 74 
rect 82 74 83 75 
rect 82 86 83 87 
rect 82 88 83 89 
rect 82 98 83 99 
rect 82 113 83 114 
rect 82 116 83 117 
rect 82 119 83 120 
rect 82 161 83 162 
rect 82 163 83 164 
rect 82 167 83 168 
rect 82 193 83 194 
rect 82 200 83 201 
rect 82 214 83 215 
rect 82 216 83 217 
rect 82 227 83 228 
rect 82 243 83 244 
rect 82 261 83 262 
rect 82 276 83 277 
rect 83 19 84 20 
rect 83 54 84 55 
rect 83 67 84 68 
rect 83 86 84 87 
rect 83 88 84 89 
rect 83 98 84 99 
rect 83 113 84 114 
rect 83 116 84 117 
rect 83 119 84 120 
rect 83 135 84 136 
rect 83 136 84 137 
rect 83 137 84 138 
rect 83 138 84 139 
rect 83 161 84 162 
rect 83 163 84 164 
rect 83 167 84 168 
rect 83 193 84 194 
rect 83 200 84 201 
rect 83 214 84 215 
rect 83 216 84 217 
rect 83 227 84 228 
rect 83 243 84 244 
rect 83 261 84 262 
rect 83 276 84 277 
rect 83 278 84 279 
rect 83 279 84 280 
rect 83 280 84 281 
rect 83 281 84 282 
rect 84 19 85 20 
rect 84 54 85 55 
rect 84 67 85 68 
rect 84 86 85 87 
rect 84 98 85 99 
rect 84 113 85 114 
rect 84 116 85 117 
rect 84 119 85 120 
rect 84 161 85 162 
rect 84 163 85 164 
rect 84 193 85 194 
rect 84 214 85 215 
rect 84 216 85 217 
rect 84 227 85 228 
rect 84 243 85 244 
rect 84 261 85 262 
rect 84 276 85 277 
rect 85 19 86 20 
rect 85 54 86 55 
rect 85 67 86 68 
rect 85 86 86 87 
rect 85 98 86 99 
rect 85 100 86 101 
rect 85 101 86 102 
rect 85 102 86 103 
rect 85 103 86 104 
rect 85 104 86 105 
rect 85 105 86 106 
rect 85 106 86 107 
rect 85 107 86 108 
rect 85 108 86 109 
rect 85 109 86 110 
rect 85 113 86 114 
rect 85 116 86 117 
rect 85 119 86 120 
rect 85 161 86 162 
rect 85 163 86 164 
rect 85 193 86 194 
rect 85 197 86 198 
rect 85 198 86 199 
rect 85 199 86 200 
rect 85 200 86 201 
rect 85 201 86 202 
rect 85 202 86 203 
rect 85 203 86 204 
rect 85 204 86 205 
rect 85 205 86 206 
rect 85 206 86 207 
rect 85 207 86 208 
rect 85 208 86 209 
rect 85 209 86 210 
rect 85 210 86 211 
rect 85 211 86 212 
rect 85 212 86 213 
rect 85 213 86 214 
rect 85 214 86 215 
rect 85 216 86 217 
rect 85 227 86 228 
rect 85 243 86 244 
rect 85 261 86 262 
rect 85 276 86 277 
rect 86 19 87 20 
rect 86 54 87 55 
rect 86 67 87 68 
rect 86 86 87 87 
rect 86 98 87 99 
rect 86 113 87 114 
rect 86 116 87 117 
rect 86 119 87 120 
rect 86 145 87 146 
rect 86 161 87 162 
rect 86 163 87 164 
rect 86 193 87 194 
rect 86 197 87 198 
rect 86 216 87 217 
rect 86 227 87 228 
rect 86 243 87 244 
rect 86 261 87 262 
rect 86 276 87 277 
rect 87 19 88 20 
rect 87 51 88 52 
rect 87 54 88 55 
rect 87 67 88 68 
rect 87 69 88 70 
rect 87 86 88 87 
rect 87 98 88 99 
rect 87 113 88 114 
rect 87 116 88 117 
rect 87 119 88 120 
rect 87 145 88 146 
rect 87 161 88 162 
rect 87 163 88 164 
rect 87 193 88 194 
rect 87 197 88 198 
rect 87 216 88 217 
rect 87 227 88 228 
rect 87 243 88 244 
rect 87 261 88 262 
rect 87 276 88 277 
rect 88 19 89 20 
rect 88 40 89 41 
rect 88 51 89 52 
rect 88 54 89 55 
rect 88 67 89 68 
rect 88 69 89 70 
rect 88 86 89 87 
rect 88 98 89 99 
rect 88 113 89 114 
rect 88 116 89 117 
rect 88 119 89 120 
rect 88 134 89 135 
rect 88 135 89 136 
rect 88 136 89 137 
rect 88 137 89 138 
rect 88 145 89 146 
rect 88 161 89 162 
rect 88 163 89 164 
rect 88 193 89 194 
rect 88 197 89 198 
rect 88 216 89 217 
rect 88 227 89 228 
rect 88 243 89 244 
rect 88 261 89 262 
rect 88 276 89 277 
rect 89 19 90 20 
rect 89 40 90 41 
rect 89 51 90 52 
rect 89 54 90 55 
rect 89 67 90 68 
rect 89 69 90 70 
rect 89 86 90 87 
rect 89 98 90 99 
rect 89 102 90 103 
rect 89 113 90 114 
rect 89 116 90 117 
rect 89 119 90 120 
rect 89 131 90 132 
rect 89 145 90 146 
rect 89 161 90 162 
rect 89 163 90 164 
rect 89 193 90 194 
rect 89 197 90 198 
rect 89 216 90 217 
rect 89 225 90 226 
rect 89 227 90 228 
rect 89 243 90 244 
rect 89 261 90 262 
rect 89 276 90 277 
rect 90 19 91 20 
rect 90 40 91 41 
rect 90 51 91 52 
rect 90 54 91 55 
rect 90 67 91 68 
rect 90 69 91 70 
rect 90 86 91 87 
rect 90 98 91 99 
rect 90 102 91 103 
rect 90 113 91 114 
rect 90 116 91 117 
rect 90 119 91 120 
rect 90 131 91 132 
rect 90 145 91 146 
rect 90 161 91 162 
rect 90 163 91 164 
rect 90 193 91 194 
rect 90 196 91 197 
rect 90 197 91 198 
rect 90 216 91 217 
rect 90 225 91 226 
rect 90 227 91 228 
rect 90 243 91 244 
rect 90 261 91 262 
rect 90 276 91 277 
rect 91 19 92 20 
rect 91 40 92 41 
rect 91 51 92 52 
rect 91 54 92 55 
rect 91 67 92 68 
rect 91 69 92 70 
rect 91 86 92 87 
rect 91 98 92 99 
rect 91 102 92 103 
rect 91 113 92 114 
rect 91 116 92 117 
rect 91 119 92 120 
rect 91 131 92 132 
rect 91 145 92 146 
rect 91 161 92 162 
rect 91 163 92 164 
rect 91 193 92 194 
rect 91 216 92 217 
rect 91 225 92 226 
rect 91 227 92 228 
rect 91 243 92 244 
rect 91 261 92 262 
rect 91 276 92 277 
rect 92 19 93 20 
rect 92 40 93 41 
rect 92 51 93 52 
rect 92 54 93 55 
rect 92 67 93 68 
rect 92 69 93 70 
rect 92 86 93 87 
rect 92 98 93 99 
rect 92 102 93 103 
rect 92 113 93 114 
rect 92 116 93 117 
rect 92 119 93 120 
rect 92 131 93 132 
rect 92 145 93 146 
rect 92 161 93 162 
rect 92 163 93 164 
rect 92 193 93 194 
rect 92 216 93 217 
rect 92 225 93 226 
rect 92 227 93 228 
rect 92 243 93 244 
rect 92 261 93 262 
rect 92 276 93 277 
rect 93 19 94 20 
rect 93 40 94 41 
rect 93 51 94 52 
rect 93 54 94 55 
rect 93 65 94 66 
rect 93 67 94 68 
rect 93 69 94 70 
rect 93 86 94 87 
rect 93 98 94 99 
rect 93 102 94 103 
rect 93 113 94 114 
rect 93 116 94 117 
rect 93 119 94 120 
rect 93 131 94 132 
rect 93 145 94 146 
rect 93 161 94 162 
rect 93 163 94 164 
rect 93 193 94 194 
rect 93 216 94 217 
rect 93 225 94 226 
rect 93 227 94 228 
rect 93 243 94 244 
rect 93 261 94 262 
rect 93 276 94 277 
rect 94 19 95 20 
rect 94 20 95 21 
rect 94 40 95 41 
rect 94 51 95 52 
rect 94 54 95 55 
rect 94 65 95 66 
rect 94 67 95 68 
rect 94 69 95 70 
rect 94 86 95 87 
rect 94 98 95 99 
rect 94 102 95 103 
rect 94 113 95 114 
rect 94 116 95 117 
rect 94 119 95 120 
rect 94 131 95 132 
rect 94 145 95 146 
rect 94 161 95 162 
rect 94 163 95 164 
rect 94 193 95 194 
rect 94 216 95 217 
rect 94 225 95 226 
rect 94 227 95 228 
rect 94 243 95 244 
rect 94 261 95 262 
rect 94 276 95 277 
rect 95 20 96 21 
rect 95 40 96 41 
rect 95 51 96 52 
rect 95 54 96 55 
rect 95 65 96 66 
rect 95 67 96 68 
rect 95 69 96 70 
rect 95 84 96 85 
rect 95 86 96 87 
rect 95 98 96 99 
rect 95 100 96 101 
rect 95 102 96 103 
rect 95 113 96 114 
rect 95 116 96 117 
rect 95 119 96 120 
rect 95 131 96 132 
rect 95 145 96 146 
rect 95 161 96 162 
rect 95 163 96 164 
rect 95 193 96 194 
rect 95 216 96 217 
rect 95 225 96 226 
rect 95 227 96 228 
rect 95 243 96 244 
rect 95 261 96 262 
rect 95 276 96 277 
rect 96 20 97 21 
rect 96 40 97 41 
rect 96 51 97 52 
rect 96 54 97 55 
rect 96 65 97 66 
rect 96 67 97 68 
rect 96 69 97 70 
rect 96 84 97 85 
rect 96 86 97 87 
rect 96 88 97 89 
rect 96 98 97 99 
rect 96 100 97 101 
rect 96 102 97 103 
rect 96 113 97 114 
rect 96 116 97 117 
rect 96 119 97 120 
rect 96 131 97 132 
rect 96 144 97 145 
rect 96 145 97 146 
rect 96 161 97 162 
rect 96 163 97 164 
rect 96 193 97 194 
rect 96 216 97 217 
rect 96 217 97 218 
rect 96 225 97 226 
rect 96 227 97 228 
rect 96 243 97 244 
rect 96 246 97 247 
rect 96 247 97 248 
rect 96 248 97 249 
rect 96 249 97 250 
rect 96 261 97 262 
rect 96 263 97 264 
rect 96 276 97 277 
rect 97 40 98 41 
rect 97 51 98 52 
rect 97 54 98 55 
rect 97 65 98 66 
rect 97 67 98 68 
rect 97 84 98 85 
rect 97 86 98 87 
rect 97 88 98 89 
rect 97 98 98 99 
rect 97 100 98 101 
rect 97 102 98 103 
rect 97 113 98 114 
rect 97 116 98 117 
rect 97 119 98 120 
rect 97 131 98 132 
rect 97 144 98 145 
rect 97 160 98 161 
rect 97 161 98 162 
rect 97 163 98 164 
rect 97 193 98 194 
rect 97 217 98 218 
rect 97 218 98 219 
rect 97 225 98 226 
rect 97 227 98 228 
rect 97 243 98 244 
rect 97 261 98 262 
rect 97 263 98 264 
rect 97 276 98 277 
rect 97 303 98 304 
rect 97 304 98 305 
rect 97 305 98 306 
rect 97 306 98 307 
rect 98 40 99 41 
rect 98 51 99 52 
rect 98 54 99 55 
rect 98 65 99 66 
rect 98 67 99 68 
rect 98 84 99 85 
rect 98 86 99 87 
rect 98 88 99 89 
rect 98 98 99 99 
rect 98 100 99 101 
rect 98 102 99 103 
rect 98 113 99 114 
rect 98 116 99 117 
rect 98 119 99 120 
rect 98 131 99 132 
rect 98 163 99 164 
rect 98 183 99 184 
rect 98 184 99 185 
rect 98 185 99 186 
rect 98 186 99 187 
rect 98 187 99 188 
rect 98 188 99 189 
rect 98 189 99 190 
rect 98 193 99 194 
rect 98 198 99 199 
rect 98 199 99 200 
rect 98 200 99 201 
rect 98 201 99 202 
rect 98 225 99 226 
rect 98 227 99 228 
rect 98 243 99 244 
rect 98 261 99 262 
rect 98 263 99 264 
rect 98 276 99 277 
rect 99 40 100 41 
rect 99 51 100 52 
rect 99 54 100 55 
rect 99 65 100 66 
rect 99 67 100 68 
rect 99 84 100 85 
rect 99 86 100 87 
rect 99 88 100 89 
rect 99 98 100 99 
rect 99 100 100 101 
rect 99 102 100 103 
rect 99 113 100 114 
rect 99 116 100 117 
rect 99 131 100 132 
rect 99 163 100 164 
rect 99 182 100 183 
rect 99 183 100 184 
rect 99 193 100 194 
rect 99 197 100 198 
rect 99 198 100 199 
rect 99 225 100 226 
rect 99 227 100 228 
rect 99 243 100 244 
rect 99 261 100 262 
rect 99 263 100 264 
rect 99 276 100 277 
rect 100 40 101 41 
rect 100 51 101 52 
rect 100 54 101 55 
rect 100 65 101 66 
rect 100 67 101 68 
rect 100 88 101 89 
rect 100 100 101 101 
rect 100 113 101 114 
rect 100 116 101 117 
rect 100 131 101 132 
rect 100 163 101 164 
rect 100 182 101 183 
rect 100 193 101 194 
rect 100 197 101 198 
rect 100 225 101 226 
rect 100 227 101 228 
rect 100 243 101 244 
rect 100 261 101 262 
rect 100 263 101 264 
rect 100 276 101 277 
rect 101 40 102 41 
rect 101 51 102 52 
rect 101 54 102 55 
rect 101 65 102 66 
rect 101 67 102 68 
rect 101 88 102 89 
rect 101 100 102 101 
rect 101 113 102 114 
rect 101 116 102 117 
rect 101 131 102 132 
rect 101 163 102 164 
rect 101 177 102 178 
rect 101 182 102 183 
rect 101 184 102 185 
rect 101 193 102 194 
rect 101 195 102 196 
rect 101 197 102 198 
rect 101 199 102 200 
rect 101 225 102 226 
rect 101 227 102 228 
rect 101 243 102 244 
rect 101 261 102 262 
rect 101 263 102 264 
rect 101 276 102 277 
rect 102 40 103 41 
rect 102 51 103 52 
rect 102 54 103 55 
rect 102 65 103 66 
rect 102 67 103 68 
rect 102 88 103 89 
rect 102 100 103 101 
rect 102 113 103 114 
rect 102 131 103 132 
rect 102 133 103 134 
rect 102 134 103 135 
rect 102 135 103 136 
rect 102 136 103 137 
rect 102 137 103 138 
rect 102 138 103 139 
rect 102 139 103 140 
rect 102 140 103 141 
rect 102 141 103 142 
rect 102 142 103 143 
rect 102 143 103 144 
rect 102 144 103 145 
rect 102 145 103 146 
rect 102 163 103 164 
rect 102 177 103 178 
rect 102 182 103 183 
rect 102 184 103 185 
rect 102 193 103 194 
rect 102 195 103 196 
rect 102 197 103 198 
rect 102 199 103 200 
rect 102 211 103 212 
rect 102 212 103 213 
rect 102 213 103 214 
rect 102 214 103 215 
rect 102 215 103 216 
rect 102 216 103 217 
rect 102 217 103 218 
rect 102 218 103 219 
rect 102 225 103 226 
rect 102 227 103 228 
rect 102 243 103 244 
rect 102 261 103 262 
rect 102 263 103 264 
rect 102 276 103 277 
rect 103 40 104 41 
rect 103 51 104 52 
rect 103 54 104 55 
rect 103 65 104 66 
rect 103 67 104 68 
rect 103 88 104 89 
rect 103 100 104 101 
rect 103 113 104 114 
rect 103 131 104 132 
rect 103 145 104 146 
rect 103 146 104 147 
rect 103 163 104 164 
rect 103 177 104 178 
rect 103 182 104 183 
rect 103 184 104 185 
rect 103 193 104 194 
rect 103 195 104 196 
rect 103 197 104 198 
rect 103 199 104 200 
rect 103 210 104 211 
rect 103 211 104 212 
rect 103 225 104 226 
rect 103 227 104 228 
rect 103 243 104 244 
rect 103 261 104 262 
rect 103 263 104 264 
rect 103 276 104 277 
rect 104 40 105 41 
rect 104 51 105 52 
rect 104 54 105 55 
rect 104 65 105 66 
rect 104 67 105 68 
rect 104 88 105 89 
rect 104 100 105 101 
rect 104 113 105 114 
rect 104 114 105 115 
rect 104 115 105 116 
rect 104 116 105 117 
rect 104 117 105 118 
rect 104 118 105 119 
rect 104 131 105 132 
rect 104 132 105 133 
rect 104 133 105 134 
rect 104 134 105 135 
rect 104 135 105 136 
rect 104 136 105 137 
rect 104 137 105 138 
rect 104 138 105 139 
rect 104 139 105 140 
rect 104 140 105 141 
rect 104 141 105 142 
rect 104 142 105 143 
rect 104 143 105 144 
rect 104 144 105 145 
rect 104 146 105 147 
rect 104 147 105 148 
rect 104 163 105 164 
rect 104 177 105 178 
rect 104 182 105 183 
rect 104 184 105 185 
rect 104 193 105 194 
rect 104 195 105 196 
rect 104 197 105 198 
rect 104 199 105 200 
rect 104 210 105 211 
rect 104 213 105 214 
rect 104 214 105 215 
rect 104 215 105 216 
rect 104 216 105 217 
rect 104 217 105 218 
rect 104 218 105 219 
rect 104 225 105 226 
rect 104 227 105 228 
rect 104 243 105 244 
rect 104 261 105 262 
rect 104 263 105 264 
rect 104 276 105 277 
rect 105 40 106 41 
rect 105 51 106 52 
rect 105 54 106 55 
rect 105 65 106 66 
rect 105 67 106 68 
rect 105 88 106 89 
rect 105 100 106 101 
rect 105 144 106 145 
rect 105 145 106 146 
rect 105 147 106 148 
rect 105 163 106 164 
rect 105 177 106 178 
rect 105 182 106 183 
rect 105 184 106 185 
rect 105 193 106 194 
rect 105 195 106 196 
rect 105 197 106 198 
rect 105 199 106 200 
rect 105 210 106 211 
rect 105 225 106 226 
rect 105 227 106 228 
rect 105 243 106 244 
rect 105 261 106 262 
rect 105 263 106 264 
rect 105 276 106 277 
rect 106 40 107 41 
rect 106 51 107 52 
rect 106 54 107 55 
rect 106 65 107 66 
rect 106 67 107 68 
rect 106 88 107 89 
rect 106 100 107 101 
rect 106 145 107 146 
rect 106 147 107 148 
rect 106 163 107 164 
rect 106 177 107 178 
rect 106 182 107 183 
rect 106 184 107 185 
rect 106 193 107 194 
rect 106 195 107 196 
rect 106 197 107 198 
rect 106 199 107 200 
rect 106 210 107 211 
rect 106 225 107 226 
rect 106 227 107 228 
rect 106 243 107 244 
rect 106 261 107 262 
rect 106 263 107 264 
rect 106 276 107 277 
rect 107 40 108 41 
rect 107 51 108 52 
rect 107 54 108 55 
rect 107 65 108 66 
rect 107 67 108 68 
rect 107 88 108 89 
rect 107 100 108 101 
rect 107 145 108 146 
rect 107 147 108 148 
rect 107 163 108 164 
rect 107 177 108 178 
rect 107 182 108 183 
rect 107 184 108 185 
rect 107 193 108 194 
rect 107 197 108 198 
rect 107 199 108 200 
rect 107 210 108 211 
rect 107 225 108 226 
rect 107 227 108 228 
rect 107 243 108 244 
rect 107 261 108 262 
rect 107 263 108 264 
rect 107 276 108 277 
rect 108 40 109 41 
rect 108 51 109 52 
rect 108 54 109 55 
rect 108 65 109 66 
rect 108 67 109 68 
rect 108 88 109 89 
rect 108 100 109 101 
rect 108 145 109 146 
rect 108 147 109 148 
rect 108 163 109 164 
rect 108 177 109 178 
rect 108 182 109 183 
rect 108 184 109 185 
rect 108 193 109 194 
rect 108 197 109 198 
rect 108 199 109 200 
rect 108 210 109 211 
rect 108 225 109 226 
rect 108 227 109 228 
rect 108 243 109 244 
rect 108 261 109 262 
rect 108 263 109 264 
rect 108 276 109 277 
rect 109 40 110 41 
rect 109 51 110 52 
rect 109 54 110 55 
rect 109 65 110 66 
rect 109 67 110 68 
rect 109 88 110 89 
rect 109 100 110 101 
rect 109 145 110 146 
rect 109 147 110 148 
rect 109 163 110 164 
rect 109 177 110 178 
rect 109 182 110 183 
rect 109 184 110 185 
rect 109 193 110 194 
rect 109 197 110 198 
rect 109 199 110 200 
rect 109 210 110 211 
rect 109 225 110 226 
rect 109 227 110 228 
rect 109 243 110 244 
rect 109 261 110 262 
rect 109 263 110 264 
rect 109 276 110 277 
rect 110 40 111 41 
rect 110 51 111 52 
rect 110 54 111 55 
rect 110 65 111 66 
rect 110 67 111 68 
rect 110 88 111 89 
rect 110 100 111 101 
rect 110 145 111 146 
rect 110 147 111 148 
rect 110 148 111 149 
rect 110 163 111 164 
rect 110 177 111 178 
rect 110 182 111 183 
rect 110 184 111 185 
rect 110 193 111 194 
rect 110 197 111 198 
rect 110 199 111 200 
rect 110 210 111 211 
rect 110 225 111 226 
rect 110 227 111 228 
rect 110 243 111 244 
rect 110 261 111 262 
rect 110 263 111 264 
rect 110 276 111 277 
rect 111 40 112 41 
rect 111 48 112 49 
rect 111 49 112 50 
rect 111 50 112 51 
rect 111 51 112 52 
rect 111 54 112 55 
rect 111 65 112 66 
rect 111 67 112 68 
rect 111 88 112 89 
rect 111 100 112 101 
rect 111 145 112 146 
rect 111 163 112 164 
rect 111 177 112 178 
rect 111 182 112 183 
rect 111 184 112 185 
rect 111 193 112 194 
rect 111 197 112 198 
rect 111 199 112 200 
rect 111 210 112 211 
rect 111 225 112 226 
rect 111 227 112 228 
rect 111 228 112 229 
rect 111 243 112 244 
rect 111 261 112 262 
rect 111 263 112 264 
rect 111 276 112 277 
rect 112 40 113 41 
rect 112 48 113 49 
rect 112 54 113 55 
rect 112 65 113 66 
rect 112 67 113 68 
rect 112 69 113 70 
rect 112 88 113 89 
rect 112 100 113 101 
rect 112 145 113 146 
rect 112 163 113 164 
rect 112 177 113 178 
rect 112 184 113 185 
rect 112 193 113 194 
rect 112 197 113 198 
rect 112 199 113 200 
rect 112 210 113 211 
rect 112 225 113 226 
rect 112 226 113 227 
rect 112 228 113 229 
rect 112 241 113 242 
rect 112 243 113 244 
rect 112 261 113 262 
rect 112 263 113 264 
rect 112 276 113 277 
rect 113 40 114 41 
rect 113 48 114 49 
rect 113 54 114 55 
rect 113 65 114 66 
rect 113 67 114 68 
rect 113 69 114 70 
rect 113 71 114 72 
rect 113 88 114 89 
rect 113 100 114 101 
rect 113 134 114 135 
rect 113 135 114 136 
rect 113 136 114 137 
rect 113 137 114 138 
rect 113 145 114 146 
rect 113 163 114 164 
rect 113 177 114 178 
rect 113 184 114 185 
rect 113 193 114 194 
rect 113 197 114 198 
rect 113 199 114 200 
rect 113 210 114 211 
rect 113 214 114 215 
rect 113 215 114 216 
rect 113 216 114 217 
rect 113 217 114 218 
rect 113 218 114 219 
rect 113 219 114 220 
rect 113 220 114 221 
rect 113 221 114 222 
rect 113 222 114 223 
rect 113 223 114 224 
rect 113 226 114 227 
rect 113 228 114 229 
rect 113 241 114 242 
rect 113 243 114 244 
rect 113 245 114 246 
rect 113 246 114 247 
rect 113 247 114 248 
rect 113 248 114 249 
rect 113 261 114 262 
rect 113 263 114 264 
rect 113 276 114 277 
rect 113 277 114 278 
rect 113 278 114 279 
rect 113 279 114 280 
rect 113 280 114 281 
rect 113 281 114 282 
rect 114 36 115 37 
rect 114 38 115 39 
rect 114 40 115 41 
rect 114 48 115 49 
rect 114 50 115 51 
rect 114 52 115 53 
rect 114 54 115 55 
rect 114 56 115 57 
rect 114 65 115 66 
rect 114 67 115 68 
rect 114 69 115 70 
rect 114 71 115 72 
rect 114 88 115 89 
rect 114 100 115 101 
rect 114 145 115 146 
rect 114 163 115 164 
rect 114 177 115 178 
rect 114 184 115 185 
rect 114 193 115 194 
rect 114 197 115 198 
rect 114 199 115 200 
rect 114 210 115 211 
rect 114 214 115 215 
rect 114 226 115 227 
rect 114 228 115 229 
rect 114 241 115 242 
rect 114 243 115 244 
rect 114 261 115 262 
rect 114 263 115 264 
rect 115 16 116 17 
rect 115 17 116 18 
rect 115 18 116 19 
rect 115 19 116 20 
rect 115 20 116 21 
rect 115 21 116 22 
rect 115 22 116 23 
rect 115 23 116 24 
rect 115 24 116 25 
rect 115 36 116 37 
rect 115 38 116 39 
rect 115 40 116 41 
rect 115 48 116 49 
rect 115 50 116 51 
rect 115 52 116 53 
rect 115 54 116 55 
rect 115 56 116 57 
rect 115 65 116 66 
rect 115 67 116 68 
rect 115 69 116 70 
rect 115 71 116 72 
rect 115 84 116 85 
rect 115 88 116 89 
rect 115 100 116 101 
rect 115 132 116 133 
rect 115 133 116 134 
rect 115 134 116 135 
rect 115 135 116 136 
rect 115 136 116 137 
rect 115 137 116 138 
rect 115 145 116 146 
rect 115 163 116 164 
rect 115 177 116 178 
rect 115 184 116 185 
rect 115 193 116 194 
rect 115 197 116 198 
rect 115 199 116 200 
rect 115 210 116 211 
rect 115 214 116 215 
rect 115 226 116 227 
rect 115 228 116 229 
rect 115 241 116 242 
rect 115 243 116 244 
rect 115 246 116 247 
rect 115 247 116 248 
rect 115 248 116 249 
rect 115 249 116 250 
rect 115 261 116 262 
rect 115 263 116 264 
rect 116 36 117 37 
rect 116 38 117 39 
rect 116 40 117 41 
rect 116 48 117 49 
rect 116 50 117 51 
rect 116 52 117 53 
rect 116 54 117 55 
rect 116 56 117 57 
rect 116 65 117 66 
rect 116 67 117 68 
rect 116 69 117 70 
rect 116 71 117 72 
rect 116 84 117 85 
rect 116 86 117 87 
rect 116 88 117 89 
rect 116 100 117 101 
rect 116 145 117 146 
rect 116 163 117 164 
rect 116 177 117 178 
rect 116 184 117 185 
rect 116 193 117 194 
rect 116 197 117 198 
rect 116 199 117 200 
rect 116 210 117 211 
rect 116 214 117 215 
rect 116 226 117 227 
rect 116 228 117 229 
rect 116 241 117 242 
rect 116 243 117 244 
rect 117 36 118 37 
rect 117 38 118 39 
rect 117 40 118 41 
rect 117 48 118 49 
rect 117 50 118 51 
rect 117 52 118 53 
rect 117 54 118 55 
rect 117 56 118 57 
rect 117 65 118 66 
rect 117 67 118 68 
rect 117 69 118 70 
rect 117 71 118 72 
rect 117 84 118 85 
rect 117 86 118 87 
rect 117 88 118 89 
rect 117 100 118 101 
rect 117 145 118 146 
rect 117 163 118 164 
rect 117 177 118 178 
rect 117 181 118 182 
rect 117 184 118 185 
rect 117 193 118 194 
rect 117 197 118 198 
rect 117 199 118 200 
rect 117 210 118 211 
rect 117 214 118 215 
rect 117 226 118 227 
rect 117 228 118 229 
rect 117 241 118 242 
rect 117 243 118 244 
rect 118 37 119 38 
rect 118 38 119 39 
rect 118 40 119 41 
rect 118 48 119 49 
rect 118 50 119 51 
rect 118 52 119 53 
rect 118 54 119 55 
rect 118 56 119 57 
rect 118 65 119 66 
rect 118 67 119 68 
rect 118 69 119 70 
rect 118 71 119 72 
rect 118 84 119 85 
rect 118 86 119 87 
rect 118 88 119 89 
rect 118 97 119 98 
rect 118 100 119 101 
rect 118 102 119 103 
rect 118 104 119 105 
rect 118 145 119 146 
rect 118 163 119 164 
rect 118 177 119 178 
rect 118 181 119 182 
rect 118 184 119 185 
rect 118 193 119 194 
rect 118 195 119 196 
rect 118 197 119 198 
rect 118 199 119 200 
rect 118 210 119 211 
rect 118 214 119 215 
rect 118 228 119 229 
rect 118 241 119 242 
rect 118 243 119 244 
rect 118 276 119 277 
rect 119 36 120 37 
rect 119 37 120 38 
rect 119 40 120 41 
rect 119 48 120 49 
rect 119 50 120 51 
rect 119 52 120 53 
rect 119 54 120 55 
rect 119 56 120 57 
rect 119 65 120 66 
rect 119 67 120 68 
rect 119 69 120 70 
rect 119 71 120 72 
rect 119 84 120 85 
rect 119 86 120 87 
rect 119 88 120 89 
rect 119 97 120 98 
rect 119 99 120 100 
rect 119 100 120 101 
rect 119 102 120 103 
rect 119 104 120 105 
rect 119 145 120 146 
rect 119 163 120 164 
rect 119 177 120 178 
rect 119 181 120 182 
rect 119 184 120 185 
rect 119 193 120 194 
rect 119 195 120 196 
rect 119 197 120 198 
rect 119 199 120 200 
rect 119 210 120 211 
rect 119 214 120 215 
rect 119 228 120 229 
rect 119 241 120 242 
rect 119 243 120 244 
rect 119 276 120 277 
rect 119 278 120 279 
rect 119 279 120 280 
rect 119 280 120 281 
rect 119 281 120 282 
rect 120 36 121 37 
rect 120 40 121 41 
rect 120 48 121 49 
rect 120 50 121 51 
rect 120 52 121 53 
rect 120 54 121 55 
rect 120 56 121 57 
rect 120 65 121 66 
rect 120 67 121 68 
rect 120 69 121 70 
rect 120 71 121 72 
rect 120 84 121 85 
rect 120 86 121 87 
rect 120 88 121 89 
rect 120 97 121 98 
rect 120 99 121 100 
rect 120 102 121 103 
rect 120 104 121 105 
rect 120 145 121 146 
rect 120 163 121 164 
rect 120 177 121 178 
rect 120 181 121 182 
rect 120 184 121 185 
rect 120 193 121 194 
rect 120 195 121 196 
rect 120 197 121 198 
rect 120 199 121 200 
rect 120 210 121 211 
rect 120 214 121 215 
rect 120 228 121 229 
rect 120 241 121 242 
rect 120 243 121 244 
rect 120 276 121 277 
rect 121 36 122 37 
rect 121 40 122 41 
rect 121 48 122 49 
rect 121 50 122 51 
rect 121 52 122 53 
rect 121 54 122 55 
rect 121 56 122 57 
rect 121 65 122 66 
rect 121 67 122 68 
rect 121 69 122 70 
rect 121 71 122 72 
rect 121 84 122 85 
rect 121 86 122 87 
rect 121 88 122 89 
rect 121 97 122 98 
rect 121 99 122 100 
rect 121 102 122 103 
rect 121 104 122 105 
rect 121 145 122 146 
rect 121 163 122 164 
rect 121 177 122 178 
rect 121 184 122 185 
rect 121 193 122 194 
rect 121 195 122 196 
rect 121 199 122 200 
rect 121 210 122 211 
rect 121 214 122 215 
rect 121 228 122 229 
rect 121 241 122 242 
rect 121 243 122 244 
rect 121 276 122 277 
rect 122 36 123 37 
rect 122 40 123 41 
rect 122 50 123 51 
rect 122 52 123 53 
rect 122 54 123 55 
rect 122 56 123 57 
rect 122 65 123 66 
rect 122 67 123 68 
rect 122 71 123 72 
rect 122 84 123 85 
rect 122 86 123 87 
rect 122 88 123 89 
rect 122 97 123 98 
rect 122 99 123 100 
rect 122 102 123 103 
rect 122 104 123 105 
rect 122 145 123 146 
rect 122 163 123 164 
rect 122 177 123 178 
rect 122 184 123 185 
rect 122 193 123 194 
rect 122 199 123 200 
rect 122 210 123 211 
rect 122 214 123 215 
rect 122 276 123 277 
rect 123 36 124 37 
rect 123 40 124 41 
rect 123 50 124 51 
rect 123 52 124 53 
rect 123 54 124 55 
rect 123 56 124 57 
rect 123 65 124 66 
rect 123 67 124 68 
rect 123 71 124 72 
rect 123 84 124 85 
rect 123 86 124 87 
rect 123 88 124 89 
rect 123 97 124 98 
rect 123 99 124 100 
rect 123 102 124 103 
rect 123 104 124 105 
rect 123 145 124 146 
rect 123 163 124 164 
rect 123 177 124 178 
rect 123 184 124 185 
rect 123 193 124 194 
rect 123 199 124 200 
rect 123 210 124 211 
rect 123 214 124 215 
rect 123 276 124 277 
rect 124 36 125 37 
rect 124 40 125 41 
rect 124 50 125 51 
rect 124 52 125 53 
rect 124 54 125 55 
rect 124 56 125 57 
rect 124 65 125 66 
rect 124 67 125 68 
rect 124 71 125 72 
rect 124 84 125 85 
rect 124 86 125 87 
rect 124 88 125 89 
rect 124 97 125 98 
rect 124 99 125 100 
rect 124 102 125 103 
rect 124 104 125 105 
rect 124 145 125 146 
rect 124 163 125 164 
rect 124 177 125 178 
rect 124 184 125 185 
rect 124 193 125 194 
rect 124 199 125 200 
rect 124 210 125 211 
rect 124 214 125 215 
rect 124 276 125 277 
rect 124 289 125 290 
rect 124 290 125 291 
rect 124 291 125 292 
rect 124 292 125 293 
rect 125 36 126 37 
rect 125 40 126 41 
rect 125 50 126 51 
rect 125 52 126 53 
rect 125 54 126 55 
rect 125 56 126 57 
rect 125 65 126 66 
rect 125 67 126 68 
rect 125 71 126 72 
rect 125 84 126 85 
rect 125 86 126 87 
rect 125 88 126 89 
rect 125 97 126 98 
rect 125 99 126 100 
rect 125 102 126 103 
rect 125 104 126 105 
rect 125 145 126 146 
rect 125 163 126 164 
rect 125 166 126 167 
rect 125 167 126 168 
rect 125 177 126 178 
rect 125 184 126 185 
rect 125 193 126 194 
rect 125 199 126 200 
rect 125 210 126 211 
rect 125 214 126 215 
rect 125 276 126 277 
rect 125 289 126 290 
rect 126 36 127 37 
rect 126 40 127 41 
rect 126 50 127 51 
rect 126 52 127 53 
rect 126 54 127 55 
rect 126 56 127 57 
rect 126 65 127 66 
rect 126 67 127 68 
rect 126 71 127 72 
rect 126 84 127 85 
rect 126 86 127 87 
rect 126 88 127 89 
rect 126 97 127 98 
rect 126 99 127 100 
rect 126 102 127 103 
rect 126 104 127 105 
rect 126 145 127 146 
rect 126 163 127 164 
rect 126 167 127 168 
rect 126 177 127 178 
rect 126 184 127 185 
rect 126 193 127 194 
rect 126 199 127 200 
rect 126 210 127 211 
rect 126 214 127 215 
rect 126 276 127 277 
rect 126 289 127 290 
rect 127 36 128 37 
rect 127 40 128 41 
rect 127 50 128 51 
rect 127 52 128 53 
rect 127 54 128 55 
rect 127 56 128 57 
rect 127 65 128 66 
rect 127 67 128 68 
rect 127 71 128 72 
rect 127 84 128 85 
rect 127 86 128 87 
rect 127 88 128 89 
rect 127 97 128 98 
rect 127 99 128 100 
rect 127 102 128 103 
rect 127 104 128 105 
rect 127 145 128 146 
rect 127 163 128 164 
rect 127 167 128 168 
rect 127 177 128 178 
rect 127 184 128 185 
rect 127 193 128 194 
rect 127 199 128 200 
rect 127 210 128 211 
rect 127 214 128 215 
rect 127 276 128 277 
rect 127 289 128 290 
rect 128 32 129 33 
rect 128 33 129 34 
rect 128 34 129 35 
rect 128 35 129 36 
rect 128 36 129 37 
rect 128 40 129 41 
rect 128 50 129 51 
rect 128 52 129 53 
rect 128 54 129 55 
rect 128 56 129 57 
rect 128 65 129 66 
rect 128 67 129 68 
rect 128 71 129 72 
rect 128 84 129 85 
rect 128 86 129 87 
rect 128 88 129 89 
rect 128 97 129 98 
rect 128 99 129 100 
rect 128 102 129 103 
rect 128 104 129 105 
rect 128 145 129 146 
rect 128 163 129 164 
rect 128 167 129 168 
rect 128 177 129 178 
rect 128 184 129 185 
rect 128 193 129 194 
rect 128 199 129 200 
rect 128 210 129 211 
rect 128 214 129 215 
rect 128 257 129 258 
rect 128 261 129 262 
rect 128 276 129 277 
rect 128 288 129 289 
rect 128 289 129 290 
rect 129 16 130 17 
rect 129 17 130 18 
rect 129 18 130 19 
rect 129 19 130 20 
rect 129 20 130 21 
rect 129 21 130 22 
rect 129 22 130 23 
rect 129 23 130 24 
rect 129 24 130 25 
rect 129 25 130 26 
rect 129 27 130 28 
rect 129 28 130 29 
rect 129 29 130 30 
rect 129 30 130 31 
rect 129 31 130 32 
rect 129 32 130 33 
rect 129 40 130 41 
rect 129 48 130 49 
rect 129 50 130 51 
rect 129 52 130 53 
rect 129 54 130 55 
rect 129 56 130 57 
rect 129 65 130 66 
rect 129 67 130 68 
rect 129 71 130 72 
rect 129 73 130 74 
rect 129 74 130 75 
rect 129 75 130 76 
rect 129 76 130 77 
rect 129 77 130 78 
rect 129 78 130 79 
rect 129 79 130 80 
rect 129 80 130 81 
rect 129 81 130 82 
rect 129 84 130 85 
rect 129 86 130 87 
rect 129 88 130 89 
rect 129 97 130 98 
rect 129 99 130 100 
rect 129 102 130 103 
rect 129 104 130 105 
rect 129 145 130 146 
rect 129 163 130 164 
rect 129 167 130 168 
rect 129 177 130 178 
rect 129 184 130 185 
rect 129 193 130 194 
rect 129 199 130 200 
rect 129 210 130 211 
rect 129 214 130 215 
rect 129 240 130 241 
rect 129 241 130 242 
rect 129 242 130 243 
rect 129 243 130 244 
rect 129 244 130 245 
rect 129 245 130 246 
rect 129 246 130 247 
rect 129 247 130 248 
rect 129 248 130 249 
rect 129 249 130 250 
rect 129 250 130 251 
rect 129 251 130 252 
rect 129 252 130 253 
rect 129 257 130 258 
rect 129 261 130 262 
rect 129 276 130 277 
rect 129 278 130 279 
rect 129 279 130 280 
rect 129 280 130 281 
rect 129 281 130 282 
rect 129 282 130 283 
rect 129 283 130 284 
rect 129 284 130 285 
rect 129 285 130 286 
rect 129 286 130 287 
rect 129 287 130 288 
rect 129 288 130 289 
rect 130 26 131 27 
rect 130 27 131 28 
rect 130 40 131 41 
rect 130 48 131 49 
rect 130 50 131 51 
rect 130 52 131 53 
rect 130 54 131 55 
rect 130 56 131 57 
rect 130 65 131 66 
rect 130 67 131 68 
rect 130 71 131 72 
rect 130 81 131 82 
rect 130 84 131 85 
rect 130 86 131 87 
rect 130 88 131 89 
rect 130 97 131 98 
rect 130 99 131 100 
rect 130 102 131 103 
rect 130 104 131 105 
rect 130 112 131 113 
rect 130 113 131 114 
rect 130 114 131 115 
rect 130 115 131 116 
rect 130 116 131 117 
rect 130 117 131 118 
rect 130 118 131 119 
rect 130 119 131 120 
rect 130 120 131 121 
rect 130 121 131 122 
rect 130 122 131 123 
rect 130 123 131 124 
rect 130 124 131 125 
rect 130 125 131 126 
rect 130 126 131 127 
rect 130 127 131 128 
rect 130 128 131 129 
rect 130 129 131 130 
rect 130 130 131 131 
rect 130 131 131 132 
rect 130 132 131 133 
rect 130 133 131 134 
rect 130 134 131 135 
rect 130 135 131 136 
rect 130 136 131 137 
rect 130 137 131 138 
rect 130 138 131 139 
rect 130 139 131 140 
rect 130 140 131 141 
rect 130 145 131 146 
rect 130 163 131 164 
rect 130 167 131 168 
rect 130 177 131 178 
rect 130 184 131 185 
rect 130 193 131 194 
rect 130 199 131 200 
rect 130 210 131 211 
rect 130 214 131 215 
rect 130 252 131 253 
rect 130 257 131 258 
rect 130 261 131 262 
rect 130 276 131 277 
rect 130 278 131 279 
rect 131 18 132 19 
rect 131 19 132 20 
rect 131 20 132 21 
rect 131 21 132 22 
rect 131 22 132 23 
rect 131 23 132 24 
rect 131 24 132 25 
rect 131 25 132 26 
rect 131 26 132 27 
rect 131 40 132 41 
rect 131 48 132 49 
rect 131 50 132 51 
rect 131 52 132 53 
rect 131 54 132 55 
rect 131 56 132 57 
rect 131 65 132 66 
rect 131 67 132 68 
rect 131 71 132 72 
rect 131 81 132 82 
rect 131 84 132 85 
rect 131 86 132 87 
rect 131 88 132 89 
rect 131 97 132 98 
rect 131 99 132 100 
rect 131 102 132 103 
rect 131 104 132 105 
rect 131 145 132 146 
rect 131 163 132 164 
rect 131 167 132 168 
rect 131 177 132 178 
rect 131 184 132 185 
rect 131 193 132 194 
rect 131 199 132 200 
rect 131 210 132 211 
rect 131 214 132 215 
rect 131 252 132 253 
rect 131 257 132 258 
rect 131 261 132 262 
rect 131 276 132 277 
rect 131 278 132 279 
rect 132 18 133 19 
rect 132 40 133 41 
rect 132 48 133 49 
rect 132 50 133 51 
rect 132 52 133 53 
rect 132 54 133 55 
rect 132 56 133 57 
rect 132 65 133 66 
rect 132 67 133 68 
rect 132 71 133 72 
rect 132 81 133 82 
rect 132 84 133 85 
rect 132 86 133 87 
rect 132 88 133 89 
rect 132 97 133 98 
rect 132 99 133 100 
rect 132 102 133 103 
rect 132 104 133 105 
rect 132 134 133 135 
rect 132 135 133 136 
rect 132 136 133 137 
rect 132 137 133 138 
rect 132 145 133 146 
rect 132 148 133 149 
rect 132 163 133 164 
rect 132 167 133 168 
rect 132 177 133 178 
rect 132 184 133 185 
rect 132 193 133 194 
rect 132 199 133 200 
rect 132 210 133 211 
rect 132 214 133 215 
rect 132 216 133 217 
rect 132 217 133 218 
rect 132 218 133 219 
rect 132 219 133 220 
rect 132 220 133 221 
rect 132 228 133 229 
rect 132 229 133 230 
rect 132 230 133 231 
rect 132 231 133 232 
rect 132 232 133 233 
rect 132 233 133 234 
rect 132 234 133 235 
rect 132 235 133 236 
rect 132 236 133 237 
rect 132 237 133 238 
rect 132 238 133 239 
rect 132 239 133 240 
rect 132 240 133 241 
rect 132 241 133 242 
rect 132 242 133 243 
rect 132 243 133 244 
rect 132 244 133 245 
rect 132 245 133 246 
rect 132 246 133 247 
rect 132 247 133 248 
rect 132 248 133 249 
rect 132 249 133 250 
rect 132 252 133 253 
rect 132 257 133 258 
rect 132 261 133 262 
rect 132 276 133 277 
rect 132 278 133 279 
rect 133 18 134 19 
rect 133 40 134 41 
rect 133 50 134 51 
rect 133 52 134 53 
rect 133 54 134 55 
rect 133 56 134 57 
rect 133 65 134 66 
rect 133 67 134 68 
rect 133 71 134 72 
rect 133 81 134 82 
rect 133 84 134 85 
rect 133 88 134 89 
rect 133 99 134 100 
rect 133 102 134 103 
rect 133 104 134 105 
rect 133 116 134 117 
rect 133 134 134 135 
rect 133 145 134 146 
rect 133 148 134 149 
rect 133 163 134 164 
rect 133 167 134 168 
rect 133 177 134 178 
rect 133 184 134 185 
rect 133 193 134 194 
rect 133 199 134 200 
rect 133 210 134 211 
rect 133 214 134 215 
rect 133 216 134 217 
rect 133 228 134 229 
rect 133 252 134 253 
rect 133 257 134 258 
rect 133 261 134 262 
rect 133 276 134 277 
rect 133 278 134 279 
rect 134 18 135 19 
rect 134 40 135 41 
rect 134 50 135 51 
rect 134 52 135 53 
rect 134 54 135 55 
rect 134 56 135 57 
rect 134 65 135 66 
rect 134 67 135 68 
rect 134 69 135 70 
rect 134 71 135 72 
rect 134 81 135 82 
rect 134 88 135 89 
rect 134 99 135 100 
rect 134 102 135 103 
rect 134 104 135 105 
rect 134 112 135 113 
rect 134 113 135 114 
rect 134 114 135 115 
rect 134 116 135 117 
rect 134 118 135 119 
rect 134 134 135 135 
rect 134 145 135 146 
rect 134 148 135 149 
rect 134 163 135 164 
rect 134 165 135 166 
rect 134 167 135 168 
rect 134 177 135 178 
rect 134 182 135 183 
rect 134 184 135 185 
rect 134 193 135 194 
rect 134 199 135 200 
rect 134 210 135 211 
rect 134 212 135 213 
rect 134 214 135 215 
rect 134 216 135 217 
rect 134 228 135 229 
rect 134 230 135 231 
rect 134 242 135 243 
rect 134 243 135 244 
rect 134 257 135 258 
rect 134 261 135 262 
rect 134 276 135 277 
rect 134 278 135 279 
rect 135 18 136 19 
rect 135 40 136 41 
rect 135 50 136 51 
rect 135 52 136 53 
rect 135 54 136 55 
rect 135 56 136 57 
rect 135 65 136 66 
rect 135 67 136 68 
rect 135 69 136 70 
rect 135 71 136 72 
rect 135 81 136 82 
rect 135 88 136 89 
rect 135 97 136 98 
rect 135 99 136 100 
rect 135 102 136 103 
rect 135 104 136 105 
rect 135 114 136 115 
rect 135 116 136 117 
rect 135 118 136 119 
rect 135 132 136 133 
rect 135 134 136 135 
rect 135 136 136 137 
rect 135 145 136 146 
rect 135 148 136 149 
rect 135 152 136 153 
rect 135 161 136 162 
rect 135 163 136 164 
rect 135 165 136 166 
rect 135 167 136 168 
rect 135 177 136 178 
rect 135 182 136 183 
rect 135 184 136 185 
rect 135 193 136 194 
rect 135 195 136 196 
rect 135 199 136 200 
rect 135 210 136 211 
rect 135 212 136 213 
rect 135 214 136 215 
rect 135 216 136 217 
rect 135 228 136 229 
rect 135 230 136 231 
rect 135 232 136 233 
rect 135 243 136 244 
rect 135 246 136 247 
rect 135 248 136 249 
rect 135 257 136 258 
rect 135 259 136 260 
rect 135 261 136 262 
rect 135 276 136 277 
rect 135 278 136 279 
rect 135 280 136 281 
rect 136 18 137 19 
rect 136 40 137 41 
rect 136 50 137 51 
rect 136 52 137 53 
rect 136 54 137 55 
rect 136 56 137 57 
rect 136 65 137 66 
rect 136 67 137 68 
rect 136 69 137 70 
rect 136 71 137 72 
rect 136 81 137 82 
rect 136 88 137 89 
rect 136 97 137 98 
rect 136 99 137 100 
rect 136 102 137 103 
rect 136 104 137 105 
rect 136 114 137 115 
rect 136 116 137 117 
rect 136 118 137 119 
rect 136 132 137 133 
rect 136 134 137 135 
rect 136 136 137 137 
rect 136 145 137 146 
rect 136 148 137 149 
rect 136 152 137 153 
rect 136 161 137 162 
rect 136 163 137 164 
rect 136 165 137 166 
rect 136 167 137 168 
rect 136 177 137 178 
rect 136 182 137 183 
rect 136 184 137 185 
rect 136 193 137 194 
rect 136 195 137 196 
rect 136 199 137 200 
rect 136 210 137 211 
rect 136 212 137 213 
rect 136 214 137 215 
rect 136 216 137 217 
rect 136 228 137 229 
rect 136 230 137 231 
rect 136 232 137 233 
rect 136 243 137 244 
rect 136 246 137 247 
rect 136 248 137 249 
rect 136 257 137 258 
rect 136 259 137 260 
rect 136 261 137 262 
rect 136 276 137 277 
rect 136 278 137 279 
rect 136 280 137 281 
rect 136 289 137 290 
rect 137 18 138 19 
rect 137 40 138 41 
rect 137 50 138 51 
rect 137 52 138 53 
rect 137 54 138 55 
rect 137 56 138 57 
rect 137 65 138 66 
rect 137 67 138 68 
rect 137 69 138 70 
rect 137 71 138 72 
rect 137 81 138 82 
rect 137 88 138 89 
rect 137 97 138 98 
rect 137 99 138 100 
rect 137 102 138 103 
rect 137 104 138 105 
rect 137 114 138 115 
rect 137 116 138 117 
rect 137 118 138 119 
rect 137 132 138 133 
rect 137 134 138 135 
rect 137 136 138 137 
rect 137 145 138 146 
rect 137 148 138 149 
rect 137 152 138 153 
rect 137 161 138 162 
rect 137 163 138 164 
rect 137 165 138 166 
rect 137 167 138 168 
rect 137 177 138 178 
rect 137 182 138 183 
rect 137 184 138 185 
rect 137 193 138 194 
rect 137 195 138 196 
rect 137 199 138 200 
rect 137 210 138 211 
rect 137 212 138 213 
rect 137 214 138 215 
rect 137 216 138 217 
rect 137 228 138 229 
rect 137 230 138 231 
rect 137 232 138 233 
rect 137 243 138 244 
rect 137 246 138 247 
rect 137 248 138 249 
rect 137 257 138 258 
rect 137 259 138 260 
rect 137 261 138 262 
rect 137 276 138 277 
rect 137 278 138 279 
rect 137 280 138 281 
rect 137 289 138 290 
rect 137 291 138 292 
rect 138 18 139 19 
rect 138 40 139 41 
rect 138 50 139 51 
rect 138 52 139 53 
rect 138 54 139 55 
rect 138 56 139 57 
rect 138 65 139 66 
rect 138 67 139 68 
rect 138 69 139 70 
rect 138 71 139 72 
rect 138 81 139 82 
rect 138 88 139 89 
rect 138 97 139 98 
rect 138 99 139 100 
rect 138 102 139 103 
rect 138 104 139 105 
rect 138 114 139 115 
rect 138 116 139 117 
rect 138 132 139 133 
rect 138 134 139 135 
rect 138 136 139 137 
rect 138 145 139 146 
rect 138 148 139 149 
rect 138 152 139 153 
rect 138 161 139 162 
rect 138 163 139 164 
rect 138 165 139 166 
rect 138 167 139 168 
rect 138 177 139 178 
rect 138 182 139 183 
rect 138 184 139 185 
rect 138 193 139 194 
rect 138 195 139 196 
rect 138 199 139 200 
rect 138 210 139 211 
rect 138 212 139 213 
rect 138 214 139 215 
rect 138 216 139 217 
rect 138 228 139 229 
rect 138 230 139 231 
rect 138 232 139 233 
rect 138 243 139 244 
rect 138 246 139 247 
rect 138 248 139 249 
rect 138 257 139 258 
rect 138 259 139 260 
rect 138 261 139 262 
rect 138 276 139 277 
rect 138 278 139 279 
rect 138 280 139 281 
rect 138 289 139 290 
rect 138 291 139 292 
rect 139 18 140 19 
rect 139 40 140 41 
rect 139 50 140 51 
rect 139 52 140 53 
rect 139 54 140 55 
rect 139 56 140 57 
rect 139 65 140 66 
rect 139 67 140 68 
rect 139 69 140 70 
rect 139 71 140 72 
rect 139 81 140 82 
rect 139 88 140 89 
rect 139 97 140 98 
rect 139 99 140 100 
rect 139 102 140 103 
rect 139 104 140 105 
rect 139 114 140 115 
rect 139 115 140 116 
rect 139 132 140 133 
rect 139 152 140 153 
rect 139 163 140 164 
rect 139 165 140 166 
rect 139 167 140 168 
rect 139 177 140 178 
rect 139 182 140 183 
rect 139 184 140 185 
rect 139 193 140 194 
rect 139 195 140 196 
rect 139 199 140 200 
rect 139 210 140 211 
rect 139 212 140 213 
rect 139 214 140 215 
rect 139 216 140 217 
rect 139 228 140 229 
rect 139 230 140 231 
rect 139 243 140 244 
rect 139 246 140 247 
rect 139 257 140 258 
rect 139 261 140 262 
rect 139 276 140 277 
rect 139 278 140 279 
rect 139 289 140 290 
rect 139 291 140 292 
rect 140 18 141 19 
rect 140 40 141 41 
rect 140 50 141 51 
rect 140 52 141 53 
rect 140 54 141 55 
rect 140 56 141 57 
rect 140 65 141 66 
rect 140 67 141 68 
rect 140 69 141 70 
rect 140 71 141 72 
rect 140 81 141 82 
rect 140 88 141 89 
rect 140 97 141 98 
rect 140 99 141 100 
rect 140 102 141 103 
rect 140 104 141 105 
rect 140 115 141 116 
rect 140 116 141 117 
rect 140 117 141 118 
rect 140 118 141 119 
rect 140 119 141 120 
rect 140 132 141 133 
rect 140 152 141 153 
rect 140 163 141 164 
rect 140 165 141 166 
rect 140 167 141 168 
rect 140 177 141 178 
rect 140 182 141 183 
rect 140 184 141 185 
rect 140 193 141 194 
rect 140 195 141 196 
rect 140 199 141 200 
rect 140 210 141 211 
rect 140 212 141 213 
rect 140 214 141 215 
rect 140 216 141 217 
rect 140 228 141 229 
rect 140 243 141 244 
rect 140 246 141 247 
rect 140 257 141 258 
rect 140 261 141 262 
rect 140 276 141 277 
rect 140 278 141 279 
rect 140 289 141 290 
rect 140 291 141 292 
rect 141 18 142 19 
rect 141 40 142 41 
rect 141 50 142 51 
rect 141 52 142 53 
rect 141 54 142 55 
rect 141 56 142 57 
rect 141 65 142 66 
rect 141 67 142 68 
rect 141 69 142 70 
rect 141 71 142 72 
rect 141 81 142 82 
rect 141 88 142 89 
rect 141 97 142 98 
rect 141 99 142 100 
rect 141 102 142 103 
rect 141 104 142 105 
rect 141 119 142 120 
rect 141 132 142 133 
rect 141 152 142 153 
rect 141 165 142 166 
rect 141 167 142 168 
rect 141 177 142 178 
rect 141 182 142 183 
rect 141 184 142 185 
rect 141 193 142 194 
rect 141 195 142 196 
rect 141 199 142 200 
rect 141 210 142 211 
rect 141 212 142 213 
rect 141 214 142 215 
rect 141 216 142 217 
rect 141 246 142 247 
rect 141 257 142 258 
rect 141 261 142 262 
rect 141 276 142 277 
rect 141 277 142 278 
rect 142 18 143 19 
rect 142 40 143 41 
rect 142 50 143 51 
rect 142 52 143 53 
rect 142 54 143 55 
rect 142 56 143 57 
rect 142 65 143 66 
rect 142 67 143 68 
rect 142 69 143 70 
rect 142 71 143 72 
rect 142 81 143 82 
rect 142 88 143 89 
rect 142 97 143 98 
rect 142 99 143 100 
rect 142 102 143 103 
rect 142 104 143 105 
rect 142 119 143 120 
rect 142 132 143 133 
rect 142 152 143 153 
rect 142 162 143 163 
rect 142 163 143 164 
rect 142 164 143 165 
rect 142 165 143 166 
rect 142 167 143 168 
rect 142 177 143 178 
rect 142 182 143 183 
rect 142 184 143 185 
rect 142 193 143 194 
rect 142 195 143 196 
rect 142 199 143 200 
rect 142 210 143 211 
rect 142 212 143 213 
rect 142 214 143 215 
rect 142 216 143 217 
rect 142 246 143 247 
rect 142 257 143 258 
rect 142 261 143 262 
rect 142 277 143 278 
rect 142 278 143 279 
rect 143 18 144 19 
rect 143 40 144 41 
rect 143 50 144 51 
rect 143 52 144 53 
rect 143 54 144 55 
rect 143 56 144 57 
rect 143 65 144 66 
rect 143 67 144 68 
rect 143 69 144 70 
rect 143 71 144 72 
rect 143 81 144 82 
rect 143 88 144 89 
rect 143 97 144 98 
rect 143 99 144 100 
rect 143 102 144 103 
rect 143 104 144 105 
rect 143 119 144 120 
rect 143 132 144 133 
rect 143 152 144 153 
rect 143 167 144 168 
rect 143 177 144 178 
rect 143 182 144 183 
rect 143 184 144 185 
rect 143 193 144 194 
rect 143 195 144 196 
rect 143 199 144 200 
rect 143 210 144 211 
rect 143 212 144 213 
rect 143 214 144 215 
rect 143 216 144 217 
rect 143 246 144 247 
rect 143 257 144 258 
rect 143 261 144 262 
rect 144 18 145 19 
rect 144 40 145 41 
rect 144 50 145 51 
rect 144 52 145 53 
rect 144 54 145 55 
rect 144 56 145 57 
rect 144 65 145 66 
rect 144 67 145 68 
rect 144 69 145 70 
rect 144 71 145 72 
rect 144 81 145 82 
rect 144 88 145 89 
rect 144 97 145 98 
rect 144 99 145 100 
rect 144 102 145 103 
rect 144 104 145 105 
rect 144 119 145 120 
rect 144 132 145 133 
rect 144 152 145 153 
rect 144 153 145 154 
rect 144 176 145 177 
rect 144 177 145 178 
rect 144 182 145 183 
rect 144 184 145 185 
rect 144 193 145 194 
rect 144 195 145 196 
rect 144 199 145 200 
rect 144 210 145 211 
rect 144 212 145 213 
rect 144 214 145 215 
rect 144 216 145 217 
rect 144 246 145 247 
rect 144 257 145 258 
rect 144 261 145 262 
rect 145 18 146 19 
rect 145 40 146 41 
rect 145 50 146 51 
rect 145 52 146 53 
rect 145 54 146 55 
rect 145 56 146 57 
rect 145 65 146 66 
rect 145 67 146 68 
rect 145 69 146 70 
rect 145 71 146 72 
rect 145 81 146 82 
rect 145 88 146 89 
rect 145 97 146 98 
rect 145 99 146 100 
rect 145 102 146 103 
rect 145 104 146 105 
rect 145 119 146 120 
rect 145 120 146 121 
rect 145 121 146 122 
rect 145 122 146 123 
rect 145 123 146 124 
rect 145 124 146 125 
rect 145 125 146 126 
rect 145 126 146 127 
rect 145 127 146 128 
rect 145 128 146 129 
rect 145 129 146 130 
rect 145 130 146 131 
rect 145 132 146 133 
rect 145 153 146 154 
rect 145 154 146 155 
rect 145 155 146 156 
rect 145 156 146 157 
rect 145 157 146 158 
rect 145 158 146 159 
rect 145 159 146 160 
rect 145 160 146 161 
rect 145 161 146 162 
rect 145 162 146 163 
rect 145 163 146 164 
rect 145 164 146 165 
rect 145 165 146 166 
rect 145 166 146 167 
rect 145 167 146 168 
rect 145 168 146 169 
rect 145 169 146 170 
rect 145 170 146 171 
rect 145 171 146 172 
rect 145 173 146 174 
rect 145 174 146 175 
rect 145 175 146 176 
rect 145 176 146 177 
rect 145 182 146 183 
rect 145 184 146 185 
rect 145 193 146 194 
rect 145 195 146 196 
rect 145 199 146 200 
rect 145 210 146 211 
rect 145 212 146 213 
rect 145 214 146 215 
rect 145 216 146 217 
rect 145 223 146 224 
rect 145 224 146 225 
rect 145 225 146 226 
rect 145 226 146 227 
rect 145 227 146 228 
rect 145 228 146 229 
rect 145 229 146 230 
rect 145 230 146 231 
rect 145 231 146 232 
rect 145 232 146 233 
rect 145 233 146 234 
rect 145 234 146 235 
rect 145 235 146 236 
rect 145 236 146 237 
rect 145 237 146 238 
rect 145 238 146 239 
rect 145 239 146 240 
rect 145 240 146 241 
rect 145 241 146 242 
rect 145 242 146 243 
rect 145 246 146 247 
rect 145 257 146 258 
rect 145 261 146 262 
rect 145 287 146 288 
rect 145 288 146 289 
rect 145 289 146 290 
rect 145 290 146 291 
rect 145 291 146 292 
rect 145 292 146 293 
rect 145 293 146 294 
rect 145 294 146 295 
rect 145 295 146 296 
rect 146 40 147 41 
rect 146 50 147 51 
rect 146 52 147 53 
rect 146 54 147 55 
rect 146 56 147 57 
rect 146 65 147 66 
rect 146 67 147 68 
rect 146 69 147 70 
rect 146 71 147 72 
rect 146 81 147 82 
rect 146 88 147 89 
rect 146 97 147 98 
rect 146 99 147 100 
rect 146 102 147 103 
rect 146 104 147 105 
rect 146 130 147 131 
rect 146 132 147 133 
rect 146 172 147 173 
rect 146 173 147 174 
rect 146 182 147 183 
rect 146 184 147 185 
rect 146 193 147 194 
rect 146 195 147 196 
rect 146 199 147 200 
rect 146 210 147 211 
rect 146 212 147 213 
rect 146 214 147 215 
rect 146 216 147 217 
rect 146 246 147 247 
rect 146 257 147 258 
rect 146 261 147 262 
rect 147 40 148 41 
rect 147 50 148 51 
rect 147 52 148 53 
rect 147 54 148 55 
rect 147 56 148 57 
rect 147 65 148 66 
rect 147 67 148 68 
rect 147 69 148 70 
rect 147 71 148 72 
rect 147 81 148 82 
rect 147 88 148 89 
rect 147 97 148 98 
rect 147 99 148 100 
rect 147 102 148 103 
rect 147 104 148 105 
rect 147 130 148 131 
rect 147 132 148 133 
rect 147 158 148 159 
rect 147 159 148 160 
rect 147 160 148 161 
rect 147 161 148 162 
rect 147 162 148 163 
rect 147 163 148 164 
rect 147 164 148 165 
rect 147 165 148 166 
rect 147 167 148 168 
rect 147 168 148 169 
rect 147 169 148 170 
rect 147 170 148 171 
rect 147 171 148 172 
rect 147 172 148 173 
rect 147 182 148 183 
rect 147 193 148 194 
rect 147 195 148 196 
rect 147 199 148 200 
rect 147 212 148 213 
rect 147 214 148 215 
rect 147 216 148 217 
rect 147 238 148 239 
rect 147 239 148 240 
rect 147 240 148 241 
rect 147 241 148 242 
rect 147 242 148 243 
rect 147 243 148 244 
rect 147 246 148 247 
rect 147 248 148 249 
rect 147 257 148 258 
rect 147 259 148 260 
rect 147 261 148 262 
rect 147 263 148 264 
rect 148 40 149 41 
rect 148 50 149 51 
rect 148 52 149 53 
rect 148 54 149 55 
rect 148 65 149 66 
rect 148 67 149 68 
rect 148 69 149 70 
rect 148 71 149 72 
rect 148 81 149 82 
rect 148 88 149 89 
rect 148 97 149 98 
rect 148 99 149 100 
rect 148 102 149 103 
rect 148 130 149 131 
rect 148 132 149 133 
rect 148 182 149 183 
rect 148 183 149 184 
rect 148 184 149 185 
rect 148 185 149 186 
rect 148 186 149 187 
rect 148 187 149 188 
rect 148 188 149 189 
rect 148 189 149 190 
rect 148 193 149 194 
rect 148 195 149 196 
rect 148 199 149 200 
rect 148 211 149 212 
rect 148 212 149 213 
rect 148 214 149 215 
rect 148 216 149 217 
rect 148 246 149 247 
rect 148 248 149 249 
rect 148 257 149 258 
rect 148 259 149 260 
rect 148 261 149 262 
rect 148 263 149 264 
rect 149 40 150 41 
rect 149 50 150 51 
rect 149 52 150 53 
rect 149 54 150 55 
rect 149 57 150 58 
rect 149 65 150 66 
rect 149 67 150 68 
rect 149 69 150 70 
rect 149 71 150 72 
rect 149 81 150 82 
rect 149 88 150 89 
rect 149 97 150 98 
rect 149 99 150 100 
rect 149 102 150 103 
rect 149 130 150 131 
rect 149 132 150 133 
rect 149 157 150 158 
rect 149 158 150 159 
rect 149 159 150 160 
rect 149 160 150 161 
rect 149 161 150 162 
rect 149 162 150 163 
rect 149 163 150 164 
rect 149 164 150 165 
rect 149 165 150 166 
rect 149 166 150 167 
rect 149 167 150 168 
rect 149 168 150 169 
rect 149 169 150 170 
rect 149 170 150 171 
rect 149 189 150 190 
rect 149 193 150 194 
rect 149 195 150 196 
rect 149 199 150 200 
rect 149 210 150 211 
rect 149 211 150 212 
rect 149 214 150 215 
rect 149 216 150 217 
rect 149 246 150 247 
rect 149 248 150 249 
rect 149 257 150 258 
rect 149 259 150 260 
rect 149 261 150 262 
rect 149 263 150 264 
rect 150 40 151 41 
rect 150 50 151 51 
rect 150 52 151 53 
rect 150 54 151 55 
rect 150 57 151 58 
rect 150 65 151 66 
rect 150 67 151 68 
rect 150 69 151 70 
rect 150 71 151 72 
rect 150 81 151 82 
rect 150 88 151 89 
rect 150 97 151 98 
rect 150 99 151 100 
rect 150 102 151 103 
rect 150 130 151 131 
rect 150 132 151 133 
rect 150 193 151 194 
rect 150 195 151 196 
rect 150 197 151 198 
rect 150 199 151 200 
rect 150 210 151 211 
rect 150 214 151 215 
rect 150 216 151 217 
rect 150 246 151 247 
rect 150 248 151 249 
rect 150 257 151 258 
rect 150 259 151 260 
rect 150 261 151 262 
rect 150 263 151 264 
rect 150 269 151 270 
rect 150 270 151 271 
rect 150 271 151 272 
rect 150 272 151 273 
rect 150 273 151 274 
rect 151 40 152 41 
rect 151 50 152 51 
rect 151 52 152 53 
rect 151 54 152 55 
rect 151 57 152 58 
rect 151 65 152 66 
rect 151 67 152 68 
rect 151 69 152 70 
rect 151 71 152 72 
rect 151 81 152 82 
rect 151 88 152 89 
rect 151 97 152 98 
rect 151 99 152 100 
rect 151 102 152 103 
rect 151 130 152 131 
rect 151 132 152 133 
rect 151 193 152 194 
rect 151 195 152 196 
rect 151 197 152 198 
rect 151 199 152 200 
rect 151 210 152 211 
rect 151 214 152 215 
rect 151 216 152 217 
rect 151 246 152 247 
rect 151 248 152 249 
rect 151 257 152 258 
rect 151 259 152 260 
rect 151 261 152 262 
rect 151 263 152 264 
rect 151 269 152 270 
rect 151 273 152 274 
rect 151 274 152 275 
rect 152 40 153 41 
rect 152 50 153 51 
rect 152 52 153 53 
rect 152 54 153 55 
rect 152 56 153 57 
rect 152 57 153 58 
rect 152 65 153 66 
rect 152 67 153 68 
rect 152 69 153 70 
rect 152 71 153 72 
rect 152 81 153 82 
rect 152 88 153 89 
rect 152 97 153 98 
rect 152 99 153 100 
rect 152 102 153 103 
rect 152 130 153 131 
rect 152 132 153 133 
rect 152 137 153 138 
rect 152 138 153 139 
rect 152 139 153 140 
rect 152 140 153 141 
rect 152 141 153 142 
rect 152 142 153 143 
rect 152 143 153 144 
rect 152 144 153 145 
rect 152 145 153 146 
rect 152 146 153 147 
rect 152 147 153 148 
rect 152 148 153 149 
rect 152 149 153 150 
rect 152 150 153 151 
rect 152 151 153 152 
rect 152 152 153 153 
rect 152 153 153 154 
rect 152 154 153 155 
rect 152 155 153 156 
rect 152 156 153 157 
rect 152 157 153 158 
rect 152 158 153 159 
rect 152 159 153 160 
rect 152 160 153 161 
rect 152 161 153 162 
rect 152 162 153 163 
rect 152 163 153 164 
rect 152 164 153 165 
rect 152 165 153 166 
rect 152 166 153 167 
rect 152 167 153 168 
rect 152 168 153 169 
rect 152 169 153 170 
rect 152 170 153 171 
rect 152 171 153 172 
rect 152 172 153 173 
rect 152 173 153 174 
rect 152 174 153 175 
rect 152 175 153 176 
rect 152 176 153 177 
rect 152 177 153 178 
rect 152 178 153 179 
rect 152 179 153 180 
rect 152 180 153 181 
rect 152 181 153 182 
rect 152 182 153 183 
rect 152 183 153 184 
rect 152 184 153 185 
rect 152 185 153 186 
rect 152 186 153 187 
rect 152 193 153 194 
rect 152 195 153 196 
rect 152 197 153 198 
rect 152 199 153 200 
rect 152 210 153 211 
rect 152 214 153 215 
rect 152 216 153 217 
rect 152 246 153 247 
rect 152 248 153 249 
rect 152 257 153 258 
rect 152 259 153 260 
rect 152 261 153 262 
rect 152 263 153 264 
rect 152 269 153 270 
rect 152 271 153 272 
rect 152 272 153 273 
rect 152 274 153 275 
rect 152 275 153 276 
rect 152 276 153 277 
rect 152 277 153 278 
rect 152 278 153 279 
rect 152 279 153 280 
rect 152 280 153 281 
rect 152 281 153 282 
rect 152 282 153 283 
rect 152 283 153 284 
rect 152 284 153 285 
rect 152 285 153 286 
rect 152 286 153 287 
rect 152 287 153 288 
rect 152 288 153 289 
rect 153 24 154 25 
rect 153 40 154 41 
rect 153 50 154 51 
rect 153 52 154 53 
rect 153 54 154 55 
rect 153 56 154 57 
rect 153 65 154 66 
rect 153 67 154 68 
rect 153 69 154 70 
rect 153 71 154 72 
rect 153 81 154 82 
rect 153 88 154 89 
rect 153 97 154 98 
rect 153 99 154 100 
rect 153 102 154 103 
rect 153 130 154 131 
rect 153 132 154 133 
rect 153 135 154 136 
rect 153 136 154 137 
rect 153 137 154 138 
rect 153 193 154 194 
rect 153 195 154 196 
rect 153 197 154 198 
rect 153 199 154 200 
rect 153 210 154 211 
rect 153 214 154 215 
rect 153 216 154 217 
rect 153 246 154 247 
rect 153 248 154 249 
rect 153 257 154 258 
rect 153 259 154 260 
rect 153 261 154 262 
rect 153 263 154 264 
rect 153 272 154 273 
rect 153 273 154 274 
rect 153 288 154 289 
rect 153 289 154 290 
rect 154 24 155 25 
rect 154 40 155 41 
rect 154 50 155 51 
rect 154 52 155 53 
rect 154 54 155 55 
rect 154 56 155 57 
rect 154 65 155 66 
rect 154 67 155 68 
rect 154 81 155 82 
rect 154 88 155 89 
rect 154 97 155 98 
rect 154 99 155 100 
rect 154 102 155 103 
rect 154 130 155 131 
rect 154 132 155 133 
rect 154 193 155 194 
rect 154 195 155 196 
rect 154 197 155 198 
rect 154 199 155 200 
rect 154 210 155 211 
rect 154 214 155 215 
rect 154 216 155 217 
rect 154 246 155 247 
rect 154 248 155 249 
rect 154 257 155 258 
rect 154 259 155 260 
rect 154 261 155 262 
rect 154 263 155 264 
rect 154 273 155 274 
rect 154 274 155 275 
rect 154 275 155 276 
rect 154 276 155 277 
rect 154 277 155 278 
rect 154 278 155 279 
rect 154 279 155 280 
rect 154 289 155 290 
rect 155 24 156 25 
rect 155 40 156 41 
rect 155 50 156 51 
rect 155 51 156 52 
rect 155 54 156 55 
rect 155 56 156 57 
rect 155 67 156 68 
rect 155 81 156 82 
rect 155 88 156 89 
rect 155 99 156 100 
rect 155 102 156 103 
rect 155 130 156 131 
rect 155 131 156 132 
rect 155 193 156 194 
rect 155 195 156 196 
rect 155 197 156 198 
rect 155 199 156 200 
rect 155 210 156 211 
rect 155 214 156 215 
rect 155 257 156 258 
rect 155 260 156 261 
rect 155 261 156 262 
rect 155 263 156 264 
rect 155 289 156 290 
rect 156 24 157 25 
rect 156 40 157 41 
rect 156 51 157 52 
rect 156 52 157 53 
rect 156 54 157 55 
rect 156 56 157 57 
rect 156 67 157 68 
rect 156 81 157 82 
rect 156 88 157 89 
rect 156 99 157 100 
rect 156 102 157 103 
rect 156 131 157 132 
rect 156 132 157 133 
rect 156 133 157 134 
rect 156 134 157 135 
rect 156 135 157 136 
rect 156 136 157 137 
rect 156 193 157 194 
rect 156 195 157 196 
rect 156 197 157 198 
rect 156 199 157 200 
rect 156 210 157 211 
rect 156 214 157 215 
rect 156 257 157 258 
rect 156 259 157 260 
rect 156 260 157 261 
rect 156 263 157 264 
rect 156 289 157 290 
rect 157 24 158 25 
rect 157 40 158 41 
rect 157 53 158 54 
rect 157 54 158 55 
rect 157 56 158 57 
rect 157 67 158 68 
rect 157 81 158 82 
rect 157 88 158 89 
rect 157 99 158 100 
rect 157 102 158 103 
rect 157 136 158 137 
rect 157 193 158 194 
rect 157 195 158 196 
rect 157 197 158 198 
rect 157 199 158 200 
rect 157 210 158 211 
rect 157 214 158 215 
rect 157 257 158 258 
rect 157 259 158 260 
rect 157 263 158 264 
rect 157 289 158 290 
rect 158 24 159 25 
rect 158 40 159 41 
rect 158 49 159 50 
rect 158 50 159 51 
rect 158 51 159 52 
rect 158 52 159 53 
rect 158 53 159 54 
rect 158 55 159 56 
rect 158 56 159 57 
rect 158 67 159 68 
rect 158 81 159 82 
rect 158 88 159 89 
rect 158 99 159 100 
rect 158 102 159 103 
rect 158 136 159 137 
rect 158 193 159 194 
rect 158 195 159 196 
rect 158 197 159 198 
rect 158 199 159 200 
rect 158 210 159 211 
rect 158 214 159 215 
rect 158 257 159 258 
rect 158 259 159 260 
rect 158 263 159 264 
rect 158 289 159 290 
rect 159 24 160 25 
rect 159 40 160 41 
rect 159 49 160 50 
rect 159 54 160 55 
rect 159 55 160 56 
rect 159 67 160 68 
rect 159 81 160 82 
rect 159 88 160 89 
rect 159 99 160 100 
rect 159 102 160 103 
rect 159 104 160 105 
rect 159 136 160 137 
rect 159 193 160 194 
rect 159 195 160 196 
rect 159 197 160 198 
rect 159 199 160 200 
rect 159 210 160 211 
rect 159 214 160 215 
rect 159 257 160 258 
rect 159 259 160 260 
rect 159 263 160 264 
rect 159 289 160 290 
rect 160 24 161 25 
rect 160 40 161 41 
rect 160 48 161 49 
rect 160 49 161 50 
rect 160 51 161 52 
rect 160 52 161 53 
rect 160 53 161 54 
rect 160 54 161 55 
rect 160 67 161 68 
rect 160 81 161 82 
rect 160 88 161 89 
rect 160 99 161 100 
rect 160 102 161 103 
rect 160 104 161 105 
rect 160 105 161 106 
rect 160 136 161 137 
rect 160 137 161 138 
rect 160 193 161 194 
rect 160 195 161 196 
rect 160 197 161 198 
rect 160 199 161 200 
rect 160 210 161 211 
rect 160 214 161 215 
rect 160 256 161 257 
rect 160 257 161 258 
rect 160 259 161 260 
rect 160 263 161 264 
rect 160 289 161 290 
rect 161 18 162 19 
rect 161 19 162 20 
rect 161 20 162 21 
rect 161 21 162 22 
rect 161 22 162 23 
rect 161 23 162 24 
rect 161 24 162 25 
rect 161 40 162 41 
rect 161 50 162 51 
rect 161 51 162 52 
rect 161 67 162 68 
rect 161 81 162 82 
rect 161 88 162 89 
rect 161 99 162 100 
rect 161 102 162 103 
rect 161 105 162 106 
rect 161 106 162 107 
rect 161 107 162 108 
rect 161 108 162 109 
rect 161 109 162 110 
rect 161 110 162 111 
rect 161 111 162 112 
rect 161 112 162 113 
rect 161 113 162 114 
rect 161 114 162 115 
rect 161 116 162 117 
rect 161 117 162 118 
rect 161 118 162 119 
rect 161 119 162 120 
rect 161 137 162 138 
rect 161 138 162 139 
rect 161 165 162 166 
rect 161 193 162 194 
rect 161 195 162 196 
rect 161 197 162 198 
rect 161 199 162 200 
rect 161 210 162 211 
rect 161 214 162 215 
rect 161 246 162 247 
rect 161 247 162 248 
rect 161 248 162 249 
rect 161 249 162 250 
rect 161 250 162 251 
rect 161 251 162 252 
rect 161 252 162 253 
rect 161 253 162 254 
rect 161 254 162 255 
rect 161 255 162 256 
rect 161 256 162 257 
rect 161 259 162 260 
rect 161 263 162 264 
rect 161 289 162 290 
rect 162 40 163 41 
rect 162 49 163 50 
rect 162 50 163 51 
rect 162 67 163 68 
rect 162 81 163 82 
rect 162 88 163 89 
rect 162 94 163 95 
rect 162 95 163 96 
rect 162 96 163 97 
rect 162 97 163 98 
rect 162 98 163 99 
rect 162 99 163 100 
rect 162 102 163 103 
rect 162 114 163 115 
rect 162 115 163 116 
rect 162 165 163 166 
rect 162 193 163 194 
rect 162 195 163 196 
rect 162 197 163 198 
rect 162 199 163 200 
rect 162 201 163 202 
rect 162 210 163 211 
rect 162 214 163 215 
rect 162 259 163 260 
rect 162 263 163 264 
rect 162 289 163 290 
rect 163 16 164 17 
rect 163 17 164 18 
rect 163 18 164 19 
rect 163 19 164 20 
rect 163 20 164 21 
rect 163 21 164 22 
rect 163 22 164 23 
rect 163 23 164 24 
rect 163 24 164 25 
rect 163 40 164 41 
rect 163 49 164 50 
rect 163 67 164 68 
rect 163 81 164 82 
rect 163 88 164 89 
rect 163 94 164 95 
rect 163 102 164 103 
rect 163 115 164 116 
rect 163 116 164 117 
rect 163 117 164 118 
rect 163 118 164 119 
rect 163 119 164 120 
rect 163 120 164 121 
rect 163 121 164 122 
rect 163 122 164 123 
rect 163 123 164 124 
rect 163 124 164 125 
rect 163 125 164 126 
rect 163 126 164 127 
rect 163 127 164 128 
rect 163 128 164 129 
rect 163 129 164 130 
rect 163 130 164 131 
rect 163 131 164 132 
rect 163 132 164 133 
rect 163 133 164 134 
rect 163 134 164 135 
rect 163 135 164 136 
rect 163 136 164 137 
rect 163 137 164 138 
rect 163 138 164 139 
rect 163 165 164 166 
rect 163 193 164 194 
rect 163 195 164 196 
rect 163 197 164 198 
rect 163 199 164 200 
rect 163 201 164 202 
rect 163 210 164 211 
rect 163 214 164 215 
rect 163 230 164 231 
rect 163 231 164 232 
rect 163 232 164 233 
rect 163 233 164 234 
rect 163 234 164 235 
rect 163 235 164 236 
rect 163 236 164 237 
rect 163 237 164 238 
rect 163 238 164 239 
rect 163 239 164 240 
rect 163 240 164 241 
rect 163 241 164 242 
rect 163 242 164 243 
rect 163 243 164 244 
rect 163 244 164 245 
rect 163 245 164 246 
rect 163 246 164 247 
rect 163 247 164 248 
rect 163 248 164 249 
rect 163 249 164 250 
rect 163 250 164 251 
rect 163 259 164 260 
rect 163 263 164 264 
rect 163 289 164 290 
rect 164 40 165 41 
rect 164 49 165 50 
rect 164 67 165 68 
rect 164 81 165 82 
rect 164 88 165 89 
rect 164 95 165 96 
rect 164 96 165 97 
rect 164 97 165 98 
rect 164 98 165 99 
rect 164 102 165 103 
rect 164 165 165 166 
rect 164 193 165 194 
rect 164 195 165 196 
rect 164 197 165 198 
rect 164 199 165 200 
rect 164 201 165 202 
rect 164 210 165 211 
rect 164 214 165 215 
rect 164 263 165 264 
rect 164 289 165 290 
rect 165 40 166 41 
rect 165 49 166 50 
rect 165 67 166 68 
rect 165 81 166 82 
rect 165 88 166 89 
rect 165 102 166 103 
rect 165 116 166 117 
rect 165 117 166 118 
rect 165 118 166 119 
rect 165 119 166 120 
rect 165 120 166 121 
rect 165 121 166 122 
rect 165 122 166 123 
rect 165 123 166 124 
rect 165 124 166 125 
rect 165 125 166 126 
rect 165 126 166 127 
rect 165 127 166 128 
rect 165 128 166 129 
rect 165 129 166 130 
rect 165 130 166 131 
rect 165 131 166 132 
rect 165 132 166 133 
rect 165 133 166 134 
rect 165 134 166 135 
rect 165 135 166 136 
rect 165 136 166 137 
rect 165 137 166 138 
rect 165 138 166 139 
rect 165 139 166 140 
rect 165 140 166 141 
rect 165 141 166 142 
rect 165 142 166 143 
rect 165 143 166 144 
rect 165 144 166 145 
rect 165 145 166 146 
rect 165 146 166 147 
rect 165 147 166 148 
rect 165 148 166 149 
rect 165 149 166 150 
rect 165 150 166 151 
rect 165 151 166 152 
rect 165 152 166 153 
rect 165 153 166 154 
rect 165 193 166 194 
rect 165 195 166 196 
rect 165 199 166 200 
rect 165 201 166 202 
rect 165 210 166 211 
rect 165 214 166 215 
rect 165 263 166 264 
rect 165 271 166 272 
rect 165 272 166 273 
rect 165 273 166 274 
rect 165 274 166 275 
rect 165 275 166 276 
rect 165 276 166 277 
rect 165 277 166 278 
rect 165 278 166 279 
rect 165 279 166 280 
rect 165 280 166 281 
rect 165 281 166 282 
rect 165 282 166 283 
rect 165 289 166 290 
rect 166 40 167 41 
rect 166 49 167 50 
rect 166 67 167 68 
rect 166 81 167 82 
rect 166 88 167 89 
rect 166 102 167 103 
rect 166 163 167 164 
rect 166 164 167 165 
rect 166 165 167 166 
rect 166 166 167 167 
rect 166 167 167 168 
rect 166 168 167 169 
rect 166 193 167 194 
rect 166 198 167 199 
rect 166 199 167 200 
rect 166 210 167 211 
rect 166 262 167 263 
rect 166 263 167 264 
rect 166 289 167 290 
rect 167 40 168 41 
rect 167 49 168 50 
rect 167 65 168 66 
rect 167 67 168 68 
rect 167 81 168 82 
rect 167 88 168 89 
rect 167 193 168 194 
rect 167 195 168 196 
rect 167 196 168 197 
rect 167 197 168 198 
rect 167 198 168 199 
rect 167 210 168 211 
rect 167 261 168 262 
rect 167 262 168 263 
rect 167 289 168 290 
rect 168 25 169 26 
rect 168 26 169 27 
rect 168 27 169 28 
rect 168 28 169 29 
rect 168 29 169 30 
rect 168 30 169 31 
rect 168 31 169 32 
rect 168 32 169 33 
rect 168 33 169 34 
rect 168 34 169 35 
rect 168 35 169 36 
rect 168 36 169 37 
rect 168 37 169 38 
rect 168 38 169 39 
rect 168 39 169 40 
rect 168 40 169 41 
rect 168 49 169 50 
rect 168 65 169 66 
rect 168 67 169 68 
rect 168 81 169 82 
rect 168 88 169 89 
rect 168 144 169 145 
rect 168 145 169 146 
rect 168 146 169 147 
rect 168 147 169 148 
rect 168 148 169 149 
rect 168 149 169 150 
rect 168 150 169 151 
rect 168 151 169 152 
rect 168 152 169 153 
rect 168 153 169 154 
rect 168 154 169 155 
rect 168 155 169 156 
rect 168 156 169 157 
rect 168 157 169 158 
rect 168 158 169 159 
rect 168 159 169 160 
rect 168 160 169 161 
rect 168 161 169 162 
rect 168 162 169 163 
rect 168 163 169 164 
rect 168 164 169 165 
rect 168 165 169 166 
rect 168 166 169 167 
rect 168 167 169 168 
rect 168 168 169 169 
rect 168 169 169 170 
rect 168 170 169 171 
rect 168 171 169 172 
rect 168 172 169 173 
rect 168 173 169 174 
rect 168 174 169 175 
rect 168 175 169 176 
rect 168 176 169 177 
rect 168 177 169 178 
rect 168 178 169 179 
rect 168 179 169 180 
rect 168 180 169 181 
rect 168 181 169 182 
rect 168 182 169 183 
rect 168 183 169 184 
rect 168 184 169 185 
rect 168 193 169 194 
rect 168 195 169 196 
rect 168 210 169 211 
rect 168 217 169 218 
rect 168 218 169 219 
rect 168 249 169 250 
rect 168 250 169 251 
rect 168 251 169 252 
rect 168 252 169 253 
rect 168 253 169 254 
rect 168 254 169 255 
rect 168 255 169 256 
rect 168 256 169 257 
rect 168 257 169 258 
rect 168 258 169 259 
rect 168 259 169 260 
rect 168 260 169 261 
rect 168 261 169 262 
rect 168 263 169 264 
rect 168 264 169 265 
rect 168 265 169 266 
rect 168 266 169 267 
rect 168 267 169 268 
rect 168 268 169 269 
rect 168 269 169 270 
rect 168 270 169 271 
rect 168 271 169 272 
rect 168 272 169 273 
rect 168 273 169 274 
rect 168 274 169 275 
rect 168 275 169 276 
rect 168 276 169 277 
rect 168 277 169 278 
rect 168 278 169 279 
rect 168 279 169 280 
rect 168 280 169 281 
rect 168 281 169 282 
rect 168 289 169 290 
rect 169 24 170 25 
rect 169 25 170 26 
rect 169 49 170 50 
rect 169 65 170 66 
rect 169 67 170 68 
rect 169 81 170 82 
rect 169 88 170 89 
rect 169 184 170 185 
rect 169 193 170 194 
rect 169 195 170 196 
rect 169 210 170 211 
rect 169 216 170 217 
rect 169 217 170 218 
rect 169 248 170 249 
rect 169 249 170 250 
rect 169 263 170 264 
rect 169 289 170 290 
rect 170 24 171 25 
rect 170 49 171 50 
rect 170 65 171 66 
rect 170 67 171 68 
rect 170 81 171 82 
rect 170 88 171 89 
rect 170 184 171 185 
rect 170 193 171 194 
rect 170 195 171 196 
rect 170 210 171 211 
rect 170 216 171 217 
rect 170 248 171 249 
rect 170 257 171 258 
rect 170 258 171 259 
rect 170 259 171 260 
rect 170 260 171 261 
rect 170 261 171 262 
rect 170 262 171 263 
rect 170 263 171 264 
rect 170 289 171 290 
rect 171 24 172 25 
rect 171 49 172 50 
rect 171 67 172 68 
rect 171 81 172 82 
rect 171 88 172 89 
rect 171 184 172 185 
rect 171 193 172 194 
rect 171 195 172 196 
rect 171 210 172 211 
rect 171 216 172 217 
rect 171 248 172 249 
rect 171 257 172 258 
rect 171 289 172 290 
rect 172 24 173 25 
rect 172 49 173 50 
rect 172 67 173 68 
rect 172 81 173 82 
rect 172 88 173 89 
rect 172 184 173 185 
rect 172 193 173 194 
rect 172 195 173 196 
rect 172 210 173 211 
rect 172 216 173 217 
rect 172 248 173 249 
rect 172 257 173 258 
rect 172 289 173 290 
rect 173 24 174 25 
rect 173 49 174 50 
rect 173 67 174 68 
rect 173 81 174 82 
rect 173 88 174 89 
rect 173 184 174 185 
rect 173 193 174 194 
rect 173 195 174 196 
rect 173 210 174 211 
rect 173 216 174 217 
rect 173 248 174 249 
rect 173 257 174 258 
rect 173 289 174 290 
rect 174 24 175 25 
rect 174 49 175 50 
rect 174 67 175 68 
rect 174 81 175 82 
rect 174 88 175 89 
rect 174 184 175 185 
rect 174 193 175 194 
rect 174 195 175 196 
rect 174 210 175 211 
rect 174 216 175 217 
rect 174 248 175 249 
rect 174 257 175 258 
rect 174 289 175 290 
rect 175 24 176 25 
rect 175 34 176 35 
rect 175 35 176 36 
rect 175 36 176 37 
rect 175 37 176 38 
rect 175 38 176 39 
rect 175 39 176 40 
rect 175 49 176 50 
rect 175 67 176 68 
rect 175 81 176 82 
rect 175 88 176 89 
rect 175 114 176 115 
rect 175 115 176 116 
rect 175 116 176 117 
rect 175 117 176 118 
rect 175 118 176 119 
rect 175 119 176 120 
rect 175 120 176 121 
rect 175 184 176 185 
rect 175 193 176 194 
rect 175 195 176 196 
rect 175 210 176 211 
rect 175 216 176 217 
rect 175 248 176 249 
rect 175 257 176 258 
rect 175 289 176 290 
rect 176 24 177 25 
rect 176 25 177 26 
rect 176 48 177 49 
rect 176 49 177 50 
rect 176 67 177 68 
rect 176 70 177 71 
rect 176 71 177 72 
rect 176 72 177 73 
rect 176 73 177 74 
rect 176 81 177 82 
rect 176 88 177 89 
rect 176 184 177 185 
rect 176 193 177 194 
rect 176 195 177 196 
rect 176 197 177 198 
rect 176 210 177 211 
rect 176 216 177 217 
rect 176 248 177 249 
rect 176 257 177 258 
rect 176 289 177 290 
rect 177 67 178 68 
rect 177 81 178 82 
rect 177 88 178 89 
rect 177 95 178 96 
rect 177 96 178 97 
rect 177 97 178 98 
rect 177 98 178 99 
rect 177 99 178 100 
rect 177 100 178 101 
rect 177 101 178 102 
rect 177 102 178 103 
rect 177 103 178 104 
rect 177 104 178 105 
rect 177 105 178 106 
rect 177 106 178 107 
rect 177 107 178 108 
rect 177 108 178 109 
rect 177 109 178 110 
rect 177 110 178 111 
rect 177 111 178 112 
rect 177 112 178 113 
rect 177 113 178 114 
rect 177 114 178 115 
rect 177 115 178 116 
rect 177 116 178 117 
rect 177 117 178 118 
rect 177 118 178 119 
rect 177 119 178 120 
rect 177 120 178 121 
rect 177 121 178 122 
rect 177 122 178 123 
rect 177 123 178 124 
rect 177 124 178 125 
rect 177 125 178 126 
rect 177 126 178 127 
rect 177 127 178 128 
rect 177 128 178 129 
rect 177 129 178 130 
rect 177 130 178 131 
rect 177 131 178 132 
rect 177 132 178 133 
rect 177 133 178 134 
rect 177 134 178 135 
rect 177 135 178 136 
rect 177 136 178 137 
rect 177 137 178 138 
rect 177 138 178 139 
rect 177 139 178 140 
rect 177 140 178 141 
rect 177 141 178 142 
rect 177 142 178 143 
rect 177 143 178 144 
rect 177 144 178 145 
rect 177 145 178 146 
rect 177 146 178 147 
rect 177 147 178 148 
rect 177 148 178 149 
rect 177 149 178 150 
rect 177 150 178 151 
rect 177 151 178 152 
rect 177 152 178 153 
rect 177 153 178 154 
rect 177 154 178 155 
rect 177 155 178 156 
rect 177 156 178 157 
rect 177 157 178 158 
rect 177 158 178 159 
rect 177 159 178 160 
rect 177 160 178 161 
rect 177 161 178 162 
rect 177 162 178 163 
rect 177 163 178 164 
rect 177 164 178 165 
rect 177 165 178 166 
rect 177 166 178 167 
rect 177 167 178 168 
rect 177 168 178 169 
rect 177 184 178 185 
rect 177 193 178 194 
rect 177 195 178 196 
rect 177 197 178 198 
rect 177 210 178 211 
rect 177 216 178 217 
rect 177 248 178 249 
rect 177 257 178 258 
rect 177 262 178 263 
rect 177 263 178 264 
rect 177 264 178 265 
rect 177 265 178 266 
rect 177 266 178 267 
rect 177 267 178 268 
rect 177 268 178 269 
rect 177 269 178 270 
rect 177 270 178 271 
rect 177 271 178 272 
rect 177 272 178 273 
rect 177 273 178 274 
rect 177 274 178 275 
rect 177 275 178 276 
rect 177 276 178 277 
rect 177 277 178 278 
rect 177 278 178 279 
rect 177 279 178 280 
rect 177 280 178 281 
rect 177 281 178 282 
rect 177 282 178 283 
rect 177 289 178 290 
rect 178 57 179 58 
rect 178 67 179 68 
rect 178 81 179 82 
rect 178 88 179 89 
rect 178 184 179 185 
rect 178 193 179 194 
rect 178 195 179 196 
rect 178 197 179 198 
rect 178 216 179 217 
rect 178 248 179 249 
rect 178 257 179 258 
rect 178 289 179 290 
rect 179 57 180 58 
rect 179 65 180 66 
rect 179 67 180 68 
rect 179 70 180 71 
rect 179 71 180 72 
rect 179 72 180 73 
rect 179 73 180 74 
rect 179 74 180 75 
rect 179 75 180 76 
rect 179 76 180 77 
rect 179 81 180 82 
rect 179 88 180 89 
rect 179 184 180 185 
rect 179 193 180 194 
rect 179 195 180 196 
rect 179 197 180 198 
rect 179 216 180 217 
rect 179 248 180 249 
rect 179 257 180 258 
rect 179 289 180 290 
rect 180 57 181 58 
rect 180 65 181 66 
rect 180 67 181 68 
rect 180 81 181 82 
rect 180 88 181 89 
rect 180 184 181 185 
rect 180 193 181 194 
rect 180 197 181 198 
rect 180 216 181 217 
rect 180 247 181 248 
rect 180 248 181 249 
rect 180 251 181 252 
rect 180 257 181 258 
rect 180 289 181 290 
rect 181 57 182 58 
rect 181 65 182 66 
rect 181 67 182 68 
rect 181 81 182 82 
rect 181 88 182 89 
rect 181 184 182 185 
rect 181 193 182 194 
rect 181 197 182 198 
rect 181 216 182 217 
rect 181 246 182 247 
rect 181 247 182 248 
rect 181 250 182 251 
rect 181 251 182 252 
rect 181 256 182 257 
rect 181 257 182 258 
rect 181 289 182 290 
rect 182 57 183 58 
rect 182 65 183 66 
rect 182 67 183 68 
rect 182 81 183 82 
rect 182 88 183 89 
rect 182 112 183 113 
rect 182 113 183 114 
rect 182 114 183 115 
rect 182 115 183 116 
rect 182 116 183 117 
rect 182 117 183 118 
rect 182 118 183 119 
rect 182 119 183 120 
rect 182 120 183 121 
rect 182 121 183 122 
rect 182 122 183 123 
rect 182 123 183 124 
rect 182 124 183 125 
rect 182 125 183 126 
rect 182 126 183 127 
rect 182 127 183 128 
rect 182 128 183 129 
rect 182 129 183 130 
rect 182 130 183 131 
rect 182 131 183 132 
rect 182 132 183 133 
rect 182 133 183 134 
rect 182 134 183 135 
rect 182 135 183 136 
rect 182 136 183 137 
rect 182 137 183 138 
rect 182 138 183 139 
rect 182 139 183 140 
rect 182 140 183 141 
rect 182 141 183 142 
rect 182 142 183 143 
rect 182 143 183 144 
rect 182 144 183 145 
rect 182 145 183 146 
rect 182 146 183 147 
rect 182 147 183 148 
rect 182 148 183 149 
rect 182 149 183 150 
rect 182 150 183 151 
rect 182 151 183 152 
rect 182 152 183 153 
rect 182 153 183 154 
rect 182 154 183 155 
rect 182 155 183 156 
rect 182 156 183 157 
rect 182 157 183 158 
rect 182 158 183 159 
rect 182 159 183 160 
rect 182 160 183 161 
rect 182 161 183 162 
rect 182 162 183 163 
rect 182 163 183 164 
rect 182 184 183 185 
rect 182 193 183 194 
rect 182 197 183 198 
rect 182 216 183 217 
rect 182 232 183 233 
rect 182 233 183 234 
rect 182 234 183 235 
rect 182 246 183 247 
rect 182 248 183 249 
rect 182 249 183 250 
rect 182 250 183 251 
rect 182 256 183 257 
rect 182 262 183 263 
rect 182 263 183 264 
rect 182 264 183 265 
rect 182 265 183 266 
rect 182 266 183 267 
rect 182 267 183 268 
rect 182 268 183 269 
rect 182 269 183 270 
rect 182 270 183 271 
rect 182 271 183 272 
rect 182 272 183 273 
rect 182 273 183 274 
rect 182 289 183 290 
rect 183 35 184 36 
rect 183 36 184 37 
rect 183 37 184 38 
rect 183 38 184 39 
rect 183 39 184 40 
rect 183 40 184 41 
rect 183 41 184 42 
rect 183 42 184 43 
rect 183 43 184 44 
rect 183 44 184 45 
rect 183 45 184 46 
rect 183 46 184 47 
rect 183 47 184 48 
rect 183 48 184 49 
rect 183 49 184 50 
rect 183 50 184 51 
rect 183 51 184 52 
rect 183 52 184 53 
rect 183 57 184 58 
rect 183 65 184 66 
rect 183 67 184 68 
rect 183 81 184 82 
rect 183 83 184 84 
rect 183 85 184 86 
rect 183 88 184 89 
rect 183 111 184 112 
rect 183 112 184 113 
rect 183 184 184 185 
rect 183 193 184 194 
rect 183 197 184 198 
rect 183 216 184 217 
rect 183 231 184 232 
rect 183 232 184 233 
rect 183 246 184 247 
rect 183 248 184 249 
rect 183 256 184 257 
rect 183 289 184 290 
rect 184 16 185 17 
rect 184 17 185 18 
rect 184 32 185 33 
rect 184 57 185 58 
rect 184 65 185 66 
rect 184 67 185 68 
rect 184 81 185 82 
rect 184 83 185 84 
rect 184 85 185 86 
rect 184 88 185 89 
rect 184 96 185 97 
rect 184 97 185 98 
rect 184 98 185 99 
rect 184 99 185 100 
rect 184 100 185 101 
rect 184 101 185 102 
rect 184 102 185 103 
rect 184 103 185 104 
rect 184 104 185 105 
rect 184 105 185 106 
rect 184 106 185 107 
rect 184 107 185 108 
rect 184 108 185 109 
rect 184 109 185 110 
rect 184 110 185 111 
rect 184 111 185 112 
rect 184 114 185 115 
rect 184 115 185 116 
rect 184 116 185 117 
rect 184 117 185 118 
rect 184 118 185 119 
rect 184 119 185 120 
rect 184 120 185 121 
rect 184 141 185 142 
rect 184 142 185 143 
rect 184 143 185 144 
rect 184 144 185 145 
rect 184 145 185 146 
rect 184 146 185 147 
rect 184 147 185 148 
rect 184 148 185 149 
rect 184 149 185 150 
rect 184 150 185 151 
rect 184 151 185 152 
rect 184 152 185 153 
rect 184 153 185 154 
rect 184 154 185 155 
rect 184 155 185 156 
rect 184 156 185 157 
rect 184 157 185 158 
rect 184 158 185 159 
rect 184 159 185 160 
rect 184 160 185 161 
rect 184 161 185 162 
rect 184 162 185 163 
rect 184 163 185 164 
rect 184 164 185 165 
rect 184 165 185 166 
rect 184 166 185 167 
rect 184 167 185 168 
rect 184 168 185 169 
rect 184 169 185 170 
rect 184 170 185 171 
rect 184 171 185 172 
rect 184 172 185 173 
rect 184 173 185 174 
rect 184 174 185 175 
rect 184 175 185 176 
rect 184 176 185 177 
rect 184 177 185 178 
rect 184 178 185 179 
rect 184 179 185 180 
rect 184 184 185 185 
rect 184 193 185 194 
rect 184 197 185 198 
rect 184 216 185 217 
rect 184 226 185 227 
rect 184 229 185 230 
rect 184 230 185 231 
rect 184 231 185 232 
rect 184 233 185 234 
rect 184 234 185 235 
rect 184 235 185 236 
rect 184 236 185 237 
rect 184 237 185 238 
rect 184 238 185 239 
rect 184 239 185 240 
rect 184 240 185 241 
rect 184 241 185 242 
rect 184 242 185 243 
rect 184 243 185 244 
rect 184 246 185 247 
rect 184 248 185 249 
rect 184 256 185 257 
rect 184 259 185 260 
rect 184 260 185 261 
rect 184 261 185 262 
rect 184 262 185 263 
rect 184 263 185 264 
rect 184 264 185 265 
rect 184 265 185 266 
rect 184 266 185 267 
rect 184 289 185 290 
rect 185 17 186 18 
rect 185 32 186 33 
rect 185 33 186 34 
rect 185 34 186 35 
rect 185 35 186 36 
rect 185 36 186 37 
rect 185 37 186 38 
rect 185 57 186 58 
rect 185 65 186 66 
rect 185 67 186 68 
rect 185 81 186 82 
rect 185 83 186 84 
rect 185 85 186 86 
rect 185 88 186 89 
rect 185 184 186 185 
rect 185 193 186 194 
rect 185 197 186 198 
rect 185 216 186 217 
rect 185 226 186 227 
rect 185 228 186 229 
rect 185 229 186 230 
rect 185 232 186 233 
rect 185 233 186 234 
rect 185 246 186 247 
rect 185 248 186 249 
rect 185 256 186 257 
rect 185 289 186 290 
rect 186 17 187 18 
rect 186 37 187 38 
rect 186 38 187 39 
rect 186 39 187 40 
rect 186 40 187 41 
rect 186 65 187 66 
rect 186 67 187 68 
rect 186 81 187 82 
rect 186 83 187 84 
rect 186 85 187 86 
rect 186 88 187 89 
rect 186 184 187 185 
rect 186 193 187 194 
rect 186 197 187 198 
rect 186 216 187 217 
rect 186 226 187 227 
rect 186 228 187 229 
rect 186 231 187 232 
rect 186 232 187 233 
rect 186 246 187 247 
rect 186 248 187 249 
rect 186 289 187 290 
rect 187 17 188 18 
rect 187 40 188 41 
rect 187 65 188 66 
rect 187 67 188 68 
rect 187 81 188 82 
rect 187 83 188 84 
rect 187 85 188 86 
rect 187 88 188 89 
rect 187 184 188 185 
rect 187 193 188 194 
rect 187 197 188 198 
rect 187 216 188 217 
rect 187 226 188 227 
rect 187 228 188 229 
rect 187 246 188 247 
rect 187 248 188 249 
rect 187 289 188 290 
rect 188 17 189 18 
rect 188 40 189 41 
rect 188 65 189 66 
rect 188 67 189 68 
rect 188 81 189 82 
rect 188 83 189 84 
rect 188 85 189 86 
rect 188 88 189 89 
rect 188 184 189 185 
rect 188 193 189 194 
rect 188 197 189 198 
rect 188 216 189 217 
rect 188 226 189 227 
rect 188 228 189 229 
rect 188 246 189 247 
rect 188 248 189 249 
rect 188 289 189 290 
rect 189 17 190 18 
rect 189 40 190 41 
rect 189 65 190 66 
rect 189 67 190 68 
rect 189 81 190 82 
rect 189 83 190 84 
rect 189 85 190 86 
rect 189 88 190 89 
rect 189 184 190 185 
rect 189 193 190 194 
rect 189 197 190 198 
rect 189 216 190 217 
rect 189 226 190 227 
rect 189 228 190 229 
rect 189 246 190 247 
rect 189 248 190 249 
rect 189 289 190 290 
rect 190 17 191 18 
rect 190 40 191 41 
rect 190 65 191 66 
rect 190 67 191 68 
rect 190 81 191 82 
rect 190 83 191 84 
rect 190 85 191 86 
rect 190 88 191 89 
rect 190 184 191 185 
rect 190 193 191 194 
rect 190 197 191 198 
rect 190 216 191 217 
rect 190 226 191 227 
rect 190 228 191 229 
rect 190 246 191 247 
rect 190 248 191 249 
rect 190 289 191 290 
rect 191 17 192 18 
rect 191 22 192 23 
rect 191 23 192 24 
rect 191 24 192 25 
rect 191 40 192 41 
rect 191 65 192 66 
rect 191 67 192 68 
rect 191 81 192 82 
rect 191 83 192 84 
rect 191 85 192 86 
rect 191 86 192 87 
rect 191 88 192 89 
rect 191 162 192 163 
rect 191 184 192 185 
rect 191 193 192 194 
rect 191 197 192 198 
rect 191 216 192 217 
rect 191 226 192 227 
rect 191 228 192 229 
rect 191 246 192 247 
rect 191 248 192 249 
rect 191 289 192 290 
rect 192 17 193 18 
rect 192 24 193 25 
rect 192 25 193 26 
rect 192 34 193 35 
rect 192 35 193 36 
rect 192 36 193 37 
rect 192 37 193 38 
rect 192 40 193 41 
rect 192 41 193 42 
rect 192 65 193 66 
rect 192 67 193 68 
rect 192 70 193 71 
rect 192 71 193 72 
rect 192 72 193 73 
rect 192 73 193 74 
rect 192 81 193 82 
rect 192 83 193 84 
rect 192 86 193 87 
rect 192 88 193 89 
rect 192 89 193 90 
rect 192 161 193 162 
rect 192 162 193 163 
rect 192 184 193 185 
rect 192 193 193 194 
rect 192 197 193 198 
rect 192 216 193 217 
rect 192 226 193 227 
rect 192 228 193 229 
rect 192 246 193 247 
rect 192 248 193 249 
rect 192 258 193 259 
rect 192 259 193 260 
rect 192 260 193 261 
rect 192 261 193 262 
rect 192 277 193 278 
rect 192 279 193 280 
rect 192 289 193 290 
rect 192 291 193 292 
rect 192 293 193 294 
rect 193 41 194 42 
rect 193 42 194 43 
rect 193 65 194 66 
rect 193 67 194 68 
rect 193 68 194 69 
rect 193 81 194 82 
rect 193 83 194 84 
rect 193 86 194 87 
rect 193 87 194 88 
rect 193 89 194 90 
rect 193 90 194 91 
rect 193 92 194 93 
rect 193 93 194 94 
rect 193 94 194 95 
rect 193 95 194 96 
rect 193 96 194 97 
rect 193 97 194 98 
rect 193 98 194 99 
rect 193 99 194 100 
rect 193 100 194 101 
rect 193 101 194 102 
rect 193 102 194 103 
rect 193 103 194 104 
rect 193 104 194 105 
rect 193 105 194 106 
rect 193 106 194 107 
rect 193 107 194 108 
rect 193 108 194 109 
rect 193 109 194 110 
rect 193 110 194 111 
rect 193 111 194 112 
rect 193 112 194 113 
rect 193 113 194 114 
rect 193 114 194 115 
rect 193 115 194 116 
rect 193 116 194 117 
rect 193 117 194 118 
rect 193 118 194 119 
rect 193 119 194 120 
rect 193 152 194 153 
rect 193 161 194 162 
rect 193 163 194 164 
rect 193 164 194 165 
rect 193 165 194 166 
rect 193 166 194 167 
rect 193 167 194 168 
rect 193 168 194 169 
rect 193 169 194 170 
rect 193 170 194 171 
rect 193 171 194 172 
rect 193 172 194 173 
rect 193 184 194 185 
rect 193 193 194 194 
rect 193 197 194 198 
rect 193 216 194 217 
rect 193 226 194 227 
rect 193 228 194 229 
rect 193 230 194 231 
rect 193 231 194 232 
rect 193 232 194 233 
rect 193 233 194 234 
rect 193 246 194 247 
rect 193 248 194 249 
rect 193 258 194 259 
rect 193 272 194 273 
rect 193 273 194 274 
rect 193 274 194 275 
rect 193 275 194 276 
rect 193 277 194 278 
rect 193 279 194 280 
rect 193 289 194 290 
rect 193 291 194 292 
rect 193 293 194 294 
rect 193 303 194 304 
rect 193 304 194 305 
rect 193 305 194 306 
rect 193 306 194 307 
rect 194 81 195 82 
rect 194 83 195 84 
rect 194 87 195 88 
rect 194 88 195 89 
rect 194 90 195 91 
rect 194 152 195 153 
rect 194 161 195 162 
rect 194 162 195 163 
rect 194 184 195 185 
rect 194 193 195 194 
rect 194 197 195 198 
rect 194 216 195 217 
rect 194 225 195 226 
rect 194 226 195 227 
rect 194 246 195 247 
rect 194 248 195 249 
rect 194 258 195 259 
rect 194 276 195 277 
rect 194 277 195 278 
rect 194 279 195 280 
rect 194 289 195 290 
rect 194 291 195 292 
rect 194 293 195 294 
rect 195 81 196 82 
rect 195 83 196 84 
rect 195 88 196 89 
rect 195 90 196 91 
rect 195 93 196 94 
rect 195 94 196 95 
rect 195 95 196 96 
rect 195 96 196 97 
rect 195 97 196 98 
rect 195 98 196 99 
rect 195 99 196 100 
rect 195 152 196 153 
rect 195 162 196 163 
rect 195 163 196 164 
rect 195 184 196 185 
rect 195 193 196 194 
rect 195 197 196 198 
rect 195 216 196 217 
rect 195 224 196 225 
rect 195 225 196 226 
rect 195 246 196 247 
rect 195 248 196 249 
rect 195 258 196 259 
rect 195 260 196 261 
rect 195 271 196 272 
rect 195 272 196 273 
rect 195 273 196 274 
rect 195 274 196 275 
rect 195 275 196 276 
rect 195 276 196 277 
rect 195 278 196 279 
rect 195 279 196 280 
rect 195 289 196 290 
rect 195 291 196 292 
rect 195 293 196 294 
rect 196 81 197 82 
rect 196 83 197 84 
rect 196 88 197 89 
rect 196 90 197 91 
rect 196 152 197 153 
rect 196 163 197 164 
rect 196 193 197 194 
rect 196 197 197 198 
rect 196 216 197 217 
rect 196 224 197 225 
rect 196 226 197 227 
rect 196 227 197 228 
rect 196 228 197 229 
rect 196 229 197 230 
rect 196 230 197 231 
rect 196 231 197 232 
rect 196 232 197 233 
rect 196 233 197 234 
rect 196 246 197 247 
rect 196 248 197 249 
rect 196 258 197 259 
rect 196 260 197 261 
rect 196 277 197 278 
rect 196 278 197 279 
rect 196 291 197 292 
rect 196 293 197 294 
rect 197 81 198 82 
rect 197 83 198 84 
rect 197 88 198 89 
rect 197 90 198 91 
rect 197 91 198 92 
rect 197 92 198 93 
rect 197 93 198 94 
rect 197 94 198 95 
rect 197 95 198 96 
rect 197 96 198 97 
rect 197 97 198 98 
rect 197 98 198 99 
rect 197 99 198 100 
rect 197 152 198 153 
rect 197 163 198 164 
rect 197 193 198 194 
rect 197 197 198 198 
rect 197 216 198 217 
rect 197 224 198 225 
rect 197 225 198 226 
rect 197 246 198 247 
rect 197 248 198 249 
rect 197 258 198 259 
rect 197 260 198 261 
rect 197 262 198 263 
rect 197 263 198 264 
rect 197 264 198 265 
rect 197 265 198 266 
rect 197 266 198 267 
rect 197 267 198 268 
rect 197 268 198 269 
rect 197 269 198 270 
rect 197 270 198 271 
rect 197 271 198 272 
rect 197 272 198 273 
rect 197 273 198 274 
rect 197 274 198 275 
rect 197 275 198 276 
rect 197 276 198 277 
rect 197 277 198 278 
rect 197 291 198 292 
rect 197 293 198 294 
rect 198 83 199 84 
rect 198 88 199 89 
rect 198 89 199 90 
rect 198 152 199 153 
rect 198 163 199 164 
rect 198 193 199 194 
rect 198 197 199 198 
rect 198 216 199 217 
rect 198 225 199 226 
rect 198 226 199 227 
rect 198 227 199 228 
rect 198 228 199 229 
rect 198 229 199 230 
rect 198 230 199 231 
rect 198 231 199 232 
rect 198 232 199 233 
rect 198 233 199 234 
rect 198 234 199 235 
rect 198 235 199 236 
rect 198 236 199 237 
rect 198 237 199 238 
rect 198 238 199 239 
rect 198 239 199 240 
rect 198 240 199 241 
rect 198 241 199 242 
rect 198 242 199 243 
rect 198 243 199 244 
rect 198 244 199 245 
rect 198 246 199 247 
rect 198 248 199 249 
rect 198 258 199 259 
rect 198 260 199 261 
rect 198 261 199 262 
rect 198 291 199 292 
rect 198 293 199 294 
rect 199 83 200 84 
rect 199 89 200 90 
rect 199 90 200 91 
rect 199 91 200 92 
rect 199 92 200 93 
rect 199 93 200 94 
rect 199 94 200 95 
rect 199 95 200 96 
rect 199 96 200 97 
rect 199 97 200 98 
rect 199 98 200 99 
rect 199 99 200 100 
rect 199 100 200 101 
rect 199 101 200 102 
rect 199 102 200 103 
rect 199 152 200 153 
rect 199 161 200 162 
rect 199 163 200 164 
rect 199 193 200 194 
rect 199 197 200 198 
rect 199 216 200 217 
rect 199 248 200 249 
rect 199 261 200 262 
rect 199 262 200 263 
rect 199 263 200 264 
rect 199 264 200 265 
rect 199 291 200 292 
rect 199 293 200 294 
rect 200 83 201 84 
rect 200 152 201 153 
rect 200 161 201 162 
rect 200 163 201 164 
rect 200 193 201 194 
rect 200 197 201 198 
rect 200 216 201 217 
rect 200 248 201 249 
rect 200 264 201 265 
rect 200 291 201 292 
rect 200 293 201 294 
rect 201 83 202 84 
rect 201 152 202 153 
rect 201 161 202 162 
rect 201 163 202 164 
rect 201 193 202 194 
rect 201 197 202 198 
rect 201 216 202 217 
rect 201 248 202 249 
rect 201 264 202 265 
rect 201 291 202 292 
rect 201 293 202 294 
rect 202 83 203 84 
rect 202 152 203 153 
rect 202 161 203 162 
rect 202 163 203 164 
rect 202 193 203 194 
rect 202 197 203 198 
rect 202 216 203 217 
rect 202 248 203 249 
rect 202 264 203 265 
rect 202 291 203 292 
rect 202 293 203 294 
rect 203 83 204 84 
rect 203 152 204 153 
rect 203 161 204 162 
rect 203 163 204 164 
rect 203 193 204 194 
rect 203 197 204 198 
rect 203 216 204 217 
rect 203 248 204 249 
rect 203 264 204 265 
rect 203 291 204 292 
rect 203 293 204 294 
rect 204 83 205 84 
rect 204 152 205 153 
rect 204 161 205 162 
rect 204 163 205 164 
rect 204 193 205 194 
rect 204 197 205 198 
rect 204 216 205 217 
rect 204 248 205 249 
rect 204 291 205 292 
rect 204 293 205 294 
rect 205 83 206 84 
rect 205 152 206 153 
rect 205 161 206 162 
rect 205 163 206 164 
rect 205 193 206 194 
rect 205 197 206 198 
rect 205 216 206 217 
rect 205 248 206 249 
rect 205 291 206 292 
rect 205 293 206 294 
rect 206 83 207 84 
rect 206 152 207 153 
rect 206 161 207 162 
rect 206 163 207 164 
rect 206 193 207 194 
rect 206 197 207 198 
rect 206 216 207 217 
rect 206 248 207 249 
rect 206 273 207 274 
rect 206 274 207 275 
rect 206 291 207 292 
rect 206 293 207 294 
rect 207 83 208 84 
rect 207 152 208 153 
rect 207 161 208 162 
rect 207 163 208 164 
rect 207 193 208 194 
rect 207 197 208 198 
rect 207 216 208 217 
rect 207 248 208 249 
rect 207 273 208 274 
rect 207 291 208 292 
rect 207 293 208 294 
rect 208 83 209 84 
rect 208 152 209 153 
rect 208 161 209 162 
rect 208 163 209 164 
rect 208 193 209 194 
rect 208 197 209 198 
rect 208 216 209 217 
rect 208 248 209 249 
rect 208 273 209 274 
rect 208 291 209 292 
rect 208 293 209 294 
rect 209 83 210 84 
rect 209 152 210 153 
rect 209 161 210 162 
rect 209 163 210 164 
rect 209 165 210 166 
rect 209 184 210 185 
rect 209 193 210 194 
rect 209 197 210 198 
rect 209 216 210 217 
rect 209 248 210 249 
rect 209 273 210 274 
rect 209 291 210 292 
rect 209 293 210 294 
rect 210 83 211 84 
rect 210 152 211 153 
rect 210 161 211 162 
rect 210 163 211 164 
rect 210 165 211 166 
rect 210 183 211 184 
rect 210 184 211 185 
rect 210 193 211 194 
rect 210 197 211 198 
rect 210 216 211 217 
rect 210 248 211 249 
rect 210 271 211 272 
rect 210 272 211 273 
rect 210 273 211 274 
rect 210 291 211 292 
rect 210 293 211 294 
rect 210 294 211 295 
rect 210 295 211 296 
rect 210 296 211 297 
rect 210 297 211 298 
rect 210 298 211 299 
rect 210 299 211 300 
rect 210 300 211 301 
rect 210 301 211 302 
rect 210 303 211 304 
rect 210 304 211 305 
rect 210 305 211 306 
rect 210 306 211 307 
rect 211 83 212 84 
rect 211 152 212 153 
rect 211 161 212 162 
rect 211 163 212 164 
rect 211 165 212 166 
rect 211 183 212 184 
rect 211 193 212 194 
rect 211 197 212 198 
rect 211 216 212 217 
rect 211 248 212 249 
rect 211 291 212 292 
rect 211 301 212 302 
rect 211 302 212 303 
rect 212 83 213 84 
rect 212 152 213 153 
rect 212 161 213 162 
rect 212 163 213 164 
rect 212 165 213 166 
rect 212 183 213 184 
rect 212 193 213 194 
rect 212 197 213 198 
rect 212 216 213 217 
rect 212 225 213 226 
rect 212 226 213 227 
rect 212 227 213 228 
rect 212 228 213 229 
rect 212 229 213 230 
rect 212 230 213 231 
rect 212 231 213 232 
rect 212 232 213 233 
rect 212 233 213 234 
rect 212 234 213 235 
rect 212 235 213 236 
rect 212 236 213 237 
rect 212 237 213 238 
rect 212 238 213 239 
rect 212 239 213 240 
rect 212 240 213 241 
rect 212 241 213 242 
rect 212 242 213 243 
rect 212 248 213 249 
rect 212 254 213 255 
rect 212 255 213 256 
rect 212 256 213 257 
rect 212 257 213 258 
rect 212 258 213 259 
rect 212 259 213 260 
rect 212 260 213 261 
rect 212 261 213 262 
rect 212 262 213 263 
rect 212 263 213 264 
rect 212 264 213 265 
rect 212 265 213 266 
rect 212 266 213 267 
rect 212 267 213 268 
rect 212 268 213 269 
rect 212 269 213 270 
rect 212 270 213 271 
rect 212 271 213 272 
rect 212 272 213 273 
rect 212 273 213 274 
rect 212 274 213 275 
rect 212 275 213 276 
rect 212 276 213 277 
rect 212 277 213 278 
rect 212 278 213 279 
rect 212 291 213 292 
rect 212 302 213 303 
rect 212 303 213 304 
rect 212 304 213 305 
rect 212 305 213 306 
rect 212 306 213 307 
rect 212 307 213 308 
rect 212 308 213 309 
rect 212 309 213 310 
rect 213 83 214 84 
rect 213 152 214 153 
rect 213 161 214 162 
rect 213 163 214 164 
rect 213 165 214 166 
rect 213 183 214 184 
rect 213 193 214 194 
rect 213 197 214 198 
rect 213 216 214 217 
rect 213 225 214 226 
rect 213 248 214 249 
rect 213 291 214 292 
rect 213 309 214 310 
rect 214 83 215 84 
rect 214 115 215 116 
rect 214 116 215 117 
rect 214 117 215 118 
rect 214 118 215 119 
rect 214 119 215 120 
rect 214 120 215 121 
rect 214 121 215 122 
rect 214 122 215 123 
rect 214 123 215 124 
rect 214 124 215 125 
rect 214 125 215 126 
rect 214 126 215 127 
rect 214 127 215 128 
rect 214 128 215 129 
rect 214 129 215 130 
rect 214 130 215 131 
rect 214 131 215 132 
rect 214 132 215 133 
rect 214 133 215 134 
rect 214 134 215 135 
rect 214 135 215 136 
rect 214 136 215 137 
rect 214 137 215 138 
rect 214 138 215 139 
rect 214 139 215 140 
rect 214 140 215 141 
rect 214 141 215 142 
rect 214 142 215 143 
rect 214 143 215 144 
rect 214 144 215 145 
rect 214 145 215 146 
rect 214 146 215 147 
rect 214 147 215 148 
rect 214 148 215 149 
rect 214 149 215 150 
rect 214 150 215 151 
rect 214 152 215 153 
rect 214 161 215 162 
rect 214 163 215 164 
rect 214 165 215 166 
rect 214 183 215 184 
rect 214 193 215 194 
rect 214 197 215 198 
rect 214 216 215 217 
rect 214 225 215 226 
rect 214 231 215 232 
rect 214 232 215 233 
rect 214 233 215 234 
rect 214 234 215 235 
rect 214 235 215 236 
rect 214 236 215 237 
rect 214 237 215 238 
rect 214 238 215 239 
rect 214 239 215 240 
rect 214 240 215 241 
rect 214 241 215 242 
rect 214 242 215 243 
rect 214 243 215 244 
rect 214 248 215 249 
rect 214 253 215 254 
rect 214 254 215 255 
rect 214 255 215 256 
rect 214 256 215 257 
rect 214 257 215 258 
rect 214 258 215 259 
rect 214 259 215 260 
rect 214 260 215 261 
rect 214 261 215 262 
rect 214 262 215 263 
rect 214 263 215 264 
rect 214 264 215 265 
rect 214 265 215 266 
rect 214 291 215 292 
rect 214 309 215 310 
rect 215 83 216 84 
rect 215 152 216 153 
rect 215 165 216 166 
rect 215 183 216 184 
rect 215 193 216 194 
rect 215 197 216 198 
rect 215 216 216 217 
rect 215 225 216 226 
rect 215 248 216 249 
rect 215 291 216 292 
rect 216 83 217 84 
rect 216 115 217 116 
rect 216 116 217 117 
rect 216 117 217 118 
rect 216 118 217 119 
rect 216 119 217 120 
rect 216 120 217 121 
rect 216 152 217 153 
rect 216 165 217 166 
rect 216 183 217 184 
rect 216 193 217 194 
rect 216 197 217 198 
rect 216 216 217 217 
rect 216 225 217 226 
rect 216 240 217 241 
rect 216 241 217 242 
rect 216 242 217 243 
rect 216 248 217 249 
rect 216 256 217 257 
rect 216 257 217 258 
rect 216 291 217 292 
rect 217 83 218 84 
rect 217 152 218 153 
rect 217 165 218 166 
rect 217 183 218 184 
rect 217 193 218 194 
rect 217 216 218 217 
rect 217 225 218 226 
rect 217 242 218 243 
rect 217 248 218 249 
rect 217 257 218 258 
rect 217 291 218 292 
rect 218 83 219 84 
rect 218 152 219 153 
rect 218 165 219 166 
rect 218 183 219 184 
rect 218 193 219 194 
rect 218 216 219 217 
rect 218 225 219 226 
rect 218 242 219 243 
rect 218 248 219 249 
rect 218 257 219 258 
rect 218 291 219 292 
rect 218 293 219 294 
rect 218 294 219 295 
rect 218 295 219 296 
rect 219 83 220 84 
rect 219 152 220 153 
rect 219 165 220 166 
rect 219 183 220 184 
rect 219 193 220 194 
rect 219 216 220 217 
rect 219 225 220 226 
rect 219 242 220 243 
rect 219 248 220 249 
rect 219 257 220 258 
rect 219 291 220 292 
rect 219 293 220 294 
rect 220 82 221 83 
rect 220 83 221 84 
rect 220 152 221 153 
rect 220 165 221 166 
rect 220 183 221 184 
rect 220 193 221 194 
rect 220 216 221 217 
rect 220 225 221 226 
rect 220 242 221 243 
rect 220 248 221 249 
rect 220 257 221 258 
rect 220 291 221 292 
rect 220 293 221 294 
rect 221 82 222 83 
rect 221 152 222 153 
rect 221 165 222 166 
rect 221 183 222 184 
rect 221 193 222 194 
rect 221 216 222 217 
rect 221 225 222 226 
rect 221 242 222 243 
rect 221 248 222 249 
rect 221 257 222 258 
rect 221 292 222 293 
rect 221 293 222 294 
rect 222 82 223 83 
rect 222 84 223 85 
rect 222 152 223 153 
rect 222 165 223 166 
rect 222 183 223 184 
rect 222 193 223 194 
rect 222 216 223 217 
rect 222 225 223 226 
rect 222 242 223 243 
rect 222 248 223 249 
rect 222 257 223 258 
rect 222 289 223 290 
rect 222 290 223 291 
rect 222 291 223 292 
rect 222 292 223 293 
rect 223 82 224 83 
rect 223 84 224 85 
rect 223 152 224 153 
rect 223 165 224 166 
rect 223 183 224 184 
rect 223 193 224 194 
rect 223 216 224 217 
rect 223 225 224 226 
rect 223 242 224 243 
rect 223 248 224 249 
rect 223 257 224 258 
rect 223 289 224 290 
rect 224 56 225 57 
rect 224 82 225 83 
rect 224 84 225 85 
rect 224 152 225 153 
rect 224 165 225 166 
rect 224 168 225 169 
rect 224 183 225 184 
rect 224 193 225 194 
rect 224 200 225 201 
rect 224 216 225 217 
rect 224 224 225 225 
rect 224 225 225 226 
rect 224 242 225 243 
rect 224 248 225 249 
rect 224 257 225 258 
rect 224 288 225 289 
rect 224 289 225 290 
rect 225 29 226 30 
rect 225 30 226 31 
rect 225 31 226 32 
rect 225 32 226 33 
rect 225 33 226 34 
rect 225 34 226 35 
rect 225 35 226 36 
rect 225 36 226 37 
rect 225 37 226 38 
rect 225 38 226 39 
rect 225 39 226 40 
rect 225 40 226 41 
rect 225 41 226 42 
rect 225 42 226 43 
rect 225 43 226 44 
rect 225 44 226 45 
rect 225 45 226 46 
rect 225 46 226 47 
rect 225 47 226 48 
rect 225 48 226 49 
rect 225 49 226 50 
rect 225 50 226 51 
rect 225 52 226 53 
rect 225 54 226 55 
rect 225 56 226 57 
rect 225 82 226 83 
rect 225 84 226 85 
rect 225 117 226 118 
rect 225 118 226 119 
rect 225 119 226 120 
rect 225 120 226 121 
rect 225 152 226 153 
rect 225 165 226 166 
rect 225 168 226 169 
rect 225 183 226 184 
rect 225 186 226 187 
rect 225 187 226 188 
rect 225 188 226 189 
rect 225 189 226 190 
rect 225 190 226 191 
rect 225 191 226 192 
rect 225 193 226 194 
rect 225 200 226 201 
rect 225 216 226 217 
rect 225 223 226 224 
rect 225 224 226 225 
rect 225 230 226 231 
rect 225 231 226 232 
rect 225 232 226 233 
rect 225 233 226 234 
rect 225 242 226 243 
rect 225 248 226 249 
rect 225 257 226 258 
rect 225 261 226 262 
rect 225 262 226 263 
rect 225 263 226 264 
rect 225 264 226 265 
rect 225 265 226 266 
rect 225 266 226 267 
rect 225 267 226 268 
rect 225 268 226 269 
rect 225 269 226 270 
rect 225 270 226 271 
rect 225 271 226 272 
rect 225 272 226 273 
rect 225 273 226 274 
rect 225 274 226 275 
rect 225 275 226 276 
rect 225 276 226 277 
rect 225 277 226 278 
rect 225 278 226 279 
rect 225 279 226 280 
rect 225 280 226 281 
rect 225 281 226 282 
rect 225 282 226 283 
rect 225 283 226 284 
rect 225 284 226 285 
rect 225 285 226 286 
rect 225 286 226 287 
rect 225 287 226 288 
rect 225 288 226 289 
rect 226 52 227 53 
rect 226 54 227 55 
rect 226 56 227 57 
rect 226 65 227 66 
rect 226 66 227 67 
rect 226 67 227 68 
rect 226 68 227 69 
rect 226 69 227 70 
rect 226 70 227 71 
rect 226 71 227 72 
rect 226 72 227 73 
rect 226 73 227 74 
rect 226 82 227 83 
rect 226 84 227 85 
rect 226 148 227 149 
rect 226 152 227 153 
rect 226 165 227 166 
rect 226 168 227 169 
rect 226 183 227 184 
rect 226 191 227 192 
rect 226 193 227 194 
rect 226 200 227 201 
rect 226 216 227 217 
rect 226 223 227 224 
rect 226 248 227 249 
rect 226 257 227 258 
rect 226 293 227 294 
rect 226 294 227 295 
rect 226 295 227 296 
rect 226 296 227 297 
rect 226 297 227 298 
rect 226 298 227 299 
rect 226 299 227 300 
rect 226 300 227 301 
rect 226 301 227 302 
rect 226 302 227 303 
rect 226 303 227 304 
rect 226 304 227 305 
rect 226 305 227 306 
rect 226 306 227 307 
rect 227 52 228 53 
rect 227 54 228 55 
rect 227 56 228 57 
rect 227 82 228 83 
rect 227 84 228 85 
rect 227 148 228 149 
rect 227 152 228 153 
rect 227 165 228 166 
rect 227 168 228 169 
rect 227 183 228 184 
rect 227 186 228 187 
rect 227 187 228 188 
rect 227 188 228 189 
rect 227 189 228 190 
rect 227 191 228 192 
rect 227 193 228 194 
rect 227 200 228 201 
rect 227 216 228 217 
rect 227 223 228 224 
rect 227 225 228 226 
rect 227 226 228 227 
rect 227 227 228 228 
rect 227 228 228 229 
rect 227 229 228 230 
rect 227 230 228 231 
rect 227 231 228 232 
rect 227 232 228 233 
rect 227 233 228 234 
rect 227 234 228 235 
rect 227 235 228 236 
rect 227 236 228 237 
rect 227 237 228 238 
rect 227 238 228 239 
rect 227 239 228 240 
rect 227 240 228 241 
rect 227 241 228 242 
rect 227 242 228 243 
rect 227 243 228 244 
rect 227 244 228 245 
rect 227 245 228 246 
rect 227 246 228 247 
rect 227 248 228 249 
rect 227 257 228 258 
rect 228 52 229 53 
rect 228 54 229 55 
rect 228 56 229 57 
rect 228 65 229 66 
rect 228 66 229 67 
rect 228 67 229 68 
rect 228 68 229 69 
rect 228 69 229 70 
rect 228 70 229 71 
rect 228 71 229 72 
rect 228 72 229 73 
rect 228 73 229 74 
rect 228 82 229 83 
rect 228 84 229 85 
rect 228 111 229 112 
rect 228 112 229 113 
rect 228 113 229 114 
rect 228 114 229 115 
rect 228 148 229 149 
rect 228 152 229 153 
rect 228 165 229 166 
rect 228 168 229 169 
rect 228 183 229 184 
rect 228 191 229 192 
rect 228 193 229 194 
rect 228 200 229 201 
rect 228 216 229 217 
rect 228 223 229 224 
rect 228 225 229 226 
rect 228 247 229 248 
rect 228 248 229 249 
rect 228 257 229 258 
rect 229 54 230 55 
rect 229 56 230 57 
rect 229 82 230 83 
rect 229 84 230 85 
rect 229 111 230 112 
rect 229 114 230 115 
rect 229 115 230 116 
rect 229 148 230 149 
rect 229 152 230 153 
rect 229 165 230 166 
rect 229 168 230 169 
rect 229 183 230 184 
rect 229 191 230 192 
rect 229 193 230 194 
rect 229 200 230 201 
rect 229 216 230 217 
rect 229 223 230 224 
rect 229 227 230 228 
rect 229 228 230 229 
rect 229 229 230 230 
rect 229 230 230 231 
rect 229 231 230 232 
rect 229 232 230 233 
rect 229 233 230 234 
rect 229 234 230 235 
rect 229 235 230 236 
rect 229 236 230 237 
rect 229 237 230 238 
rect 229 238 230 239 
rect 229 239 230 240 
rect 229 240 230 241 
rect 229 241 230 242 
rect 229 242 230 243 
rect 229 243 230 244 
rect 229 246 230 247 
rect 229 247 230 248 
rect 229 257 230 258 
rect 230 54 231 55 
rect 230 56 231 57 
rect 230 82 231 83 
rect 230 84 231 85 
rect 230 94 231 95 
rect 230 95 231 96 
rect 230 96 231 97 
rect 230 97 231 98 
rect 230 98 231 99 
rect 230 99 231 100 
rect 230 113 231 114 
rect 230 115 231 116 
rect 230 118 231 119 
rect 230 119 231 120 
rect 230 148 231 149 
rect 230 152 231 153 
rect 230 165 231 166 
rect 230 168 231 169 
rect 230 184 231 185 
rect 230 185 231 186 
rect 230 186 231 187 
rect 230 193 231 194 
rect 230 200 231 201 
rect 230 216 231 217 
rect 230 223 231 224 
rect 230 245 231 246 
rect 230 246 231 247 
rect 230 257 231 258 
rect 231 54 232 55 
rect 231 56 232 57 
rect 231 82 232 83 
rect 231 84 232 85 
rect 231 93 232 94 
rect 231 94 232 95 
rect 231 113 232 114 
rect 231 115 232 116 
rect 231 118 232 119 
rect 231 148 232 149 
rect 231 152 232 153 
rect 231 165 232 166 
rect 231 168 232 169 
rect 231 184 232 185 
rect 231 193 232 194 
rect 231 200 232 201 
rect 231 216 232 217 
rect 231 223 232 224 
rect 231 242 232 243 
rect 231 243 232 244 
rect 231 244 232 245 
rect 231 245 232 246 
rect 231 257 232 258 
rect 232 54 233 55 
rect 232 56 233 57 
rect 232 82 233 83 
rect 232 84 233 85 
rect 232 96 233 97 
rect 232 97 233 98 
rect 232 98 233 99 
rect 232 99 233 100 
rect 232 100 233 101 
rect 232 101 233 102 
rect 232 113 233 114 
rect 232 115 233 116 
rect 232 118 233 119 
rect 232 148 233 149 
rect 232 152 233 153 
rect 232 165 233 166 
rect 232 168 233 169 
rect 232 184 233 185 
rect 232 193 233 194 
rect 232 200 233 201 
rect 232 216 233 217 
rect 232 242 233 243 
rect 232 257 233 258 
rect 233 54 234 55 
rect 233 56 234 57 
rect 233 82 234 83 
rect 233 84 234 85 
rect 233 101 234 102 
rect 233 113 234 114 
rect 233 115 234 116 
rect 233 118 234 119 
rect 233 148 234 149 
rect 233 152 234 153 
rect 233 165 234 166 
rect 233 168 234 169 
rect 233 184 234 185 
rect 233 193 234 194 
rect 233 200 234 201 
rect 233 216 234 217 
rect 233 242 234 243 
rect 233 257 234 258 
rect 234 54 235 55 
rect 234 56 235 57 
rect 234 82 235 83 
rect 234 84 235 85 
rect 234 101 235 102 
rect 234 113 235 114 
rect 234 118 235 119 
rect 234 148 235 149 
rect 234 152 235 153 
rect 234 165 235 166 
rect 234 168 235 169 
rect 234 184 235 185 
rect 234 193 235 194 
rect 234 200 235 201 
rect 234 216 235 217 
rect 234 242 235 243 
rect 234 257 235 258 
rect 235 54 236 55 
rect 235 56 236 57 
rect 235 82 236 83 
rect 235 84 236 85 
rect 235 101 236 102 
rect 235 113 236 114 
rect 235 118 236 119 
rect 235 148 236 149 
rect 235 152 236 153 
rect 235 165 236 166 
rect 235 168 236 169 
rect 235 184 236 185 
rect 235 193 236 194 
rect 235 200 236 201 
rect 235 216 236 217 
rect 235 242 236 243 
rect 235 257 236 258 
rect 236 54 237 55 
rect 236 56 237 57 
rect 236 82 237 83 
rect 236 84 237 85 
rect 236 101 237 102 
rect 236 113 237 114 
rect 236 118 237 119 
rect 236 148 237 149 
rect 236 152 237 153 
rect 236 165 237 166 
rect 236 168 237 169 
rect 236 184 237 185 
rect 236 193 237 194 
rect 236 200 237 201 
rect 236 216 237 217 
rect 236 242 237 243 
rect 236 257 237 258 
rect 237 54 238 55 
rect 237 56 238 57 
rect 237 82 238 83 
rect 237 84 238 85 
rect 237 101 238 102 
rect 237 113 238 114 
rect 237 118 238 119 
rect 237 148 238 149 
rect 237 152 238 153 
rect 237 165 238 166 
rect 237 168 238 169 
rect 237 184 238 185 
rect 237 193 238 194 
rect 237 200 238 201 
rect 237 216 238 217 
rect 237 242 238 243 
rect 237 257 238 258 
rect 238 54 239 55 
rect 238 56 239 57 
rect 238 82 239 83 
rect 238 84 239 85 
rect 238 101 239 102 
rect 238 113 239 114 
rect 238 118 239 119 
rect 238 148 239 149 
rect 238 152 239 153 
rect 238 165 239 166 
rect 238 168 239 169 
rect 238 184 239 185 
rect 238 193 239 194 
rect 238 200 239 201 
rect 238 216 239 217 
rect 238 242 239 243 
rect 238 244 239 245 
rect 238 257 239 258 
rect 239 2 240 3 
rect 239 3 240 4 
rect 239 4 240 5 
rect 239 5 240 6 
rect 239 6 240 7 
rect 239 7 240 8 
rect 239 8 240 9 
rect 239 37 240 38 
rect 239 54 240 55 
rect 239 56 240 57 
rect 239 82 240 83 
rect 239 84 240 85 
rect 239 88 240 89 
rect 239 99 240 100 
rect 239 101 240 102 
rect 239 113 240 114 
rect 239 118 240 119 
rect 239 148 240 149 
rect 239 152 240 153 
rect 239 165 240 166 
rect 239 168 240 169 
rect 239 184 240 185 
rect 239 193 240 194 
rect 239 200 240 201 
rect 239 216 240 217 
rect 239 241 240 242 
rect 239 242 240 243 
rect 239 244 240 245 
rect 239 257 240 258 
rect 240 8 241 9 
rect 240 9 241 10 
rect 240 37 241 38 
rect 240 40 241 41 
rect 240 54 241 55 
rect 240 56 241 57 
rect 240 66 241 67 
rect 240 68 241 69 
rect 240 82 241 83 
rect 240 84 241 85 
rect 240 88 241 89 
rect 240 97 241 98 
rect 240 99 241 100 
rect 240 101 241 102 
rect 240 113 241 114 
rect 240 118 241 119 
rect 240 120 241 121 
rect 240 121 241 122 
rect 240 148 241 149 
rect 240 152 241 153 
rect 240 165 241 166 
rect 240 168 241 169 
rect 240 184 241 185 
rect 240 185 241 186 
rect 240 193 241 194 
rect 240 200 241 201 
rect 240 209 241 210 
rect 240 211 241 212 
rect 240 216 241 217 
rect 240 217 241 218 
rect 240 241 241 242 
rect 240 244 241 245 
rect 240 257 241 258 
rect 240 304 241 305 
rect 240 305 241 306 
rect 240 306 241 307 
rect 241 9 242 10 
rect 241 10 242 11 
rect 241 37 242 38 
rect 241 40 242 41 
rect 241 54 242 55 
rect 241 56 242 57 
rect 241 66 242 67 
rect 241 68 242 69 
rect 241 82 242 83 
rect 241 84 242 85 
rect 241 88 242 89 
rect 241 97 242 98 
rect 241 99 242 100 
rect 241 101 242 102 
rect 241 113 242 114 
rect 241 118 242 119 
rect 241 121 242 122 
rect 241 122 242 123 
rect 241 123 242 124 
rect 241 124 242 125 
rect 241 125 242 126 
rect 241 126 242 127 
rect 241 127 242 128 
rect 241 128 242 129 
rect 241 129 242 130 
rect 241 148 242 149 
rect 241 152 242 153 
rect 241 165 242 166 
rect 241 168 242 169 
rect 241 185 242 186 
rect 241 186 242 187 
rect 241 193 242 194 
rect 241 200 242 201 
rect 241 209 242 210 
rect 241 211 242 212 
rect 241 217 242 218 
rect 241 218 242 219 
rect 241 219 242 220 
rect 241 220 242 221 
rect 241 221 242 222 
rect 241 222 242 223 
rect 241 223 242 224 
rect 241 224 242 225 
rect 241 225 242 226 
rect 241 226 242 227 
rect 241 227 242 228 
rect 241 228 242 229 
rect 241 229 242 230 
rect 241 230 242 231 
rect 241 231 242 232 
rect 241 232 242 233 
rect 241 233 242 234 
rect 241 234 242 235 
rect 241 241 242 242 
rect 241 244 242 245 
rect 241 257 242 258 
rect 241 261 242 262 
rect 241 262 242 263 
rect 241 263 242 264 
rect 241 264 242 265 
rect 241 303 242 304 
rect 241 304 242 305 
rect 242 37 243 38 
rect 242 40 243 41 
rect 242 54 243 55 
rect 242 56 243 57 
rect 242 66 243 67 
rect 242 68 243 69 
rect 242 82 243 83 
rect 242 84 243 85 
rect 242 88 243 89 
rect 242 97 243 98 
rect 242 99 243 100 
rect 242 101 243 102 
rect 242 113 243 114 
rect 242 118 243 119 
rect 242 129 243 130 
rect 242 148 243 149 
rect 242 152 243 153 
rect 242 165 243 166 
rect 242 168 243 169 
rect 242 193 243 194 
rect 242 200 243 201 
rect 242 209 243 210 
rect 242 211 243 212 
rect 242 241 243 242 
rect 242 244 243 245 
rect 242 257 243 258 
rect 243 37 244 38 
rect 243 40 244 41 
rect 243 54 244 55 
rect 243 56 244 57 
rect 243 66 244 67 
rect 243 68 244 69 
rect 243 82 244 83 
rect 243 84 244 85 
rect 243 88 244 89 
rect 243 97 244 98 
rect 243 99 244 100 
rect 243 101 244 102 
rect 243 113 244 114 
rect 243 118 244 119 
rect 243 129 244 130 
rect 243 148 244 149 
rect 243 152 244 153 
rect 243 165 244 166 
rect 243 168 244 169 
rect 243 193 244 194 
rect 243 200 244 201 
rect 243 209 244 210 
rect 243 211 244 212 
rect 243 241 244 242 
rect 243 244 244 245 
rect 243 248 244 249 
rect 243 257 244 258 
rect 244 31 245 32 
rect 244 32 245 33 
rect 244 33 245 34 
rect 244 34 245 35 
rect 244 37 245 38 
rect 244 54 245 55 
rect 244 56 245 57 
rect 244 68 245 69 
rect 244 82 245 83 
rect 244 84 245 85 
rect 244 88 245 89 
rect 244 99 245 100 
rect 244 113 245 114 
rect 244 118 245 119 
rect 244 129 245 130 
rect 244 148 245 149 
rect 244 152 245 153 
rect 244 165 245 166 
rect 244 168 245 169 
rect 244 193 245 194 
rect 244 200 245 201 
rect 244 209 245 210 
rect 244 211 245 212 
rect 244 228 245 229 
rect 244 229 245 230 
rect 244 230 245 231 
rect 244 231 245 232 
rect 244 232 245 233 
rect 244 233 245 234 
rect 244 241 245 242 
rect 244 244 245 245 
rect 244 248 245 249 
rect 245 31 246 32 
rect 245 37 246 38 
rect 245 40 246 41 
rect 245 41 246 42 
rect 245 42 246 43 
rect 245 43 246 44 
rect 245 54 246 55 
rect 245 56 246 57 
rect 245 68 246 69 
rect 245 82 246 83 
rect 245 84 246 85 
rect 245 88 246 89 
rect 245 89 246 90 
rect 245 90 246 91 
rect 245 91 246 92 
rect 245 92 246 93 
rect 245 93 246 94 
rect 245 94 246 95 
rect 245 95 246 96 
rect 245 99 246 100 
rect 245 113 246 114 
rect 245 118 246 119 
rect 245 129 246 130 
rect 245 148 246 149 
rect 245 152 246 153 
rect 245 165 246 166 
rect 245 168 246 169 
rect 245 193 246 194 
rect 245 200 246 201 
rect 245 209 246 210 
rect 245 211 246 212 
rect 245 241 246 242 
rect 245 244 246 245 
rect 245 248 246 249 
rect 245 256 246 257 
rect 245 257 246 258 
rect 245 258 246 259 
rect 245 259 246 260 
rect 245 260 246 261 
rect 245 261 246 262 
rect 245 262 246 263 
rect 245 263 246 264 
rect 245 264 246 265 
rect 245 265 246 266 
rect 245 266 246 267 
rect 245 267 246 268 
rect 245 268 246 269 
rect 245 269 246 270 
rect 245 270 246 271 
rect 245 271 246 272 
rect 245 272 246 273 
rect 245 273 246 274 
rect 245 274 246 275 
rect 245 275 246 276 
rect 245 276 246 277 
rect 245 277 246 278 
rect 245 278 246 279 
rect 245 279 246 280 
rect 245 280 246 281 
rect 245 281 246 282 
rect 246 37 247 38 
rect 246 54 247 55 
rect 246 56 247 57 
rect 246 68 247 69 
rect 246 82 247 83 
rect 246 84 247 85 
rect 246 99 247 100 
rect 246 113 247 114 
rect 246 118 247 119 
rect 246 129 247 130 
rect 246 148 247 149 
rect 246 152 247 153 
rect 246 165 247 166 
rect 246 193 247 194 
rect 246 200 247 201 
rect 246 209 247 210 
rect 246 211 247 212 
rect 246 241 247 242 
rect 246 244 247 245 
rect 246 248 247 249 
rect 247 32 248 33 
rect 247 37 248 38 
rect 247 54 248 55 
rect 247 56 248 57 
rect 247 65 248 66 
rect 247 68 248 69 
rect 247 82 248 83 
rect 247 84 248 85 
rect 247 87 248 88 
rect 247 88 248 89 
rect 247 89 248 90 
rect 247 90 248 91 
rect 247 91 248 92 
rect 247 92 248 93 
rect 247 93 248 94 
rect 247 94 248 95 
rect 247 95 248 96 
rect 247 96 248 97 
rect 247 97 248 98 
rect 247 98 248 99 
rect 247 99 248 100 
rect 247 101 248 102 
rect 247 113 248 114 
rect 247 118 248 119 
rect 247 129 248 130 
rect 247 148 248 149 
rect 247 152 248 153 
rect 247 165 248 166 
rect 247 193 248 194 
rect 247 200 248 201 
rect 247 211 248 212 
rect 247 241 248 242 
rect 247 244 248 245 
rect 247 248 248 249 
rect 248 32 249 33 
rect 248 37 249 38 
rect 248 40 249 41 
rect 248 41 249 42 
rect 248 42 249 43 
rect 248 43 249 44 
rect 248 54 249 55 
rect 248 56 249 57 
rect 248 65 249 66 
rect 248 68 249 69 
rect 248 82 249 83 
rect 248 84 249 85 
rect 248 85 249 86 
rect 248 100 249 101 
rect 248 101 249 102 
rect 248 113 249 114 
rect 248 118 249 119 
rect 248 129 249 130 
rect 248 148 249 149 
rect 248 152 249 153 
rect 248 165 249 166 
rect 248 180 249 181 
rect 248 182 249 183 
rect 248 183 249 184 
rect 248 184 249 185 
rect 248 185 249 186 
rect 248 193 249 194 
rect 248 200 249 201 
rect 248 211 249 212 
rect 248 228 249 229 
rect 248 229 249 230 
rect 248 230 249 231 
rect 248 231 249 232 
rect 248 232 249 233 
rect 248 233 249 234 
rect 248 241 249 242 
rect 248 244 249 245 
rect 248 248 249 249 
rect 248 256 249 257 
rect 248 257 249 258 
rect 248 258 249 259 
rect 248 259 249 260 
rect 248 260 249 261 
rect 248 261 249 262 
rect 248 262 249 263 
rect 248 263 249 264 
rect 248 264 249 265 
rect 248 265 249 266 
rect 248 266 249 267 
rect 248 267 249 268 
rect 248 268 249 269 
rect 248 269 249 270 
rect 248 270 249 271 
rect 248 271 249 272 
rect 248 272 249 273 
rect 248 273 249 274 
rect 248 274 249 275 
rect 248 275 249 276 
rect 248 276 249 277 
rect 248 277 249 278 
rect 248 278 249 279 
rect 248 279 249 280 
rect 248 280 249 281 
rect 248 281 249 282 
rect 249 32 250 33 
rect 249 33 250 34 
rect 249 37 250 38 
rect 249 54 250 55 
rect 249 56 250 57 
rect 249 65 250 66 
rect 249 68 250 69 
rect 249 82 250 83 
rect 249 85 250 86 
rect 249 86 250 87 
rect 249 87 250 88 
rect 249 88 250 89 
rect 249 97 250 98 
rect 249 98 250 99 
rect 249 99 250 100 
rect 249 100 250 101 
rect 249 113 250 114 
rect 249 118 250 119 
rect 249 129 250 130 
rect 249 148 250 149 
rect 249 152 250 153 
rect 249 165 250 166 
rect 249 180 250 181 
rect 249 181 250 182 
rect 249 193 250 194 
rect 249 200 250 201 
rect 249 211 250 212 
rect 249 241 250 242 
rect 249 244 250 245 
rect 249 248 250 249 
rect 250 33 251 34 
rect 250 37 251 38 
rect 250 54 251 55 
rect 250 56 251 57 
rect 250 65 251 66 
rect 250 68 251 69 
rect 250 82 251 83 
rect 250 88 251 89 
rect 250 97 251 98 
rect 250 113 251 114 
rect 250 118 251 119 
rect 250 129 251 130 
rect 250 148 251 149 
rect 250 152 251 153 
rect 250 165 251 166 
rect 250 181 251 182 
rect 250 182 251 183 
rect 250 183 251 184 
rect 250 184 251 185 
rect 250 193 251 194 
rect 250 200 251 201 
rect 250 211 251 212 
rect 250 241 251 242 
rect 250 244 251 245 
rect 250 248 251 249 
rect 251 54 252 55 
rect 251 65 252 66 
rect 251 68 252 69 
rect 251 88 252 89 
rect 251 97 252 98 
rect 251 113 252 114 
rect 251 118 252 119 
rect 251 129 252 130 
rect 251 152 252 153 
rect 251 165 252 166 
rect 251 184 252 185 
rect 251 193 252 194 
rect 251 200 252 201 
rect 251 211 252 212 
rect 251 241 252 242 
rect 251 244 252 245 
rect 251 248 252 249 
rect 252 65 253 66 
rect 252 68 253 69 
rect 252 88 253 89 
rect 252 97 253 98 
rect 252 113 253 114 
rect 252 118 253 119 
rect 252 129 253 130 
rect 252 152 253 153 
rect 252 184 253 185 
rect 252 193 253 194 
rect 252 200 253 201 
rect 252 211 253 212 
rect 252 241 253 242 
rect 252 244 253 245 
rect 252 248 253 249 
rect 253 65 254 66 
rect 253 68 254 69 
rect 253 88 254 89 
rect 253 97 254 98 
rect 253 113 254 114 
rect 253 118 254 119 
rect 253 129 254 130 
rect 253 152 254 153 
rect 253 184 254 185 
rect 253 193 254 194 
rect 253 200 254 201 
rect 253 211 254 212 
rect 253 241 254 242 
rect 253 244 254 245 
rect 253 248 254 249 
rect 254 65 255 66 
rect 254 68 255 69 
rect 254 88 255 89 
rect 254 97 255 98 
rect 254 113 255 114 
rect 254 118 255 119 
rect 254 129 255 130 
rect 254 152 255 153 
rect 254 184 255 185 
rect 254 193 255 194 
rect 254 200 255 201 
rect 254 211 255 212 
rect 254 226 255 227 
rect 254 241 255 242 
rect 254 244 255 245 
rect 254 248 255 249 
rect 255 65 256 66 
rect 255 68 256 69 
rect 255 88 256 89 
rect 255 97 256 98 
rect 255 113 256 114 
rect 255 118 256 119 
rect 255 129 256 130 
rect 255 152 256 153 
rect 255 184 256 185 
rect 255 193 256 194 
rect 255 200 256 201 
rect 255 211 256 212 
rect 255 226 256 227 
rect 255 241 256 242 
rect 255 244 256 245 
rect 255 248 256 249 
rect 256 65 257 66 
rect 256 68 257 69 
rect 256 88 257 89 
rect 256 89 257 90 
rect 256 96 257 97 
rect 256 97 257 98 
rect 256 113 257 114 
rect 256 118 257 119 
rect 256 121 257 122 
rect 256 129 257 130 
rect 256 152 257 153 
rect 256 184 257 185 
rect 256 185 257 186 
rect 256 192 257 193 
rect 256 193 257 194 
rect 256 198 257 199 
rect 256 200 257 201 
rect 256 208 257 209 
rect 256 209 257 210 
rect 256 211 257 212 
rect 256 226 257 227 
rect 256 240 257 241 
rect 256 241 257 242 
rect 256 244 257 245 
rect 256 248 257 249 
rect 256 249 257 250 
rect 257 7 258 8 
rect 257 8 258 9 
rect 257 9 258 10 
rect 257 10 258 11 
rect 257 65 258 66 
rect 257 68 258 69 
rect 257 83 258 84 
rect 257 84 258 85 
rect 257 85 258 86 
rect 257 86 258 87 
rect 257 89 258 90 
rect 257 90 258 91 
rect 257 91 258 92 
rect 257 92 258 93 
rect 257 93 258 94 
rect 257 94 258 95 
rect 257 96 258 97 
rect 257 113 258 114 
rect 257 115 258 116 
rect 257 118 258 119 
rect 257 121 258 122 
rect 257 122 258 123 
rect 257 123 258 124 
rect 257 129 258 130 
rect 257 152 258 153 
rect 257 185 258 186 
rect 257 186 258 187 
rect 257 187 258 188 
rect 257 188 258 189 
rect 257 189 258 190 
rect 257 190 258 191 
rect 257 191 258 192 
rect 257 198 258 199 
rect 257 200 258 201 
rect 257 202 258 203 
rect 257 203 258 204 
rect 257 204 258 205 
rect 257 205 258 206 
rect 257 206 258 207 
rect 257 207 258 208 
rect 257 208 258 209 
rect 257 211 258 212 
rect 257 226 258 227 
rect 257 229 258 230 
rect 257 230 258 231 
rect 257 231 258 232 
rect 257 232 258 233 
rect 257 233 258 234 
rect 257 234 258 235 
rect 257 235 258 236 
rect 257 236 258 237 
rect 257 237 258 238 
rect 257 239 258 240 
rect 257 240 258 241 
rect 257 244 258 245 
rect 257 249 258 250 
rect 257 250 258 251 
rect 257 251 258 252 
rect 257 252 258 253 
rect 257 253 258 254 
rect 257 254 258 255 
rect 257 255 258 256 
rect 257 256 258 257 
rect 257 257 258 258 
rect 257 258 258 259 
rect 257 259 258 260 
rect 257 260 258 261 
rect 257 261 258 262 
rect 257 262 258 263 
rect 257 263 258 264 
rect 257 264 258 265 
rect 258 65 259 66 
rect 258 68 259 69 
rect 258 94 259 95 
rect 258 96 259 97 
rect 258 113 259 114 
rect 258 115 259 116 
rect 258 118 259 119 
rect 258 129 259 130 
rect 258 152 259 153 
rect 258 191 259 192 
rect 258 192 259 193 
rect 258 193 259 194 
rect 258 194 259 195 
rect 258 195 259 196 
rect 258 196 259 197 
rect 258 198 259 199 
rect 258 200 259 201 
rect 258 202 259 203 
rect 258 211 259 212 
rect 258 226 259 227 
rect 258 239 259 240 
rect 258 244 259 245 
rect 259 37 260 38 
rect 259 38 260 39 
rect 259 39 260 40 
rect 259 40 260 41 
rect 259 41 260 42 
rect 259 42 260 43 
rect 259 43 260 44 
rect 259 44 260 45 
rect 259 45 260 46 
rect 259 65 260 66 
rect 259 68 260 69 
rect 259 94 260 95 
rect 259 96 260 97 
rect 259 113 260 114 
rect 259 115 260 116 
rect 259 118 260 119 
rect 259 129 260 130 
rect 259 143 260 144 
rect 259 144 260 145 
rect 259 145 260 146 
rect 259 146 260 147 
rect 259 152 260 153 
rect 259 163 260 164 
rect 259 164 260 165 
rect 259 165 260 166 
rect 259 166 260 167 
rect 259 197 260 198 
rect 259 198 260 199 
rect 259 200 260 201 
rect 259 202 260 203 
rect 259 211 260 212 
rect 259 226 260 227 
rect 259 230 260 231 
rect 259 231 260 232 
rect 259 232 260 233 
rect 259 233 260 234 
rect 259 234 260 235 
rect 259 235 260 236 
rect 259 236 260 237 
rect 259 237 260 238 
rect 259 238 260 239 
rect 259 239 260 240 
rect 260 65 261 66 
rect 260 68 261 69 
rect 260 95 261 96 
rect 260 96 261 97 
rect 260 113 261 114 
rect 260 115 261 116 
rect 260 118 261 119 
rect 260 152 261 153 
rect 260 185 261 186 
rect 260 186 261 187 
rect 260 187 261 188 
rect 260 188 261 189 
rect 260 189 261 190 
rect 260 190 261 191 
rect 260 191 261 192 
rect 260 192 261 193 
rect 260 193 261 194 
rect 260 194 261 195 
rect 260 195 261 196 
rect 260 196 261 197 
rect 260 197 261 198 
rect 260 200 261 201 
rect 260 202 261 203 
rect 261 36 262 37 
rect 261 37 262 38 
rect 261 38 262 39 
rect 261 39 262 40 
rect 261 40 262 41 
rect 261 41 262 42 
rect 261 42 262 43 
rect 261 43 262 44 
rect 261 44 262 45 
rect 261 45 262 46 
rect 261 46 262 47 
rect 261 65 262 66 
rect 261 68 262 69 
rect 261 83 262 84 
rect 261 84 262 85 
rect 261 85 262 86 
rect 261 86 262 87 
rect 261 87 262 88 
rect 261 88 262 89 
rect 261 89 262 90 
rect 261 90 262 91 
rect 261 91 262 92 
rect 261 92 262 93 
rect 261 93 262 94 
rect 261 94 262 95 
rect 261 95 262 96 
rect 261 114 262 115 
rect 261 115 262 116 
rect 261 118 262 119 
rect 261 121 262 122 
rect 261 122 262 123 
rect 261 123 262 124 
rect 261 124 262 125 
rect 261 125 262 126 
rect 261 126 262 127 
rect 261 127 262 128 
rect 261 128 262 129 
rect 261 129 262 130 
rect 261 130 262 131 
rect 261 131 262 132 
rect 261 132 262 133 
rect 261 133 262 134 
rect 261 134 262 135 
rect 261 135 262 136 
rect 261 136 262 137 
rect 261 137 262 138 
rect 261 138 262 139 
rect 261 139 262 140 
rect 261 140 262 141 
rect 261 141 262 142 
rect 261 142 262 143 
rect 261 143 262 144 
rect 261 144 262 145 
rect 261 145 262 146 
rect 261 146 262 147 
rect 261 152 262 153 
rect 261 200 262 201 
rect 261 202 262 203 
rect 262 65 263 66 
rect 262 68 263 69 
rect 262 112 263 113 
rect 262 113 263 114 
rect 262 114 263 115 
rect 262 118 263 119 
rect 262 152 263 153 
rect 262 163 263 164 
rect 262 164 263 165 
rect 262 165 263 166 
rect 262 166 263 167 
rect 262 167 263 168 
rect 262 168 263 169 
rect 262 169 263 170 
rect 262 170 263 171 
rect 262 171 263 172 
rect 262 172 263 173 
rect 262 173 263 174 
rect 262 174 263 175 
rect 262 175 263 176 
rect 262 176 263 177 
rect 262 177 263 178 
rect 262 178 263 179 
rect 262 179 263 180 
rect 262 180 263 181 
rect 262 181 263 182 
rect 262 182 263 183 
rect 262 183 263 184 
rect 262 184 263 185 
rect 262 185 263 186 
rect 262 186 263 187 
rect 262 187 263 188 
rect 262 188 263 189 
rect 262 189 263 190 
rect 262 190 263 191 
rect 262 191 263 192 
rect 262 192 263 193 
rect 262 193 263 194 
rect 262 194 263 195 
rect 262 195 263 196 
rect 262 200 263 201 
rect 262 202 263 203 
rect 263 68 264 69 
rect 263 95 264 96 
rect 263 96 264 97 
rect 263 97 264 98 
rect 263 98 264 99 
rect 263 118 264 119 
rect 263 144 264 145 
rect 263 145 264 146 
rect 263 146 264 147 
rect 263 147 264 148 
rect 263 152 264 153 
rect 263 200 264 201 
rect 263 202 264 203 
rect 264 68 265 69 
rect 264 84 265 85 
rect 264 85 265 86 
rect 264 86 265 87 
rect 264 87 265 88 
rect 264 118 265 119 
rect 264 152 265 153 
rect 264 185 265 186 
rect 264 186 265 187 
rect 264 187 265 188 
rect 264 188 265 189 
rect 264 189 265 190 
rect 264 190 265 191 
rect 264 191 265 192 
rect 264 192 265 193 
rect 264 193 265 194 
rect 264 194 265 195 
rect 264 195 265 196 
rect 264 201 265 202 
rect 264 202 265 203 
rect 264 229 265 230 
rect 264 230 265 231 
rect 264 231 265 232 
rect 264 232 265 233 
rect 264 233 265 234 
rect 264 234 265 235 
rect 264 235 265 236 
rect 264 236 265 237 
rect 264 237 265 238 
rect 264 238 265 239 
rect 264 239 265 240 
rect 264 240 265 241 
rect 264 241 265 242 
rect 264 242 265 243 
rect 264 243 265 244 
rect 264 244 265 245 
rect 264 245 265 246 
rect 265 68 266 69 
rect 265 118 266 119 
rect 265 152 266 153 
rect 265 200 266 201 
rect 265 201 266 202 
rect 266 68 267 69 
rect 266 115 267 116 
rect 266 118 267 119 
rect 266 152 267 153 
rect 266 200 267 201 
rect 267 68 268 69 
rect 267 115 268 116 
rect 267 118 268 119 
rect 267 152 268 153 
rect 267 200 268 201 
rect 268 68 269 69 
rect 268 115 269 116 
rect 268 117 269 118 
rect 268 118 269 119 
rect 268 152 269 153 
rect 268 200 269 201 
rect 269 68 270 69 
rect 269 115 270 116 
rect 269 117 270 118 
rect 269 152 270 153 
rect 269 200 270 201 
rect 270 68 271 69 
rect 270 115 271 116 
rect 270 117 271 118 
rect 270 152 271 153 
rect 270 200 271 201 
rect 271 68 272 69 
rect 271 115 272 116 
rect 271 117 272 118 
rect 271 152 272 153 
rect 271 200 272 201 
rect 272 68 273 69 
rect 272 85 273 86 
rect 272 104 273 105 
rect 272 115 273 116 
rect 272 117 273 118 
rect 272 119 273 120 
rect 272 152 273 153 
rect 272 198 273 199 
rect 272 200 273 201 
rect 272 240 273 241 
rect 272 241 273 242 
rect 272 243 273 244 
rect 272 246 273 247 
rect 272 258 273 259 
rect 273 68 274 69 
rect 273 85 274 86 
rect 273 104 274 105 
rect 273 115 274 116 
rect 273 117 274 118 
rect 273 119 274 120 
rect 273 152 274 153 
rect 273 192 274 193 
rect 273 193 274 194 
rect 273 194 274 195 
rect 273 195 274 196 
rect 273 198 274 199 
rect 273 200 274 201 
rect 273 232 274 233 
rect 273 233 274 234 
rect 273 234 274 235 
rect 273 235 274 236 
rect 273 236 274 237 
rect 273 237 274 238 
rect 273 238 274 239 
rect 273 239 274 240 
rect 273 240 274 241 
rect 273 243 274 244 
rect 273 246 274 247 
rect 273 258 274 259 
rect 273 261 274 262 
rect 273 262 274 263 
rect 273 263 274 264 
rect 273 264 274 265 
rect 274 68 275 69 
rect 274 85 275 86 
rect 274 104 275 105 
rect 274 115 275 116 
rect 274 117 275 118 
rect 274 119 275 120 
rect 274 152 275 153 
rect 274 197 275 198 
rect 274 198 275 199 
rect 274 200 275 201 
rect 274 232 275 233 
rect 274 243 275 244 
rect 274 246 275 247 
rect 274 258 275 259 
rect 275 68 276 69 
rect 275 85 276 86 
rect 275 104 276 105 
rect 275 115 276 116 
rect 275 117 276 118 
rect 275 119 276 120 
rect 275 152 276 153 
rect 275 183 276 184 
rect 275 184 276 185 
rect 275 185 276 186 
rect 275 186 276 187 
rect 275 187 276 188 
rect 275 188 276 189 
rect 275 189 276 190 
rect 275 190 276 191 
rect 275 191 276 192 
rect 275 192 276 193 
rect 275 193 276 194 
rect 275 194 276 195 
rect 275 195 276 196 
rect 275 196 276 197 
rect 275 197 276 198 
rect 275 199 276 200 
rect 275 200 276 201 
rect 275 232 276 233 
rect 275 243 276 244 
rect 275 246 276 247 
rect 275 258 276 259 
rect 276 115 277 116 
rect 276 117 277 118 
rect 276 119 277 120 
rect 276 152 277 153 
rect 276 164 277 165 
rect 276 165 277 166 
rect 276 166 277 167 
rect 276 167 277 168 
rect 276 168 277 169 
rect 276 169 277 170 
rect 276 170 277 171 
rect 276 171 277 172 
rect 276 172 277 173 
rect 276 173 277 174 
rect 276 174 277 175 
rect 276 175 277 176 
rect 276 176 277 177 
rect 276 198 277 199 
rect 276 199 277 200 
rect 276 232 277 233 
rect 276 243 277 244 
rect 276 246 277 247 
rect 277 115 278 116 
rect 277 117 278 118 
rect 277 119 278 120 
rect 277 152 278 153 
rect 277 162 278 163 
rect 277 163 278 164 
rect 277 192 278 193 
rect 277 193 278 194 
rect 277 194 278 195 
rect 277 195 278 196 
rect 277 196 278 197 
rect 277 197 278 198 
rect 277 198 278 199 
rect 277 232 278 233 
rect 277 243 278 244 
rect 277 246 278 247 
rect 277 257 278 258 
rect 277 258 278 259 
rect 277 259 278 260 
rect 277 260 278 261 
rect 277 261 278 262 
rect 277 262 278 263 
rect 277 263 278 264 
rect 277 264 278 265 
rect 277 265 278 266 
rect 277 266 278 267 
rect 277 267 278 268 
rect 277 268 278 269 
rect 277 269 278 270 
rect 277 270 278 271 
rect 277 271 278 272 
rect 277 272 278 273 
rect 277 273 278 274 
rect 277 274 278 275 
rect 277 275 278 276 
rect 277 276 278 277 
rect 277 277 278 278 
rect 277 278 278 279 
rect 277 279 278 280 
rect 277 280 278 281 
rect 277 281 278 282 
rect 278 115 279 116 
rect 278 117 279 118 
rect 278 119 279 120 
rect 278 152 279 153 
rect 278 163 279 164 
rect 278 164 279 165 
rect 278 165 279 166 
rect 278 166 279 167 
rect 278 167 279 168 
rect 278 168 279 169 
rect 278 169 279 170 
rect 278 170 279 171 
rect 278 171 279 172 
rect 278 172 279 173 
rect 278 173 279 174 
rect 278 174 279 175 
rect 278 175 279 176 
rect 278 199 279 200 
rect 278 232 279 233 
rect 278 243 279 244 
rect 278 246 279 247 
rect 279 115 280 116 
rect 279 117 280 118 
rect 279 119 280 120 
rect 279 152 280 153 
rect 279 175 280 176 
rect 279 176 280 177 
rect 279 177 280 178 
rect 279 178 280 179 
rect 279 179 280 180 
rect 279 180 280 181 
rect 279 181 280 182 
rect 279 182 280 183 
rect 279 183 280 184 
rect 279 184 280 185 
rect 279 185 280 186 
rect 279 186 280 187 
rect 279 187 280 188 
rect 279 188 280 189 
rect 279 189 280 190 
rect 279 190 280 191 
rect 279 191 280 192 
rect 279 192 280 193 
rect 279 193 280 194 
rect 279 194 280 195 
rect 279 195 280 196 
rect 279 196 280 197 
rect 279 197 280 198 
rect 279 198 280 199 
rect 279 199 280 200 
rect 279 232 280 233 
rect 279 243 280 244 
rect 279 246 280 247 
rect 280 119 281 120 
rect 280 152 281 153 
rect 280 232 281 233 
rect 280 243 281 244 
rect 280 246 281 247 
rect 280 248 281 249 
rect 280 249 281 250 
rect 280 250 281 251 
rect 280 251 281 252 
rect 280 252 281 253 
rect 280 253 281 254 
rect 280 254 281 255 
rect 280 255 281 256 
rect 280 256 281 257 
rect 280 257 281 258 
rect 280 258 281 259 
rect 280 259 281 260 
rect 280 260 281 261 
rect 280 261 281 262 
rect 280 262 281 263 
rect 280 263 281 264 
rect 280 264 281 265 
rect 280 265 281 266 
rect 280 266 281 267 
rect 280 267 281 268 
rect 280 268 281 269 
rect 280 269 281 270 
rect 280 270 281 271 
rect 280 271 281 272 
rect 280 272 281 273 
rect 280 273 281 274 
rect 280 274 281 275 
rect 280 275 281 276 
rect 280 276 281 277 
rect 281 119 282 120 
rect 281 232 282 233 
rect 281 243 282 244 
rect 281 246 282 247 
rect 281 248 282 249 
rect 282 119 283 120 
rect 282 232 283 233 
rect 282 243 283 244 
rect 282 246 283 247 
rect 282 248 283 249 
rect 283 119 284 120 
rect 283 243 284 244 
rect 283 246 284 247 
rect 283 247 284 248 
rect 284 119 285 120 
rect 284 243 285 244 
rect 284 247 285 248 
rect 285 119 286 120 
rect 285 225 286 226 
rect 285 243 286 244 
rect 286 119 287 120 
rect 286 225 287 226 
rect 286 243 287 244 
rect 287 119 288 120 
rect 287 166 288 167 
rect 287 225 288 226 
rect 287 243 288 244 
rect 287 259 288 260 
rect 287 262 288 263 
rect 288 119 289 120 
rect 288 166 289 167 
rect 288 168 289 169 
rect 288 225 289 226 
rect 288 243 289 244 
rect 288 259 289 260 
rect 288 262 289 263 
rect 289 119 290 120 
rect 289 120 290 121 
rect 289 121 290 122 
rect 289 122 290 123 
rect 289 123 290 124 
rect 289 166 290 167 
rect 289 168 290 169 
rect 289 225 290 226 
rect 289 243 290 244 
rect 289 259 290 260 
rect 289 262 290 263 
rect 289 264 290 265 
rect 289 265 290 266 
rect 289 266 290 267 
rect 289 267 290 268 
rect 289 268 290 269 
rect 289 269 290 270 
rect 289 270 290 271 
rect 289 271 290 272 
rect 289 272 290 273 
rect 289 273 290 274 
rect 289 274 290 275 
rect 289 275 290 276 
rect 289 276 290 277 
rect 290 166 291 167 
rect 290 168 291 169 
rect 290 225 291 226 
rect 290 243 291 244 
rect 290 259 291 260 
rect 290 262 291 263 
rect 290 264 291 265 
rect 291 41 292 42 
rect 291 42 292 43 
rect 291 43 292 44 
rect 291 44 292 45 
rect 291 166 292 167 
rect 291 168 292 169 
rect 291 225 292 226 
rect 291 243 292 244 
rect 291 258 292 259 
rect 291 259 292 260 
rect 291 263 292 264 
rect 291 264 292 265 
rect 292 166 293 167 
rect 292 168 293 169 
rect 292 225 293 226 
rect 292 243 293 244 
rect 292 258 293 259 
rect 292 260 293 261 
rect 292 261 293 262 
rect 292 262 293 263 
rect 292 263 293 264 
rect 292 274 293 275 
rect 293 156 294 157 
rect 293 157 294 158 
rect 293 158 294 159 
rect 293 159 294 160 
rect 293 166 294 167 
rect 293 168 294 169 
rect 293 170 294 171 
rect 293 171 294 172 
rect 293 172 294 173 
rect 293 173 294 174 
rect 293 174 294 175 
rect 293 175 294 176 
rect 293 176 294 177 
rect 293 177 294 178 
rect 293 225 294 226 
rect 293 243 294 244 
rect 293 258 294 259 
rect 293 268 294 269 
rect 293 269 294 270 
rect 293 270 294 271 
rect 293 271 294 272 
rect 293 274 294 275 
rect 294 156 295 157 
rect 294 166 295 167 
rect 294 167 295 168 
rect 294 169 295 170 
rect 294 170 295 171 
rect 294 243 295 244 
rect 294 258 295 259 
rect 294 273 295 274 
rect 294 274 295 275 
rect 295 156 296 157 
rect 295 167 296 168 
rect 295 168 296 169 
rect 295 169 296 170 
rect 295 243 296 244 
rect 295 258 296 259 
rect 295 268 296 269 
rect 295 269 296 270 
rect 295 270 296 271 
rect 295 271 296 272 
rect 295 272 296 273 
rect 295 273 296 274 
rect 296 38 297 39 
rect 296 243 297 244 
rect 296 258 297 259 
rect 297 38 298 39 
rect 297 243 298 244 
rect 297 258 298 259 
rect 297 259 298 260 
rect 298 38 299 39 
rect 298 243 299 244 
rect 298 259 299 260 
rect 299 38 300 39 
rect 299 243 300 244 
rect 299 259 300 260 
rect 300 243 301 244 
rect 301 243 302 244 
rect 302 243 303 244 
rect 303 243 304 244 
rect 304 243 305 244 
rect 305 243 306 244 
rect 306 243 307 244 
rect 307 243 308 244 
<< m2contact >>
rect 2 134 3 135 
rect 17 218 18 219 
rect 17 288 18 289 
rect 19 165 20 166 
rect 20 168 21 169 
rect 20 219 21 220 
rect 22 161 23 162 
rect 24 138 25 139 
rect 24 170 25 171 
rect 24 205 25 206 
rect 26 101 27 102 
rect 30 123 31 124 
rect 36 157 37 158 
rect 36 165 37 166 
rect 38 84 39 85 
rect 38 134 39 135 
rect 38 165 39 166 
rect 39 193 40 194 
rect 40 145 41 146 
rect 40 161 41 162 
rect 42 104 43 105 
rect 45 56 46 57 
rect 47 116 48 117 
rect 49 101 50 102 
rect 49 161 50 162 
rect 49 230 50 231 
rect 50 80 51 81 
rect 50 215 51 216 
rect 51 49 52 50 
rect 51 101 52 102 
rect 51 161 52 162 
rect 51 234 52 235 
rect 52 80 53 81 
rect 53 195 54 196 
rect 54 129 55 130 
rect 54 246 55 247 
rect 56 161 57 162 
rect 56 234 57 235 
rect 56 271 57 272 
rect 56 309 57 310 
rect 63 225 64 226 
rect 65 84 66 85 
rect 66 245 67 246 
rect 67 168 68 169 
rect 67 197 68 198 
rect 67 212 68 213 
rect 68 88 69 89 
rect 69 218 70 219 
rect 70 257 71 258 
rect 70 276 71 277 
rect 72 38 73 39 
rect 74 56 75 57 
rect 74 65 75 66 
rect 74 70 75 71 
rect 74 72 75 73 
rect 74 103 75 104 
rect 74 131 75 132 
rect 74 133 75 134 
rect 74 136 75 137 
rect 74 152 75 153 
rect 74 165 75 166 
rect 74 210 75 211 
rect 74 232 75 233 
rect 74 241 75 242 
rect 74 245 75 246 
rect 76 100 77 101 
rect 81 21 82 22 
rect 81 127 82 128 
rect 81 231 82 232 
rect 81 309 82 310 
rect 82 71 83 72 
rect 83 138 84 139 
rect 83 167 84 168 
rect 83 200 84 201 
rect 83 278 84 279 
rect 85 100 86 101 
rect 86 145 87 146 
rect 88 134 89 135 
rect 95 84 96 85 
rect 95 100 96 101 
rect 96 20 97 21 
rect 96 69 97 70 
rect 96 249 97 250 
rect 97 218 98 219 
rect 97 303 98 304 
rect 98 189 99 190 
rect 98 201 99 202 
rect 99 86 100 87 
rect 99 98 100 99 
rect 99 102 100 103 
rect 102 133 103 134 
rect 102 218 103 219 
rect 104 218 105 219 
rect 106 195 107 196 
rect 113 71 114 72 
rect 113 134 114 135 
rect 113 245 114 246 
rect 115 16 116 17 
rect 115 84 116 85 
rect 115 132 116 133 
rect 115 249 116 250 
rect 115 261 116 262 
rect 115 263 116 264 
rect 117 36 118 37 
rect 117 181 118 182 
rect 117 226 118 227 
rect 119 278 120 279 
rect 121 48 122 49 
rect 121 69 122 70 
rect 121 195 122 196 
rect 121 228 122 229 
rect 121 241 122 242 
rect 121 243 122 244 
rect 125 166 126 167 
rect 129 25 130 26 
rect 130 140 131 141 
rect 132 48 133 49 
rect 132 86 133 87 
rect 132 97 133 98 
rect 133 252 134 253 
rect 134 69 135 70 
rect 134 118 135 119 
rect 134 165 135 166 
rect 134 182 135 183 
rect 134 212 135 213 
rect 134 230 135 231 
rect 138 116 139 117 
rect 138 134 139 135 
rect 138 136 139 137 
rect 138 145 139 146 
rect 138 148 139 149 
rect 138 161 139 162 
rect 138 232 139 233 
rect 138 248 139 249 
rect 138 259 139 260 
rect 138 280 139 281 
rect 140 163 141 164 
rect 140 228 141 229 
rect 140 243 141 244 
rect 140 278 141 279 
rect 140 289 141 290 
rect 140 291 141 292 
rect 142 278 143 279 
rect 145 18 146 19 
rect 145 171 146 172 
rect 145 242 146 243 
rect 145 295 146 296 
rect 146 184 147 185 
rect 147 56 148 57 
rect 147 104 148 105 
rect 147 165 148 166 
rect 147 167 148 168 
rect 147 238 148 239 
rect 149 157 150 158 
rect 150 197 151 198 
rect 152 186 153 187 
rect 152 271 153 272 
rect 154 52 155 53 
rect 154 65 155 66 
rect 154 97 155 98 
rect 154 132 155 133 
rect 154 216 155 217 
rect 154 246 155 247 
rect 154 248 155 249 
rect 154 259 155 260 
rect 156 52 157 53 
rect 160 48 161 49 
rect 161 18 162 19 
rect 161 116 162 117 
rect 161 138 162 139 
rect 161 246 162 247 
rect 163 16 164 17 
rect 163 138 164 139 
rect 163 230 164 231 
rect 163 259 164 260 
rect 164 95 165 96 
rect 164 165 165 166 
rect 165 116 166 117 
rect 165 195 166 196 
rect 165 201 166 202 
rect 165 214 166 215 
rect 165 282 166 283 
rect 166 102 167 103 
rect 166 163 167 164 
rect 170 65 171 66 
rect 175 34 176 35 
rect 175 120 176 121 
rect 176 25 177 26 
rect 176 48 177 49 
rect 176 73 177 74 
rect 177 95 178 96 
rect 177 282 178 283 
rect 179 65 180 66 
rect 179 76 180 77 
rect 179 195 180 196 
rect 182 163 183 164 
rect 182 234 183 235 
rect 182 262 183 263 
rect 183 52 184 53 
rect 184 120 185 121 
rect 184 179 185 180 
rect 184 243 185 244 
rect 184 266 185 267 
rect 185 57 186 58 
rect 185 256 186 257 
rect 192 17 193 18 
rect 192 25 193 26 
rect 192 34 193 35 
rect 192 73 193 74 
rect 193 42 194 43 
rect 193 68 194 69 
rect 193 92 194 93 
rect 193 163 194 164 
rect 193 230 194 231 
rect 193 275 194 276 
rect 193 303 194 304 
rect 195 99 196 100 
rect 195 184 196 185 
rect 195 271 196 272 
rect 195 289 196 290 
rect 196 226 197 227 
rect 197 81 198 82 
rect 197 99 198 100 
rect 197 262 198 263 
rect 198 244 199 245 
rect 198 246 199 247 
rect 198 258 199 259 
rect 199 102 200 103 
rect 203 264 204 265 
rect 210 271 211 272 
rect 210 303 211 304 
rect 212 278 213 279 
rect 214 150 215 151 
rect 214 161 215 162 
rect 214 163 215 164 
rect 214 243 215 244 
rect 214 253 215 254 
rect 214 309 215 310 
rect 216 120 217 121 
rect 216 197 217 198 
rect 218 295 219 296 
rect 220 291 221 292 
rect 224 56 225 57 
rect 225 50 226 51 
rect 225 120 226 121 
rect 225 230 226 231 
rect 225 242 226 243 
rect 226 73 227 74 
rect 226 293 227 294 
rect 227 189 228 190 
rect 227 246 228 247 
rect 228 52 229 53 
rect 228 73 229 74 
rect 229 183 230 184 
rect 229 191 230 192 
rect 229 227 230 228 
rect 230 99 231 100 
rect 231 223 232 224 
rect 233 115 234 116 
rect 239 88 240 89 
rect 239 99 240 100 
rect 241 10 242 11 
rect 241 186 242 187 
rect 241 234 242 235 
rect 241 264 242 265 
rect 241 303 242 304 
rect 243 40 244 41 
rect 243 66 244 67 
rect 243 97 244 98 
rect 243 101 244 102 
rect 243 257 244 258 
rect 244 34 245 35 
rect 244 228 245 229 
rect 245 43 246 44 
rect 245 168 246 169 
rect 245 256 246 257 
rect 246 209 247 210 
rect 248 43 249 44 
rect 248 182 249 183 
rect 248 228 249 229 
rect 248 256 249 257 
rect 250 33 251 34 
rect 250 37 251 38 
rect 250 82 251 83 
rect 250 148 251 149 
rect 251 54 252 55 
rect 251 165 252 166 
rect 256 121 257 122 
rect 256 192 257 193 
rect 257 10 258 11 
rect 257 83 258 84 
rect 257 237 258 238 
rect 257 264 258 265 
rect 258 196 259 197 
rect 258 244 259 245 
rect 259 45 260 46 
rect 259 94 260 95 
rect 259 129 260 130 
rect 259 143 260 144 
rect 259 163 260 164 
rect 259 211 260 212 
rect 259 226 260 227 
rect 259 230 260 231 
rect 260 113 261 114 
rect 260 185 261 186 
rect 261 36 262 37 
rect 261 83 262 84 
rect 261 121 262 122 
rect 262 65 263 66 
rect 262 112 263 113 
rect 262 163 263 164 
rect 263 95 264 96 
rect 263 147 264 148 
rect 263 200 264 201 
rect 264 87 265 88 
rect 264 185 265 186 
rect 264 245 265 246 
rect 273 192 274 193 
rect 273 264 274 265 
rect 275 68 276 69 
rect 275 85 276 86 
rect 275 104 276 105 
rect 275 183 276 184 
rect 275 258 276 259 
rect 276 164 277 165 
rect 277 192 278 193 
rect 277 281 278 282 
rect 278 199 279 200 
rect 279 115 280 116 
rect 279 117 280 118 
rect 280 152 281 153 
rect 282 232 283 233 
rect 282 248 283 249 
rect 284 247 285 248 
rect 287 166 288 167 
rect 289 123 290 124 
rect 290 262 291 263 
rect 291 41 292 42 
rect 292 260 293 261 
rect 293 168 294 169 
rect 293 225 294 226 
rect 293 268 294 269 
rect 295 156 296 157 
rect 295 268 296 269 
rect 299 38 300 39 
rect 299 259 300 260 
rect 307 243 308 244 
rect 8 205 9 206 
rect 17 214 18 215 
rect 17 284 18 285 
rect 18 172 19 173 
rect 19 161 20 162 
rect 22 97 23 98 
rect 22 165 23 166 
rect 24 168 25 169 
rect 24 199 25 200 
rect 24 219 25 220 
rect 25 132 26 133 
rect 26 97 27 98 
rect 31 161 32 162 
rect 34 67 35 68 
rect 34 99 35 100 
rect 34 130 35 131 
rect 34 134 35 135 
rect 34 136 35 137 
rect 34 145 35 146 
rect 35 200 36 201 
rect 38 80 39 81 
rect 38 132 39 133 
rect 38 161 39 162 
rect 40 165 41 166 
rect 42 97 43 98 
rect 42 113 43 114 
rect 46 145 47 146 
rect 46 212 47 213 
rect 46 215 47 216 
rect 46 228 47 229 
rect 47 49 48 50 
rect 47 54 48 55 
rect 47 193 48 194 
rect 47 197 48 198 
rect 48 97 49 98 
rect 49 165 50 166 
rect 49 246 50 247 
rect 50 84 51 85 
rect 51 105 52 106 
rect 51 165 52 166 
rect 53 152 54 153 
rect 54 165 55 166 
rect 54 230 55 231 
rect 56 103 57 104 
rect 56 165 57 166 
rect 56 261 57 262 
rect 56 275 57 276 
rect 56 302 57 303 
rect 57 57 58 58 
rect 57 80 58 81 
rect 61 51 62 52 
rect 63 98 64 99 
rect 63 163 64 164 
rect 65 73 66 74 
rect 66 239 67 240 
rect 67 210 68 211 
rect 68 65 69 66 
rect 68 75 69 76 
rect 68 131 69 132 
rect 68 259 69 260 
rect 70 165 71 166 
rect 70 216 71 217 
rect 70 227 71 228 
rect 70 241 71 242 
rect 70 243 71 244 
rect 70 245 71 246 
rect 72 27 73 28 
rect 74 129 75 130 
rect 74 148 75 149 
rect 74 257 75 258 
rect 76 225 77 226 
rect 80 38 81 39 
rect 81 25 82 26 
rect 81 237 82 238 
rect 81 302 82 303 
rect 82 75 83 76 
rect 82 229 83 230 
rect 83 134 84 135 
rect 83 282 84 283 
rect 84 88 85 89 
rect 85 110 86 111 
rect 86 51 87 52 
rect 86 69 87 70 
rect 87 40 88 41 
rect 88 102 89 103 
rect 88 131 89 132 
rect 88 138 89 139 
rect 89 224 90 225 
rect 90 195 91 196 
rect 92 65 93 66 
rect 95 88 96 89 
rect 95 263 96 264 
rect 96 245 97 246 
rect 97 143 98 144 
rect 97 159 98 160 
rect 97 307 98 308 
rect 99 119 100 120 
rect 100 84 101 85 
rect 100 177 101 178 
rect 100 184 101 185 
rect 100 195 101 196 
rect 100 199 101 200 
rect 102 116 103 117 
rect 104 119 105 120 
rect 104 212 105 213 
rect 110 149 111 150 
rect 111 69 112 70 
rect 111 181 112 182 
rect 111 241 112 242 
rect 113 36 114 37 
rect 113 38 114 39 
rect 113 50 114 51 
rect 113 52 114 53 
rect 113 56 114 57 
rect 113 138 114 139 
rect 113 224 114 225 
rect 113 249 114 250 
rect 113 282 114 283 
rect 115 25 116 26 
rect 115 86 116 87 
rect 115 138 116 139 
rect 115 245 116 246 
rect 117 97 118 98 
rect 117 102 118 103 
rect 117 104 118 105 
rect 117 195 118 196 
rect 117 276 118 277 
rect 119 282 120 283 
rect 121 181 122 182 
rect 121 197 122 198 
rect 124 293 125 294 
rect 127 257 128 258 
rect 127 261 128 262 
rect 128 48 129 49 
rect 128 73 129 74 
rect 129 15 130 16 
rect 129 239 130 240 
rect 130 111 131 112 
rect 131 148 132 149 
rect 132 116 133 117 
rect 132 138 133 139 
rect 132 221 133 222 
rect 132 250 133 251 
rect 134 84 135 85 
rect 134 97 135 98 
rect 134 111 135 112 
rect 134 132 135 133 
rect 134 136 135 137 
rect 134 152 135 153 
rect 134 161 135 162 
rect 134 195 135 196 
rect 134 232 135 233 
rect 134 241 135 242 
rect 134 246 135 247 
rect 134 248 135 249 
rect 134 259 135 260 
rect 134 280 135 281 
rect 135 289 136 290 
rect 136 291 137 292 
rect 138 118 139 119 
rect 140 230 141 231 
rect 142 161 143 162 
rect 143 166 144 167 
rect 145 222 146 223 
rect 145 286 146 287 
rect 146 248 147 249 
rect 146 259 147 260 
rect 146 263 147 264 
rect 147 157 148 158 
rect 147 210 148 211 
rect 147 244 148 245 
rect 148 57 149 58 
rect 149 171 150 172 
rect 150 189 151 190 
rect 152 268 153 269 
rect 153 25 154 26 
rect 153 134 154 135 
rect 154 69 155 70 
rect 154 71 155 72 
rect 154 280 155 281 
rect 158 104 159 105 
rect 160 165 161 166 
rect 161 120 162 121 
rect 161 201 162 202 
rect 163 25 164 26 
rect 163 93 164 94 
rect 163 251 164 252 
rect 164 99 165 100 
rect 165 154 166 155 
rect 165 197 166 198 
rect 165 270 166 271 
rect 166 65 167 66 
rect 166 169 167 170 
rect 168 143 169 144 
rect 168 219 169 220 
rect 168 282 169 283 
rect 175 40 176 41 
rect 175 113 176 114 
rect 175 197 176 198 
rect 176 69 177 70 
rect 177 57 178 58 
rect 177 169 178 170 
rect 177 261 178 262 
rect 178 210 179 211 
rect 179 69 180 70 
rect 179 251 180 252 
rect 182 83 183 84 
rect 182 85 183 86 
rect 182 274 183 275 
rect 183 34 184 35 
rect 184 15 185 16 
rect 184 31 185 32 
rect 184 95 185 96 
rect 184 113 185 114 
rect 184 140 185 141 
rect 184 227 185 228 
rect 184 258 185 259 
rect 186 230 187 231 
rect 191 21 192 22 
rect 191 163 192 164 
rect 191 277 192 278 
rect 191 279 192 280 
rect 191 291 192 292 
rect 191 293 192 294 
rect 192 38 193 39 
rect 192 69 193 70 
rect 192 262 193 263 
rect 193 64 194 65 
rect 193 120 194 121 
rect 193 151 194 152 
rect 193 173 194 174 
rect 193 234 194 235 
rect 193 271 194 272 
rect 193 307 194 308 
rect 194 228 195 229 
rect 194 260 195 261 
rect 195 92 196 93 
rect 196 234 197 235 
rect 198 161 199 162 
rect 206 275 207 276 
rect 208 165 209 166 
rect 208 184 209 185 
rect 210 307 211 308 
rect 212 243 213 244 
rect 212 253 213 254 
rect 214 114 215 115 
rect 214 230 215 231 
rect 214 266 215 267 
rect 216 114 217 115 
rect 216 239 217 240 
rect 216 255 217 256 
rect 221 84 222 85 
rect 223 168 224 169 
rect 223 200 224 201 
rect 224 52 225 53 
rect 224 54 225 55 
rect 225 28 226 29 
rect 225 116 226 117 
rect 225 148 226 149 
rect 225 185 226 186 
rect 225 234 226 235 
rect 225 260 226 261 
rect 226 64 227 65 
rect 226 307 227 308 
rect 227 185 228 186 
rect 228 64 229 65 
rect 229 110 230 111 
rect 229 225 230 226 
rect 229 244 230 245 
rect 230 112 231 113 
rect 230 120 231 121 
rect 230 187 231 188 
rect 232 93 233 94 
rect 232 95 233 96 
rect 237 244 238 245 
rect 239 1 240 2 
rect 239 38 240 39 
rect 239 40 240 41 
rect 239 66 240 67 
rect 239 68 240 69 
rect 239 97 240 98 
rect 239 120 240 121 
rect 239 209 240 210 
rect 239 211 240 212 
rect 240 307 241 308 
rect 241 260 242 261 
rect 242 248 243 249 
rect 244 234 245 235 
rect 245 30 246 31 
rect 245 39 246 40 
rect 245 96 246 97 
rect 245 282 246 283 
rect 246 32 247 33 
rect 246 65 247 66 
rect 246 101 247 102 
rect 247 86 248 87 
rect 247 180 248 181 
rect 248 39 249 40 
rect 248 186 249 187 
rect 248 234 249 235 
rect 248 282 249 283 
rect 251 56 252 57 
rect 253 226 254 227 
rect 255 198 256 199 
rect 255 209 256 210 
rect 256 115 257 116 
rect 257 6 258 7 
rect 257 87 258 88 
rect 257 124 258 125 
rect 257 228 258 229 
rect 259 36 260 37 
rect 259 147 260 148 
rect 259 167 260 168 
rect 261 47 262 48 
rect 261 147 262 148 
rect 262 196 263 197 
rect 263 99 264 100 
rect 263 143 264 144 
rect 264 83 265 84 
rect 264 196 265 197 
rect 264 228 265 229 
rect 266 116 267 117 
rect 271 85 272 86 
rect 271 104 272 105 
rect 271 119 272 120 
rect 271 198 272 199 
rect 271 241 272 242 
rect 271 243 272 244 
rect 271 246 272 247 
rect 271 258 272 259 
rect 273 196 274 197 
rect 273 260 274 261 
rect 276 162 277 163 
rect 277 176 278 177 
rect 277 256 278 257 
rect 280 277 281 278 
rect 284 225 285 226 
rect 286 259 287 260 
rect 286 262 287 263 
rect 287 168 288 169 
rect 289 277 290 278 
rect 291 45 292 46 
rect 291 274 292 275 
rect 293 160 294 161 
rect 293 178 294 179 
rect 293 272 294 273 
rect 295 38 296 39 
<< end >>
3.99seconds.
