magic
tech scmos
timestamp1555213304
<< pdiffusion >>
<< polysilicon >>
rect 0 0 3 3 
rect 0 3 3 6 
rect 0 6 3 9 
rect 0 9 3 12 
rect 0 12 3 15 
rect 0 15 3 18 
rect 0 18 3 21 
rect 0 21 3 24 
rect 0 24 3 27 
rect 0 27 3 30 
rect 0 30 3 33 
rect 0 33 3 36 
rect 0 36 3 39 
rect 0 39 3 42 
rect 0 42 3 45 
rect 0 45 3 48 
rect 0 48 3 51 
rect 0 51 3 54 
rect 0 54 3 57 
rect 0 57 3 60 
rect 0 60 3 63 
rect 0 63 3 66 
rect 0 66 3 69 
rect 0 69 3 72 
rect 0 72 3 75 
rect 0 75 3 78 
rect 0 78 3 81 
rect 0 81 3 84 
rect 0 84 3 87 
rect 0 87 3 90 
rect 0 90 3 93 
rect 0 93 3 96 
rect 0 96 3 99 
rect 0 99 3 102 
rect 0 102 3 105 
rect 0 105 3 108 
rect 0 108 3 111 
rect 0 111 3 114 
rect 0 114 3 117 
rect 0 117 3 120 
rect 0 120 3 123 
rect 0 123 3 126 
rect 0 126 3 129 
rect 0 129 3 132 
rect 0 132 3 135 
rect 0 135 3 138 
rect 0 138 3 141 
rect 0 141 3 144 
rect 0 144 3 147 
rect 0 147 3 150 
rect 0 150 3 153 
rect 0 153 3 156 
rect 0 156 3 159 
rect 0 159 3 162 
rect 0 162 3 165 
rect 0 165 3 168 
rect 0 168 3 171 
rect 0 171 3 174 
rect 0 174 3 177 
rect 0 177 3 180 
rect 0 180 3 183 
rect 0 183 3 186 
rect 0 186 3 189 
rect 0 189 3 192 
rect 0 192 3 195 
rect 0 195 3 198 
rect 0 198 3 201 
rect 0 201 3 204 
rect 0 204 3 207 
rect 0 207 3 210 
rect 0 210 3 213 
rect 0 213 3 216 
rect 0 216 3 219 
rect 0 219 3 222 
rect 0 222 3 225 
rect 0 225 3 228 
rect 0 228 3 231 
rect 0 231 3 234 
rect 0 234 3 237 
rect 0 237 3 240 
rect 0 240 3 243 
rect 0 243 3 246 
rect 0 246 3 249 
rect 0 249 3 252 
rect 0 252 3 255 
rect 0 255 3 258 
rect 0 258 3 261 
rect 0 261 3 264 
rect 0 264 3 267 
rect 0 267 3 270 
rect 0 270 3 273 
rect 0 273 3 276 
rect 0 276 3 279 
rect 0 279 3 282 
rect 0 282 3 285 
rect 0 285 3 288 
rect 0 288 3 291 
rect 0 291 3 294 
rect 0 294 3 297 
rect 0 297 3 300 
rect 0 300 3 303 
rect 0 303 3 306 
rect 0 306 3 309 
rect 0 309 3 312 
rect 0 312 3 315 
rect 0 315 3 318 
rect 0 318 3 321 
rect 0 321 3 324 
rect 0 324 3 327 
rect 0 327 3 330 
rect 0 330 3 333 
rect 0 333 3 336 
rect 0 336 3 339 
rect 0 339 3 342 
rect 0 342 3 345 
rect 0 345 3 348 
rect 0 348 3 351 
rect 0 351 3 354 
rect 0 354 3 357 
rect 0 357 3 360 
rect 0 360 3 363 
rect 0 363 3 366 
rect 0 366 3 369 
rect 0 369 3 372 
rect 0 372 3 375 
rect 0 375 3 378 
rect 0 378 3 381 
rect 0 381 3 384 
rect 0 384 3 387 
rect 0 387 3 390 
rect 0 390 3 393 
rect 0 393 3 396 
rect 0 396 3 399 
rect 0 399 3 402 
rect 0 402 3 405 
rect 0 405 3 408 
rect 0 408 3 411 
rect 0 411 3 414 
rect 0 414 3 417 
rect 0 417 3 420 
rect 0 420 3 423 
rect 0 423 3 426 
rect 0 426 3 429 
rect 0 429 3 432 
rect 0 432 3 435 
rect 0 435 3 438 
rect 0 438 3 441 
rect 0 441 3 444 
rect 0 444 3 447 
rect 0 447 3 450 
rect 0 450 3 453 
rect 0 453 3 456 
rect 0 456 3 459 
rect 0 459 3 462 
rect 0 462 3 465 
rect 0 465 3 468 
rect 0 468 3 471 
rect 0 471 3 474 
rect 0 474 3 477 
rect 0 477 3 480 
rect 0 480 3 483 
rect 0 483 3 486 
rect 0 486 3 489 
rect 0 489 3 492 
rect 0 492 3 495 
rect 0 495 3 498 
rect 0 498 3 501 
rect 0 501 3 504 
rect 0 504 3 507 
rect 0 507 3 510 
rect 3 0 6 3 
rect 3 3 6 6 
rect 3 6 6 9 
rect 3 9 6 12 
rect 3 12 6 15 
rect 3 15 6 18 
rect 3 18 6 21 
rect 3 21 6 24 
rect 3 24 6 27 
rect 3 27 6 30 
rect 3 30 6 33 
rect 3 33 6 36 
rect 3 36 6 39 
rect 3 39 6 42 
rect 3 42 6 45 
rect 3 45 6 48 
rect 3 48 6 51 
rect 3 51 6 54 
rect 3 54 6 57 
rect 3 57 6 60 
rect 3 60 6 63 
rect 3 63 6 66 
rect 3 66 6 69 
rect 3 69 6 72 
rect 3 72 6 75 
rect 3 75 6 78 
rect 3 78 6 81 
rect 3 81 6 84 
rect 3 84 6 87 
rect 3 87 6 90 
rect 3 90 6 93 
rect 3 93 6 96 
rect 3 96 6 99 
rect 3 99 6 102 
rect 3 102 6 105 
rect 3 105 6 108 
rect 3 108 6 111 
rect 3 111 6 114 
rect 3 114 6 117 
rect 3 117 6 120 
rect 3 120 6 123 
rect 3 123 6 126 
rect 3 126 6 129 
rect 3 129 6 132 
rect 3 132 6 135 
rect 3 135 6 138 
rect 3 138 6 141 
rect 3 141 6 144 
rect 3 144 6 147 
rect 3 147 6 150 
rect 3 150 6 153 
rect 3 153 6 156 
rect 3 156 6 159 
rect 3 159 6 162 
rect 3 162 6 165 
rect 3 165 6 168 
rect 3 168 6 171 
rect 3 171 6 174 
rect 3 174 6 177 
rect 3 177 6 180 
rect 3 180 6 183 
rect 3 183 6 186 
rect 3 186 6 189 
rect 3 189 6 192 
rect 3 192 6 195 
rect 3 195 6 198 
rect 3 198 6 201 
rect 3 201 6 204 
rect 3 204 6 207 
rect 3 207 6 210 
rect 3 210 6 213 
rect 3 213 6 216 
rect 3 216 6 219 
rect 3 219 6 222 
rect 3 222 6 225 
rect 3 225 6 228 
rect 3 228 6 231 
rect 3 231 6 234 
rect 3 234 6 237 
rect 3 237 6 240 
rect 3 240 6 243 
rect 3 243 6 246 
rect 3 246 6 249 
rect 3 249 6 252 
rect 3 252 6 255 
rect 3 255 6 258 
rect 3 258 6 261 
rect 3 261 6 264 
rect 3 264 6 267 
rect 3 267 6 270 
rect 3 270 6 273 
rect 3 273 6 276 
rect 3 276 6 279 
rect 3 279 6 282 
rect 3 282 6 285 
rect 3 285 6 288 
rect 3 288 6 291 
rect 3 291 6 294 
rect 3 294 6 297 
rect 3 297 6 300 
rect 3 300 6 303 
rect 3 303 6 306 
rect 3 306 6 309 
rect 3 309 6 312 
rect 3 312 6 315 
rect 3 315 6 318 
rect 3 318 6 321 
rect 3 321 6 324 
rect 3 324 6 327 
rect 3 327 6 330 
rect 3 330 6 333 
rect 3 333 6 336 
rect 3 336 6 339 
rect 3 339 6 342 
rect 3 342 6 345 
rect 3 345 6 348 
rect 3 348 6 351 
rect 3 351 6 354 
rect 3 354 6 357 
rect 3 357 6 360 
rect 3 360 6 363 
rect 3 363 6 366 
rect 3 366 6 369 
rect 3 369 6 372 
rect 3 372 6 375 
rect 3 375 6 378 
rect 3 378 6 381 
rect 3 381 6 384 
rect 3 384 6 387 
rect 3 387 6 390 
rect 3 390 6 393 
rect 3 393 6 396 
rect 3 396 6 399 
rect 3 399 6 402 
rect 3 402 6 405 
rect 3 405 6 408 
rect 3 408 6 411 
rect 3 411 6 414 
rect 3 414 6 417 
rect 3 417 6 420 
rect 3 420 6 423 
rect 3 423 6 426 
rect 3 426 6 429 
rect 3 429 6 432 
rect 3 432 6 435 
rect 3 435 6 438 
rect 3 438 6 441 
rect 3 441 6 444 
rect 3 444 6 447 
rect 3 447 6 450 
rect 3 450 6 453 
rect 3 453 6 456 
rect 3 456 6 459 
rect 3 459 6 462 
rect 3 462 6 465 
rect 3 465 6 468 
rect 3 468 6 471 
rect 3 471 6 474 
rect 3 474 6 477 
rect 3 477 6 480 
rect 3 480 6 483 
rect 3 483 6 486 
rect 3 486 6 489 
rect 3 489 6 492 
rect 3 492 6 495 
rect 3 495 6 498 
rect 3 498 6 501 
rect 3 501 6 504 
rect 3 504 6 507 
rect 3 507 6 510 
rect 6 0 9 3 
rect 6 3 9 6 
rect 6 6 9 9 
rect 6 9 9 12 
rect 6 12 9 15 
rect 6 15 9 18 
rect 6 18 9 21 
rect 6 21 9 24 
rect 6 24 9 27 
rect 6 27 9 30 
rect 6 30 9 33 
rect 6 33 9 36 
rect 6 36 9 39 
rect 6 39 9 42 
rect 6 42 9 45 
rect 6 45 9 48 
rect 6 48 9 51 
rect 6 51 9 54 
rect 6 54 9 57 
rect 6 57 9 60 
rect 6 60 9 63 
rect 6 63 9 66 
rect 6 66 9 69 
rect 6 69 9 72 
rect 6 72 9 75 
rect 6 75 9 78 
rect 6 78 9 81 
rect 6 81 9 84 
rect 6 84 9 87 
rect 6 87 9 90 
rect 6 90 9 93 
rect 6 93 9 96 
rect 6 96 9 99 
rect 6 99 9 102 
rect 6 102 9 105 
rect 6 105 9 108 
rect 6 108 9 111 
rect 6 111 9 114 
rect 6 114 9 117 
rect 6 117 9 120 
rect 6 120 9 123 
rect 6 123 9 126 
rect 6 126 9 129 
rect 6 129 9 132 
rect 6 132 9 135 
rect 6 135 9 138 
rect 6 138 9 141 
rect 6 141 9 144 
rect 6 144 9 147 
rect 6 147 9 150 
rect 6 150 9 153 
rect 6 153 9 156 
rect 6 156 9 159 
rect 6 159 9 162 
rect 6 162 9 165 
rect 6 165 9 168 
rect 6 168 9 171 
rect 6 171 9 174 
rect 6 174 9 177 
rect 6 177 9 180 
rect 6 180 9 183 
rect 6 183 9 186 
rect 6 186 9 189 
rect 6 189 9 192 
rect 6 192 9 195 
rect 6 195 9 198 
rect 6 198 9 201 
rect 6 201 9 204 
rect 6 204 9 207 
rect 6 207 9 210 
rect 6 210 9 213 
rect 6 213 9 216 
rect 6 216 9 219 
rect 6 219 9 222 
rect 6 222 9 225 
rect 6 225 9 228 
rect 6 228 9 231 
rect 6 231 9 234 
rect 6 234 9 237 
rect 6 237 9 240 
rect 6 240 9 243 
rect 6 243 9 246 
rect 6 246 9 249 
rect 6 249 9 252 
rect 6 252 9 255 
rect 6 255 9 258 
rect 6 258 9 261 
rect 6 261 9 264 
rect 6 264 9 267 
rect 6 267 9 270 
rect 6 270 9 273 
rect 6 273 9 276 
rect 6 276 9 279 
rect 6 279 9 282 
rect 6 282 9 285 
rect 6 285 9 288 
rect 6 288 9 291 
rect 6 291 9 294 
rect 6 294 9 297 
rect 6 297 9 300 
rect 6 300 9 303 
rect 6 303 9 306 
rect 6 306 9 309 
rect 6 309 9 312 
rect 6 312 9 315 
rect 6 315 9 318 
rect 6 318 9 321 
rect 6 321 9 324 
rect 6 324 9 327 
rect 6 327 9 330 
rect 6 330 9 333 
rect 6 333 9 336 
rect 6 336 9 339 
rect 6 339 9 342 
rect 6 342 9 345 
rect 6 345 9 348 
rect 6 348 9 351 
rect 6 351 9 354 
rect 6 354 9 357 
rect 6 357 9 360 
rect 6 360 9 363 
rect 6 363 9 366 
rect 6 366 9 369 
rect 6 369 9 372 
rect 6 372 9 375 
rect 6 375 9 378 
rect 6 378 9 381 
rect 6 381 9 384 
rect 6 384 9 387 
rect 6 387 9 390 
rect 6 390 9 393 
rect 6 393 9 396 
rect 6 396 9 399 
rect 6 399 9 402 
rect 6 402 9 405 
rect 6 405 9 408 
rect 6 408 9 411 
rect 6 411 9 414 
rect 6 414 9 417 
rect 6 417 9 420 
rect 6 420 9 423 
rect 6 423 9 426 
rect 6 426 9 429 
rect 6 429 9 432 
rect 6 432 9 435 
rect 6 435 9 438 
rect 6 438 9 441 
rect 6 441 9 444 
rect 6 444 9 447 
rect 6 447 9 450 
rect 6 450 9 453 
rect 6 453 9 456 
rect 6 456 9 459 
rect 6 459 9 462 
rect 6 462 9 465 
rect 6 465 9 468 
rect 6 468 9 471 
rect 6 471 9 474 
rect 6 474 9 477 
rect 6 477 9 480 
rect 6 480 9 483 
rect 6 483 9 486 
rect 6 486 9 489 
rect 6 489 9 492 
rect 6 492 9 495 
rect 6 495 9 498 
rect 6 498 9 501 
rect 6 501 9 504 
rect 6 504 9 507 
rect 6 507 9 510 
rect 9 0 12 3 
rect 9 3 12 6 
rect 9 6 12 9 
rect 9 9 12 12 
rect 9 12 12 15 
rect 9 15 12 18 
rect 9 18 12 21 
rect 9 21 12 24 
rect 9 24 12 27 
rect 9 27 12 30 
rect 9 30 12 33 
rect 9 33 12 36 
rect 9 36 12 39 
rect 9 39 12 42 
rect 9 42 12 45 
rect 9 45 12 48 
rect 9 48 12 51 
rect 9 51 12 54 
rect 9 54 12 57 
rect 9 57 12 60 
rect 9 60 12 63 
rect 9 63 12 66 
rect 9 66 12 69 
rect 9 69 12 72 
rect 9 72 12 75 
rect 9 75 12 78 
rect 9 78 12 81 
rect 9 81 12 84 
rect 9 84 12 87 
rect 9 87 12 90 
rect 9 90 12 93 
rect 9 93 12 96 
rect 9 96 12 99 
rect 9 99 12 102 
rect 9 102 12 105 
rect 9 105 12 108 
rect 9 108 12 111 
rect 9 111 12 114 
rect 9 114 12 117 
rect 9 117 12 120 
rect 9 120 12 123 
rect 9 123 12 126 
rect 9 126 12 129 
rect 9 129 12 132 
rect 9 132 12 135 
rect 9 135 12 138 
rect 9 138 12 141 
rect 9 141 12 144 
rect 9 144 12 147 
rect 9 147 12 150 
rect 9 150 12 153 
rect 9 153 12 156 
rect 9 156 12 159 
rect 9 159 12 162 
rect 9 162 12 165 
rect 9 165 12 168 
rect 9 168 12 171 
rect 9 171 12 174 
rect 9 174 12 177 
rect 9 177 12 180 
rect 9 180 12 183 
rect 9 183 12 186 
rect 9 186 12 189 
rect 9 189 12 192 
rect 9 192 12 195 
rect 9 195 12 198 
rect 9 198 12 201 
rect 9 201 12 204 
rect 9 204 12 207 
rect 9 207 12 210 
rect 9 210 12 213 
rect 9 213 12 216 
rect 9 216 12 219 
rect 9 219 12 222 
rect 9 222 12 225 
rect 9 225 12 228 
rect 9 228 12 231 
rect 9 231 12 234 
rect 9 234 12 237 
rect 9 237 12 240 
rect 9 240 12 243 
rect 9 243 12 246 
rect 9 246 12 249 
rect 9 249 12 252 
rect 9 252 12 255 
rect 9 255 12 258 
rect 9 258 12 261 
rect 9 261 12 264 
rect 9 264 12 267 
rect 9 267 12 270 
rect 9 270 12 273 
rect 9 273 12 276 
rect 9 276 12 279 
rect 9 279 12 282 
rect 9 282 12 285 
rect 9 285 12 288 
rect 9 288 12 291 
rect 9 291 12 294 
rect 9 294 12 297 
rect 9 297 12 300 
rect 9 300 12 303 
rect 9 303 12 306 
rect 9 306 12 309 
rect 9 309 12 312 
rect 9 312 12 315 
rect 9 315 12 318 
rect 9 318 12 321 
rect 9 321 12 324 
rect 9 324 12 327 
rect 9 327 12 330 
rect 9 330 12 333 
rect 9 333 12 336 
rect 9 336 12 339 
rect 9 339 12 342 
rect 9 342 12 345 
rect 9 345 12 348 
rect 9 348 12 351 
rect 9 351 12 354 
rect 9 354 12 357 
rect 9 357 12 360 
rect 9 360 12 363 
rect 9 363 12 366 
rect 9 366 12 369 
rect 9 369 12 372 
rect 9 372 12 375 
rect 9 375 12 378 
rect 9 378 12 381 
rect 9 381 12 384 
rect 9 384 12 387 
rect 9 387 12 390 
rect 9 390 12 393 
rect 9 393 12 396 
rect 9 396 12 399 
rect 9 399 12 402 
rect 9 402 12 405 
rect 9 405 12 408 
rect 9 408 12 411 
rect 9 411 12 414 
rect 9 414 12 417 
rect 9 417 12 420 
rect 9 420 12 423 
rect 9 423 12 426 
rect 9 426 12 429 
rect 9 429 12 432 
rect 9 432 12 435 
rect 9 435 12 438 
rect 9 438 12 441 
rect 9 441 12 444 
rect 9 444 12 447 
rect 9 447 12 450 
rect 9 450 12 453 
rect 9 453 12 456 
rect 9 456 12 459 
rect 9 459 12 462 
rect 9 462 12 465 
rect 9 465 12 468 
rect 9 468 12 471 
rect 9 471 12 474 
rect 9 474 12 477 
rect 9 477 12 480 
rect 9 480 12 483 
rect 9 483 12 486 
rect 9 486 12 489 
rect 9 489 12 492 
rect 9 492 12 495 
rect 9 495 12 498 
rect 9 498 12 501 
rect 9 501 12 504 
rect 9 504 12 507 
rect 9 507 12 510 
rect 12 0 15 3 
rect 12 3 15 6 
rect 12 6 15 9 
rect 12 9 15 12 
rect 12 12 15 15 
rect 12 15 15 18 
rect 12 18 15 21 
rect 12 21 15 24 
rect 12 24 15 27 
rect 12 27 15 30 
rect 12 30 15 33 
rect 12 33 15 36 
rect 12 36 15 39 
rect 12 39 15 42 
rect 12 42 15 45 
rect 12 45 15 48 
rect 12 48 15 51 
rect 12 51 15 54 
rect 12 54 15 57 
rect 12 57 15 60 
rect 12 60 15 63 
rect 12 63 15 66 
rect 12 66 15 69 
rect 12 69 15 72 
rect 12 72 15 75 
rect 12 75 15 78 
rect 12 78 15 81 
rect 12 81 15 84 
rect 12 84 15 87 
rect 12 87 15 90 
rect 12 90 15 93 
rect 12 93 15 96 
rect 12 96 15 99 
rect 12 99 15 102 
rect 12 102 15 105 
rect 12 105 15 108 
rect 12 108 15 111 
rect 12 111 15 114 
rect 12 114 15 117 
rect 12 117 15 120 
rect 12 120 15 123 
rect 12 123 15 126 
rect 12 126 15 129 
rect 12 129 15 132 
rect 12 132 15 135 
rect 12 135 15 138 
rect 12 138 15 141 
rect 12 141 15 144 
rect 12 144 15 147 
rect 12 147 15 150 
rect 12 150 15 153 
rect 12 153 15 156 
rect 12 156 15 159 
rect 12 159 15 162 
rect 12 162 15 165 
rect 12 165 15 168 
rect 12 168 15 171 
rect 12 171 15 174 
rect 12 174 15 177 
rect 12 177 15 180 
rect 12 180 15 183 
rect 12 183 15 186 
rect 12 186 15 189 
rect 12 189 15 192 
rect 12 192 15 195 
rect 12 195 15 198 
rect 12 198 15 201 
rect 12 201 15 204 
rect 12 204 15 207 
rect 12 207 15 210 
rect 12 210 15 213 
rect 12 213 15 216 
rect 12 216 15 219 
rect 12 219 15 222 
rect 12 222 15 225 
rect 12 225 15 228 
rect 12 228 15 231 
rect 12 231 15 234 
rect 12 234 15 237 
rect 12 237 15 240 
rect 12 240 15 243 
rect 12 243 15 246 
rect 12 246 15 249 
rect 12 249 15 252 
rect 12 252 15 255 
rect 12 255 15 258 
rect 12 258 15 261 
rect 12 261 15 264 
rect 12 264 15 267 
rect 12 267 15 270 
rect 12 270 15 273 
rect 12 273 15 276 
rect 12 276 15 279 
rect 12 279 15 282 
rect 12 282 15 285 
rect 12 285 15 288 
rect 12 288 15 291 
rect 12 291 15 294 
rect 12 294 15 297 
rect 12 297 15 300 
rect 12 300 15 303 
rect 12 303 15 306 
rect 12 306 15 309 
rect 12 309 15 312 
rect 12 312 15 315 
rect 12 315 15 318 
rect 12 318 15 321 
rect 12 321 15 324 
rect 12 324 15 327 
rect 12 327 15 330 
rect 12 330 15 333 
rect 12 333 15 336 
rect 12 336 15 339 
rect 12 339 15 342 
rect 12 342 15 345 
rect 12 345 15 348 
rect 12 348 15 351 
rect 12 351 15 354 
rect 12 354 15 357 
rect 12 357 15 360 
rect 12 360 15 363 
rect 12 363 15 366 
rect 12 366 15 369 
rect 12 369 15 372 
rect 12 372 15 375 
rect 12 375 15 378 
rect 12 378 15 381 
rect 12 381 15 384 
rect 12 384 15 387 
rect 12 387 15 390 
rect 12 390 15 393 
rect 12 393 15 396 
rect 12 396 15 399 
rect 12 399 15 402 
rect 12 402 15 405 
rect 12 405 15 408 
rect 12 408 15 411 
rect 12 411 15 414 
rect 12 414 15 417 
rect 12 417 15 420 
rect 12 420 15 423 
rect 12 423 15 426 
rect 12 426 15 429 
rect 12 429 15 432 
rect 12 432 15 435 
rect 12 435 15 438 
rect 12 438 15 441 
rect 12 441 15 444 
rect 12 444 15 447 
rect 12 447 15 450 
rect 12 450 15 453 
rect 12 453 15 456 
rect 12 456 15 459 
rect 12 459 15 462 
rect 12 462 15 465 
rect 12 465 15 468 
rect 12 468 15 471 
rect 12 471 15 474 
rect 12 474 15 477 
rect 12 477 15 480 
rect 12 480 15 483 
rect 12 483 15 486 
rect 12 486 15 489 
rect 12 489 15 492 
rect 12 492 15 495 
rect 12 495 15 498 
rect 12 498 15 501 
rect 12 501 15 504 
rect 12 504 15 507 
rect 12 507 15 510 
rect 15 0 18 3 
rect 15 3 18 6 
rect 15 6 18 9 
rect 15 9 18 12 
rect 15 12 18 15 
rect 15 15 18 18 
rect 15 18 18 21 
rect 15 21 18 24 
rect 15 24 18 27 
rect 15 27 18 30 
rect 15 30 18 33 
rect 15 33 18 36 
rect 15 36 18 39 
rect 15 39 18 42 
rect 15 42 18 45 
rect 15 45 18 48 
rect 15 48 18 51 
rect 15 51 18 54 
rect 15 54 18 57 
rect 15 57 18 60 
rect 15 60 18 63 
rect 15 63 18 66 
rect 15 66 18 69 
rect 15 69 18 72 
rect 15 72 18 75 
rect 15 75 18 78 
rect 15 78 18 81 
rect 15 81 18 84 
rect 15 84 18 87 
rect 15 87 18 90 
rect 15 90 18 93 
rect 15 93 18 96 
rect 15 96 18 99 
rect 15 99 18 102 
rect 15 102 18 105 
rect 15 105 18 108 
rect 15 108 18 111 
rect 15 111 18 114 
rect 15 114 18 117 
rect 15 117 18 120 
rect 15 120 18 123 
rect 15 123 18 126 
rect 15 126 18 129 
rect 15 129 18 132 
rect 15 132 18 135 
rect 15 135 18 138 
rect 15 138 18 141 
rect 15 141 18 144 
rect 15 144 18 147 
rect 15 147 18 150 
rect 15 150 18 153 
rect 15 153 18 156 
rect 15 156 18 159 
rect 15 159 18 162 
rect 15 162 18 165 
rect 15 165 18 168 
rect 15 168 18 171 
rect 15 171 18 174 
rect 15 174 18 177 
rect 15 177 18 180 
rect 15 180 18 183 
rect 15 183 18 186 
rect 15 186 18 189 
rect 15 189 18 192 
rect 15 192 18 195 
rect 15 195 18 198 
rect 15 198 18 201 
rect 15 201 18 204 
rect 15 204 18 207 
rect 15 207 18 210 
rect 15 210 18 213 
rect 15 213 18 216 
rect 15 216 18 219 
rect 15 219 18 222 
rect 15 222 18 225 
rect 15 225 18 228 
rect 15 228 18 231 
rect 15 231 18 234 
rect 15 234 18 237 
rect 15 237 18 240 
rect 15 240 18 243 
rect 15 243 18 246 
rect 15 246 18 249 
rect 15 249 18 252 
rect 15 252 18 255 
rect 15 255 18 258 
rect 15 258 18 261 
rect 15 261 18 264 
rect 15 264 18 267 
rect 15 267 18 270 
rect 15 270 18 273 
rect 15 273 18 276 
rect 15 276 18 279 
rect 15 279 18 282 
rect 15 282 18 285 
rect 15 285 18 288 
rect 15 288 18 291 
rect 15 291 18 294 
rect 15 294 18 297 
rect 15 297 18 300 
rect 15 300 18 303 
rect 15 303 18 306 
rect 15 306 18 309 
rect 15 309 18 312 
rect 15 312 18 315 
rect 15 315 18 318 
rect 15 318 18 321 
rect 15 321 18 324 
rect 15 324 18 327 
rect 15 327 18 330 
rect 15 330 18 333 
rect 15 333 18 336 
rect 15 336 18 339 
rect 15 339 18 342 
rect 15 342 18 345 
rect 15 345 18 348 
rect 15 348 18 351 
rect 15 351 18 354 
rect 15 354 18 357 
rect 15 357 18 360 
rect 15 360 18 363 
rect 15 363 18 366 
rect 15 366 18 369 
rect 15 369 18 372 
rect 15 372 18 375 
rect 15 375 18 378 
rect 15 378 18 381 
rect 15 381 18 384 
rect 15 384 18 387 
rect 15 387 18 390 
rect 15 390 18 393 
rect 15 393 18 396 
rect 15 396 18 399 
rect 15 399 18 402 
rect 15 402 18 405 
rect 15 405 18 408 
rect 15 408 18 411 
rect 15 411 18 414 
rect 15 414 18 417 
rect 15 417 18 420 
rect 15 420 18 423 
rect 15 423 18 426 
rect 15 426 18 429 
rect 15 429 18 432 
rect 15 432 18 435 
rect 15 435 18 438 
rect 15 438 18 441 
rect 15 441 18 444 
rect 15 444 18 447 
rect 15 447 18 450 
rect 15 450 18 453 
rect 15 453 18 456 
rect 15 456 18 459 
rect 15 459 18 462 
rect 15 462 18 465 
rect 15 465 18 468 
rect 15 468 18 471 
rect 15 471 18 474 
rect 15 474 18 477 
rect 15 477 18 480 
rect 15 480 18 483 
rect 15 483 18 486 
rect 15 486 18 489 
rect 15 489 18 492 
rect 15 492 18 495 
rect 15 495 18 498 
rect 15 498 18 501 
rect 15 501 18 504 
rect 15 504 18 507 
rect 15 507 18 510 
rect 18 0 21 3 
rect 18 3 21 6 
rect 18 6 21 9 
rect 18 9 21 12 
rect 18 12 21 15 
rect 18 15 21 18 
rect 18 18 21 21 
rect 18 21 21 24 
rect 18 24 21 27 
rect 18 27 21 30 
rect 18 30 21 33 
rect 18 33 21 36 
rect 18 36 21 39 
rect 18 39 21 42 
rect 18 42 21 45 
rect 18 45 21 48 
rect 18 48 21 51 
rect 18 51 21 54 
rect 18 54 21 57 
rect 18 57 21 60 
rect 18 60 21 63 
rect 18 63 21 66 
rect 18 66 21 69 
rect 18 69 21 72 
rect 18 72 21 75 
rect 18 75 21 78 
rect 18 78 21 81 
rect 18 81 21 84 
rect 18 84 21 87 
rect 18 87 21 90 
rect 18 90 21 93 
rect 18 93 21 96 
rect 18 96 21 99 
rect 18 99 21 102 
rect 18 102 21 105 
rect 18 105 21 108 
rect 18 108 21 111 
rect 18 111 21 114 
rect 18 114 21 117 
rect 18 117 21 120 
rect 18 120 21 123 
rect 18 123 21 126 
rect 18 126 21 129 
rect 18 129 21 132 
rect 18 132 21 135 
rect 18 135 21 138 
rect 18 138 21 141 
rect 18 141 21 144 
rect 18 144 21 147 
rect 18 147 21 150 
rect 18 150 21 153 
rect 18 153 21 156 
rect 18 156 21 159 
rect 18 159 21 162 
rect 18 162 21 165 
rect 18 165 21 168 
rect 18 168 21 171 
rect 18 171 21 174 
rect 18 174 21 177 
rect 18 177 21 180 
rect 18 180 21 183 
rect 18 183 21 186 
rect 18 186 21 189 
rect 18 189 21 192 
rect 18 192 21 195 
rect 18 195 21 198 
rect 18 198 21 201 
rect 18 201 21 204 
rect 18 204 21 207 
rect 18 207 21 210 
rect 18 210 21 213 
rect 18 213 21 216 
rect 18 216 21 219 
rect 18 219 21 222 
rect 18 222 21 225 
rect 18 225 21 228 
rect 18 228 21 231 
rect 18 231 21 234 
rect 18 234 21 237 
rect 18 237 21 240 
rect 18 240 21 243 
rect 18 243 21 246 
rect 18 246 21 249 
rect 18 249 21 252 
rect 18 252 21 255 
rect 18 255 21 258 
rect 18 258 21 261 
rect 18 261 21 264 
rect 18 264 21 267 
rect 18 267 21 270 
rect 18 270 21 273 
rect 18 273 21 276 
rect 18 276 21 279 
rect 18 279 21 282 
rect 18 282 21 285 
rect 18 285 21 288 
rect 18 288 21 291 
rect 18 291 21 294 
rect 18 294 21 297 
rect 18 297 21 300 
rect 18 300 21 303 
rect 18 303 21 306 
rect 18 306 21 309 
rect 18 309 21 312 
rect 18 312 21 315 
rect 18 315 21 318 
rect 18 318 21 321 
rect 18 321 21 324 
rect 18 324 21 327 
rect 18 327 21 330 
rect 18 330 21 333 
rect 18 333 21 336 
rect 18 336 21 339 
rect 18 339 21 342 
rect 18 342 21 345 
rect 18 345 21 348 
rect 18 348 21 351 
rect 18 351 21 354 
rect 18 354 21 357 
rect 18 357 21 360 
rect 18 360 21 363 
rect 18 363 21 366 
rect 18 366 21 369 
rect 18 369 21 372 
rect 18 372 21 375 
rect 18 375 21 378 
rect 18 378 21 381 
rect 18 381 21 384 
rect 18 384 21 387 
rect 18 387 21 390 
rect 18 390 21 393 
rect 18 393 21 396 
rect 18 396 21 399 
rect 18 399 21 402 
rect 18 402 21 405 
rect 18 405 21 408 
rect 18 408 21 411 
rect 18 411 21 414 
rect 18 414 21 417 
rect 18 417 21 420 
rect 18 420 21 423 
rect 18 423 21 426 
rect 18 426 21 429 
rect 18 429 21 432 
rect 18 432 21 435 
rect 18 435 21 438 
rect 18 438 21 441 
rect 18 441 21 444 
rect 18 444 21 447 
rect 18 447 21 450 
rect 18 450 21 453 
rect 18 453 21 456 
rect 18 456 21 459 
rect 18 459 21 462 
rect 18 462 21 465 
rect 18 465 21 468 
rect 18 468 21 471 
rect 18 471 21 474 
rect 18 474 21 477 
rect 18 477 21 480 
rect 18 480 21 483 
rect 18 483 21 486 
rect 18 486 21 489 
rect 18 489 21 492 
rect 18 492 21 495 
rect 18 495 21 498 
rect 18 498 21 501 
rect 18 501 21 504 
rect 18 504 21 507 
rect 18 507 21 510 
rect 21 0 24 3 
rect 21 3 24 6 
rect 21 6 24 9 
rect 21 9 24 12 
rect 21 12 24 15 
rect 21 15 24 18 
rect 21 18 24 21 
rect 21 21 24 24 
rect 21 24 24 27 
rect 21 27 24 30 
rect 21 30 24 33 
rect 21 33 24 36 
rect 21 36 24 39 
rect 21 39 24 42 
rect 21 42 24 45 
rect 21 45 24 48 
rect 21 48 24 51 
rect 21 51 24 54 
rect 21 54 24 57 
rect 21 57 24 60 
rect 21 60 24 63 
rect 21 63 24 66 
rect 21 66 24 69 
rect 21 69 24 72 
rect 21 72 24 75 
rect 21 75 24 78 
rect 21 78 24 81 
rect 21 81 24 84 
rect 21 84 24 87 
rect 21 87 24 90 
rect 21 90 24 93 
rect 21 93 24 96 
rect 21 96 24 99 
rect 21 99 24 102 
rect 21 102 24 105 
rect 21 105 24 108 
rect 21 108 24 111 
rect 21 111 24 114 
rect 21 114 24 117 
rect 21 117 24 120 
rect 21 120 24 123 
rect 21 123 24 126 
rect 21 126 24 129 
rect 21 129 24 132 
rect 21 132 24 135 
rect 21 135 24 138 
rect 21 138 24 141 
rect 21 141 24 144 
rect 21 144 24 147 
rect 21 147 24 150 
rect 21 150 24 153 
rect 21 153 24 156 
rect 21 156 24 159 
rect 21 159 24 162 
rect 21 162 24 165 
rect 21 165 24 168 
rect 21 168 24 171 
rect 21 171 24 174 
rect 21 174 24 177 
rect 21 177 24 180 
rect 21 180 24 183 
rect 21 183 24 186 
rect 21 186 24 189 
rect 21 189 24 192 
rect 21 192 24 195 
rect 21 195 24 198 
rect 21 198 24 201 
rect 21 201 24 204 
rect 21 204 24 207 
rect 21 207 24 210 
rect 21 210 24 213 
rect 21 213 24 216 
rect 21 216 24 219 
rect 21 219 24 222 
rect 21 222 24 225 
rect 21 225 24 228 
rect 21 228 24 231 
rect 21 231 24 234 
rect 21 234 24 237 
rect 21 237 24 240 
rect 21 240 24 243 
rect 21 243 24 246 
rect 21 246 24 249 
rect 21 249 24 252 
rect 21 252 24 255 
rect 21 255 24 258 
rect 21 258 24 261 
rect 21 261 24 264 
rect 21 264 24 267 
rect 21 267 24 270 
rect 21 270 24 273 
rect 21 273 24 276 
rect 21 276 24 279 
rect 21 279 24 282 
rect 21 282 24 285 
rect 21 285 24 288 
rect 21 288 24 291 
rect 21 291 24 294 
rect 21 294 24 297 
rect 21 297 24 300 
rect 21 300 24 303 
rect 21 303 24 306 
rect 21 306 24 309 
rect 21 309 24 312 
rect 21 312 24 315 
rect 21 315 24 318 
rect 21 318 24 321 
rect 21 321 24 324 
rect 21 324 24 327 
rect 21 327 24 330 
rect 21 330 24 333 
rect 21 333 24 336 
rect 21 336 24 339 
rect 21 339 24 342 
rect 21 342 24 345 
rect 21 345 24 348 
rect 21 348 24 351 
rect 21 351 24 354 
rect 21 354 24 357 
rect 21 357 24 360 
rect 21 360 24 363 
rect 21 363 24 366 
rect 21 366 24 369 
rect 21 369 24 372 
rect 21 372 24 375 
rect 21 375 24 378 
rect 21 378 24 381 
rect 21 381 24 384 
rect 21 384 24 387 
rect 21 387 24 390 
rect 21 390 24 393 
rect 21 393 24 396 
rect 21 396 24 399 
rect 21 399 24 402 
rect 21 402 24 405 
rect 21 405 24 408 
rect 21 408 24 411 
rect 21 411 24 414 
rect 21 414 24 417 
rect 21 417 24 420 
rect 21 420 24 423 
rect 21 423 24 426 
rect 21 426 24 429 
rect 21 429 24 432 
rect 21 432 24 435 
rect 21 435 24 438 
rect 21 438 24 441 
rect 21 441 24 444 
rect 21 444 24 447 
rect 21 447 24 450 
rect 21 450 24 453 
rect 21 453 24 456 
rect 21 456 24 459 
rect 21 459 24 462 
rect 21 462 24 465 
rect 21 465 24 468 
rect 21 468 24 471 
rect 21 471 24 474 
rect 21 474 24 477 
rect 21 477 24 480 
rect 21 480 24 483 
rect 21 483 24 486 
rect 21 486 24 489 
rect 21 489 24 492 
rect 21 492 24 495 
rect 21 495 24 498 
rect 21 498 24 501 
rect 21 501 24 504 
rect 21 504 24 507 
rect 21 507 24 510 
rect 24 0 27 3 
rect 24 3 27 6 
rect 24 6 27 9 
rect 24 9 27 12 
rect 24 12 27 15 
rect 24 15 27 18 
rect 24 18 27 21 
rect 24 21 27 24 
rect 24 24 27 27 
rect 24 27 27 30 
rect 24 30 27 33 
rect 24 33 27 36 
rect 24 36 27 39 
rect 24 39 27 42 
rect 24 42 27 45 
rect 24 45 27 48 
rect 24 48 27 51 
rect 24 51 27 54 
rect 24 54 27 57 
rect 24 57 27 60 
rect 24 60 27 63 
rect 24 63 27 66 
rect 24 66 27 69 
rect 24 69 27 72 
rect 24 72 27 75 
rect 24 75 27 78 
rect 24 78 27 81 
rect 24 81 27 84 
rect 24 84 27 87 
rect 24 87 27 90 
rect 24 90 27 93 
rect 24 93 27 96 
rect 24 96 27 99 
rect 24 99 27 102 
rect 24 102 27 105 
rect 24 105 27 108 
rect 24 108 27 111 
rect 24 111 27 114 
rect 24 114 27 117 
rect 24 117 27 120 
rect 24 120 27 123 
rect 24 123 27 126 
rect 24 126 27 129 
rect 24 129 27 132 
rect 24 132 27 135 
rect 24 135 27 138 
rect 24 138 27 141 
rect 24 141 27 144 
rect 24 144 27 147 
rect 24 147 27 150 
rect 24 150 27 153 
rect 24 153 27 156 
rect 24 156 27 159 
rect 24 159 27 162 
rect 24 162 27 165 
rect 24 165 27 168 
rect 24 168 27 171 
rect 24 171 27 174 
rect 24 174 27 177 
rect 24 177 27 180 
rect 24 180 27 183 
rect 24 183 27 186 
rect 24 186 27 189 
rect 24 189 27 192 
rect 24 192 27 195 
rect 24 195 27 198 
rect 24 198 27 201 
rect 24 201 27 204 
rect 24 204 27 207 
rect 24 207 27 210 
rect 24 210 27 213 
rect 24 213 27 216 
rect 24 216 27 219 
rect 24 219 27 222 
rect 24 222 27 225 
rect 24 225 27 228 
rect 24 228 27 231 
rect 24 231 27 234 
rect 24 234 27 237 
rect 24 237 27 240 
rect 24 240 27 243 
rect 24 243 27 246 
rect 24 246 27 249 
rect 24 249 27 252 
rect 24 252 27 255 
rect 24 255 27 258 
rect 24 258 27 261 
rect 24 261 27 264 
rect 24 264 27 267 
rect 24 267 27 270 
rect 24 270 27 273 
rect 24 273 27 276 
rect 24 276 27 279 
rect 24 279 27 282 
rect 24 282 27 285 
rect 24 285 27 288 
rect 24 288 27 291 
rect 24 291 27 294 
rect 24 294 27 297 
rect 24 297 27 300 
rect 24 300 27 303 
rect 24 303 27 306 
rect 24 306 27 309 
rect 24 309 27 312 
rect 24 312 27 315 
rect 24 315 27 318 
rect 24 318 27 321 
rect 24 321 27 324 
rect 24 324 27 327 
rect 24 327 27 330 
rect 24 330 27 333 
rect 24 333 27 336 
rect 24 336 27 339 
rect 24 339 27 342 
rect 24 342 27 345 
rect 24 345 27 348 
rect 24 348 27 351 
rect 24 351 27 354 
rect 24 354 27 357 
rect 24 357 27 360 
rect 24 360 27 363 
rect 24 363 27 366 
rect 24 366 27 369 
rect 24 369 27 372 
rect 24 372 27 375 
rect 24 375 27 378 
rect 24 378 27 381 
rect 24 381 27 384 
rect 24 384 27 387 
rect 24 387 27 390 
rect 24 390 27 393 
rect 24 393 27 396 
rect 24 396 27 399 
rect 24 399 27 402 
rect 24 402 27 405 
rect 24 405 27 408 
rect 24 408 27 411 
rect 24 411 27 414 
rect 24 414 27 417 
rect 24 417 27 420 
rect 24 420 27 423 
rect 24 423 27 426 
rect 24 426 27 429 
rect 24 429 27 432 
rect 24 432 27 435 
rect 24 435 27 438 
rect 24 438 27 441 
rect 24 441 27 444 
rect 24 444 27 447 
rect 24 447 27 450 
rect 24 450 27 453 
rect 24 453 27 456 
rect 24 456 27 459 
rect 24 459 27 462 
rect 24 462 27 465 
rect 24 465 27 468 
rect 24 468 27 471 
rect 24 471 27 474 
rect 24 474 27 477 
rect 24 477 27 480 
rect 24 480 27 483 
rect 24 483 27 486 
rect 24 486 27 489 
rect 24 489 27 492 
rect 24 492 27 495 
rect 24 495 27 498 
rect 24 498 27 501 
rect 24 501 27 504 
rect 24 504 27 507 
rect 24 507 27 510 
rect 27 0 30 3 
rect 27 3 30 6 
rect 27 6 30 9 
rect 27 9 30 12 
rect 27 12 30 15 
rect 27 15 30 18 
rect 27 18 30 21 
rect 27 21 30 24 
rect 27 24 30 27 
rect 27 27 30 30 
rect 27 30 30 33 
rect 27 33 30 36 
rect 27 36 30 39 
rect 27 39 30 42 
rect 27 42 30 45 
rect 27 45 30 48 
rect 27 48 30 51 
rect 27 51 30 54 
rect 27 54 30 57 
rect 27 57 30 60 
rect 27 60 30 63 
rect 27 63 30 66 
rect 27 66 30 69 
rect 27 69 30 72 
rect 27 72 30 75 
rect 27 75 30 78 
rect 27 78 30 81 
rect 27 81 30 84 
rect 27 84 30 87 
rect 27 87 30 90 
rect 27 90 30 93 
rect 27 93 30 96 
rect 27 96 30 99 
rect 27 99 30 102 
rect 27 102 30 105 
rect 27 105 30 108 
rect 27 108 30 111 
rect 27 111 30 114 
rect 27 114 30 117 
rect 27 117 30 120 
rect 27 120 30 123 
rect 27 123 30 126 
rect 27 126 30 129 
rect 27 129 30 132 
rect 27 132 30 135 
rect 27 135 30 138 
rect 27 138 30 141 
rect 27 141 30 144 
rect 27 144 30 147 
rect 27 147 30 150 
rect 27 150 30 153 
rect 27 153 30 156 
rect 27 156 30 159 
rect 27 159 30 162 
rect 27 162 30 165 
rect 27 165 30 168 
rect 27 168 30 171 
rect 27 171 30 174 
rect 27 174 30 177 
rect 27 177 30 180 
rect 27 180 30 183 
rect 27 183 30 186 
rect 27 186 30 189 
rect 27 189 30 192 
rect 27 192 30 195 
rect 27 195 30 198 
rect 27 198 30 201 
rect 27 201 30 204 
rect 27 204 30 207 
rect 27 207 30 210 
rect 27 210 30 213 
rect 27 213 30 216 
rect 27 216 30 219 
rect 27 219 30 222 
rect 27 222 30 225 
rect 27 225 30 228 
rect 27 228 30 231 
rect 27 231 30 234 
rect 27 234 30 237 
rect 27 237 30 240 
rect 27 240 30 243 
rect 27 243 30 246 
rect 27 246 30 249 
rect 27 249 30 252 
rect 27 252 30 255 
rect 27 255 30 258 
rect 27 258 30 261 
rect 27 261 30 264 
rect 27 264 30 267 
rect 27 267 30 270 
rect 27 270 30 273 
rect 27 273 30 276 
rect 27 276 30 279 
rect 27 279 30 282 
rect 27 282 30 285 
rect 27 285 30 288 
rect 27 288 30 291 
rect 27 291 30 294 
rect 27 294 30 297 
rect 27 297 30 300 
rect 27 300 30 303 
rect 27 303 30 306 
rect 27 306 30 309 
rect 27 309 30 312 
rect 27 312 30 315 
rect 27 315 30 318 
rect 27 318 30 321 
rect 27 321 30 324 
rect 27 324 30 327 
rect 27 327 30 330 
rect 27 330 30 333 
rect 27 333 30 336 
rect 27 336 30 339 
rect 27 339 30 342 
rect 27 342 30 345 
rect 27 345 30 348 
rect 27 348 30 351 
rect 27 351 30 354 
rect 27 354 30 357 
rect 27 357 30 360 
rect 27 360 30 363 
rect 27 363 30 366 
rect 27 366 30 369 
rect 27 369 30 372 
rect 27 372 30 375 
rect 27 375 30 378 
rect 27 378 30 381 
rect 27 381 30 384 
rect 27 384 30 387 
rect 27 387 30 390 
rect 27 390 30 393 
rect 27 393 30 396 
rect 27 396 30 399 
rect 27 399 30 402 
rect 27 402 30 405 
rect 27 405 30 408 
rect 27 408 30 411 
rect 27 411 30 414 
rect 27 414 30 417 
rect 27 417 30 420 
rect 27 420 30 423 
rect 27 423 30 426 
rect 27 426 30 429 
rect 27 429 30 432 
rect 27 432 30 435 
rect 27 435 30 438 
rect 27 438 30 441 
rect 27 441 30 444 
rect 27 444 30 447 
rect 27 447 30 450 
rect 27 450 30 453 
rect 27 453 30 456 
rect 27 456 30 459 
rect 27 459 30 462 
rect 27 462 30 465 
rect 27 465 30 468 
rect 27 468 30 471 
rect 27 471 30 474 
rect 27 474 30 477 
rect 27 477 30 480 
rect 27 480 30 483 
rect 27 483 30 486 
rect 27 486 30 489 
rect 27 489 30 492 
rect 27 492 30 495 
rect 27 495 30 498 
rect 27 498 30 501 
rect 27 501 30 504 
rect 27 504 30 507 
rect 27 507 30 510 
rect 30 0 33 3 
rect 30 3 33 6 
rect 30 6 33 9 
rect 30 9 33 12 
rect 30 12 33 15 
rect 30 15 33 18 
rect 30 18 33 21 
rect 30 21 33 24 
rect 30 24 33 27 
rect 30 27 33 30 
rect 30 30 33 33 
rect 30 33 33 36 
rect 30 36 33 39 
rect 30 39 33 42 
rect 30 42 33 45 
rect 30 45 33 48 
rect 30 48 33 51 
rect 30 51 33 54 
rect 30 54 33 57 
rect 30 57 33 60 
rect 30 60 33 63 
rect 30 63 33 66 
rect 30 66 33 69 
rect 30 69 33 72 
rect 30 72 33 75 
rect 30 75 33 78 
rect 30 78 33 81 
rect 30 81 33 84 
rect 30 84 33 87 
rect 30 87 33 90 
rect 30 90 33 93 
rect 30 93 33 96 
rect 30 96 33 99 
rect 30 99 33 102 
rect 30 102 33 105 
rect 30 105 33 108 
rect 30 108 33 111 
rect 30 111 33 114 
rect 30 114 33 117 
rect 30 117 33 120 
rect 30 120 33 123 
rect 30 123 33 126 
rect 30 126 33 129 
rect 30 129 33 132 
rect 30 132 33 135 
rect 30 135 33 138 
rect 30 138 33 141 
rect 30 141 33 144 
rect 30 144 33 147 
rect 30 147 33 150 
rect 30 150 33 153 
rect 30 153 33 156 
rect 30 156 33 159 
rect 30 159 33 162 
rect 30 162 33 165 
rect 30 165 33 168 
rect 30 168 33 171 
rect 30 171 33 174 
rect 30 174 33 177 
rect 30 177 33 180 
rect 30 180 33 183 
rect 30 183 33 186 
rect 30 186 33 189 
rect 30 189 33 192 
rect 30 192 33 195 
rect 30 195 33 198 
rect 30 198 33 201 
rect 30 201 33 204 
rect 30 204 33 207 
rect 30 207 33 210 
rect 30 210 33 213 
rect 30 213 33 216 
rect 30 216 33 219 
rect 30 219 33 222 
rect 30 222 33 225 
rect 30 228 33 231 
rect 30 231 33 234 
rect 30 234 33 237 
rect 30 237 33 240 
rect 30 240 33 243 
rect 30 243 33 246 
rect 30 246 33 249 
rect 30 249 33 252 
rect 30 252 33 255 
rect 30 255 33 258 
rect 30 258 33 261 
rect 30 261 33 264 
rect 30 264 33 267 
rect 30 267 33 270 
rect 30 270 33 273 
rect 30 273 33 276 
rect 30 276 33 279 
rect 30 279 33 282 
rect 30 282 33 285 
rect 30 285 33 288 
rect 30 288 33 291 
rect 30 291 33 294 
rect 30 294 33 297 
rect 30 297 33 300 
rect 30 300 33 303 
rect 30 303 33 306 
rect 30 306 33 309 
rect 30 309 33 312 
rect 30 312 33 315 
rect 30 315 33 318 
rect 30 318 33 321 
rect 30 321 33 324 
rect 30 324 33 327 
rect 30 327 33 330 
rect 30 330 33 333 
rect 30 333 33 336 
rect 30 336 33 339 
rect 30 339 33 342 
rect 30 342 33 345 
rect 30 345 33 348 
rect 30 348 33 351 
rect 30 351 33 354 
rect 30 354 33 357 
rect 30 357 33 360 
rect 30 360 33 363 
rect 30 363 33 366 
rect 30 366 33 369 
rect 30 369 33 372 
rect 30 372 33 375 
rect 30 375 33 378 
rect 30 378 33 381 
rect 30 381 33 384 
rect 30 384 33 387 
rect 30 387 33 390 
rect 30 390 33 393 
rect 30 393 33 396 
rect 30 396 33 399 
rect 30 399 33 402 
rect 30 402 33 405 
rect 30 405 33 408 
rect 30 408 33 411 
rect 30 411 33 414 
rect 30 414 33 417 
rect 30 417 33 420 
rect 30 420 33 423 
rect 30 423 33 426 
rect 30 426 33 429 
rect 30 429 33 432 
rect 30 432 33 435 
rect 30 435 33 438 
rect 30 438 33 441 
rect 30 441 33 444 
rect 30 444 33 447 
rect 30 447 33 450 
rect 30 450 33 453 
rect 30 453 33 456 
rect 30 456 33 459 
rect 30 459 33 462 
rect 30 462 33 465 
rect 30 465 33 468 
rect 30 468 33 471 
rect 30 471 33 474 
rect 30 474 33 477 
rect 30 477 33 480 
rect 30 480 33 483 
rect 30 483 33 486 
rect 30 486 33 489 
rect 30 489 33 492 
rect 30 492 33 495 
rect 30 495 33 498 
rect 30 498 33 501 
rect 30 501 33 504 
rect 30 504 33 507 
rect 30 507 33 510 
rect 33 0 36 3 
rect 33 3 36 6 
rect 33 6 36 9 
rect 33 9 36 12 
rect 33 12 36 15 
rect 33 15 36 18 
rect 33 18 36 21 
rect 33 21 36 24 
rect 33 24 36 27 
rect 33 27 36 30 
rect 33 30 36 33 
rect 33 33 36 36 
rect 33 36 36 39 
rect 33 39 36 42 
rect 33 42 36 45 
rect 33 45 36 48 
rect 33 48 36 51 
rect 33 51 36 54 
rect 33 54 36 57 
rect 33 57 36 60 
rect 33 60 36 63 
rect 33 63 36 66 
rect 33 66 36 69 
rect 33 69 36 72 
rect 33 72 36 75 
rect 33 75 36 78 
rect 33 78 36 81 
rect 33 81 36 84 
rect 33 84 36 87 
rect 33 87 36 90 
rect 33 90 36 93 
rect 33 93 36 96 
rect 33 96 36 99 
rect 33 99 36 102 
rect 33 102 36 105 
rect 33 105 36 108 
rect 33 108 36 111 
rect 33 111 36 114 
rect 33 114 36 117 
rect 33 117 36 120 
rect 33 120 36 123 
rect 33 123 36 126 
rect 33 126 36 129 
rect 33 129 36 132 
rect 33 132 36 135 
rect 33 135 36 138 
rect 33 138 36 141 
rect 33 141 36 144 
rect 33 144 36 147 
rect 33 147 36 150 
rect 33 150 36 153 
rect 33 153 36 156 
rect 33 156 36 159 
rect 33 159 36 162 
rect 33 162 36 165 
rect 33 165 36 168 
rect 33 168 36 171 
rect 33 171 36 174 
rect 33 174 36 177 
rect 33 177 36 180 
rect 33 180 36 183 
rect 33 183 36 186 
rect 33 186 36 189 
rect 33 189 36 192 
rect 33 192 36 195 
rect 33 195 36 198 
rect 33 198 36 201 
rect 33 201 36 204 
rect 33 204 36 207 
rect 33 207 36 210 
rect 33 210 36 213 
rect 33 213 36 216 
rect 33 216 36 219 
rect 33 219 36 222 
rect 33 222 36 225 
rect 33 225 36 228 
rect 33 228 36 231 
rect 33 231 36 234 
rect 33 234 36 237 
rect 33 237 36 240 
rect 33 240 36 243 
rect 33 243 36 246 
rect 33 246 36 249 
rect 33 249 36 252 
rect 33 252 36 255 
rect 33 255 36 258 
rect 33 258 36 261 
rect 33 261 36 264 
rect 33 264 36 267 
rect 33 267 36 270 
rect 33 270 36 273 
rect 33 273 36 276 
rect 33 276 36 279 
rect 33 279 36 282 
rect 33 282 36 285 
rect 33 285 36 288 
rect 33 288 36 291 
rect 33 291 36 294 
rect 33 294 36 297 
rect 33 297 36 300 
rect 33 300 36 303 
rect 33 303 36 306 
rect 33 306 36 309 
rect 33 309 36 312 
rect 33 312 36 315 
rect 33 315 36 318 
rect 33 318 36 321 
rect 33 321 36 324 
rect 33 324 36 327 
rect 33 327 36 330 
rect 33 330 36 333 
rect 33 333 36 336 
rect 33 336 36 339 
rect 33 339 36 342 
rect 33 342 36 345 
rect 33 345 36 348 
rect 33 348 36 351 
rect 33 351 36 354 
rect 33 354 36 357 
rect 33 357 36 360 
rect 33 360 36 363 
rect 33 363 36 366 
rect 33 366 36 369 
rect 33 369 36 372 
rect 33 372 36 375 
rect 33 375 36 378 
rect 33 378 36 381 
rect 33 381 36 384 
rect 33 384 36 387 
rect 33 387 36 390 
rect 33 390 36 393 
rect 33 393 36 396 
rect 33 396 36 399 
rect 33 399 36 402 
rect 33 402 36 405 
rect 33 405 36 408 
rect 33 408 36 411 
rect 33 411 36 414 
rect 33 414 36 417 
rect 33 417 36 420 
rect 33 420 36 423 
rect 33 423 36 426 
rect 33 426 36 429 
rect 33 429 36 432 
rect 33 432 36 435 
rect 33 435 36 438 
rect 33 438 36 441 
rect 33 441 36 444 
rect 33 444 36 447 
rect 33 447 36 450 
rect 33 450 36 453 
rect 33 453 36 456 
rect 33 456 36 459 
rect 33 459 36 462 
rect 33 462 36 465 
rect 33 465 36 468 
rect 33 468 36 471 
rect 33 471 36 474 
rect 33 474 36 477 
rect 33 477 36 480 
rect 33 480 36 483 
rect 33 483 36 486 
rect 33 486 36 489 
rect 33 489 36 492 
rect 33 492 36 495 
rect 33 495 36 498 
rect 33 498 36 501 
rect 33 501 36 504 
rect 33 504 36 507 
rect 33 507 36 510 
rect 36 0 39 3 
rect 36 3 39 6 
rect 36 6 39 9 
rect 36 9 39 12 
rect 36 12 39 15 
rect 36 15 39 18 
rect 36 18 39 21 
rect 36 21 39 24 
rect 36 24 39 27 
rect 36 27 39 30 
rect 36 30 39 33 
rect 36 33 39 36 
rect 36 36 39 39 
rect 36 39 39 42 
rect 36 42 39 45 
rect 36 45 39 48 
rect 36 48 39 51 
rect 36 51 39 54 
rect 36 54 39 57 
rect 36 57 39 60 
rect 36 60 39 63 
rect 36 63 39 66 
rect 36 66 39 69 
rect 36 69 39 72 
rect 36 72 39 75 
rect 36 75 39 78 
rect 36 78 39 81 
rect 36 81 39 84 
rect 36 84 39 87 
rect 36 87 39 90 
rect 36 90 39 93 
rect 36 93 39 96 
rect 36 96 39 99 
rect 36 99 39 102 
rect 36 102 39 105 
rect 36 105 39 108 
rect 36 108 39 111 
rect 36 111 39 114 
rect 36 114 39 117 
rect 36 117 39 120 
rect 36 120 39 123 
rect 36 123 39 126 
rect 36 126 39 129 
rect 36 129 39 132 
rect 36 132 39 135 
rect 36 135 39 138 
rect 36 138 39 141 
rect 36 141 39 144 
rect 36 144 39 147 
rect 36 147 39 150 
rect 36 150 39 153 
rect 36 153 39 156 
rect 36 156 39 159 
rect 36 159 39 162 
rect 36 162 39 165 
rect 36 165 39 168 
rect 36 168 39 171 
rect 36 171 39 174 
rect 36 174 39 177 
rect 36 177 39 180 
rect 36 180 39 183 
rect 36 183 39 186 
rect 36 186 39 189 
rect 36 189 39 192 
rect 36 192 39 195 
rect 36 195 39 198 
rect 36 198 39 201 
rect 36 201 39 204 
rect 36 204 39 207 
rect 36 207 39 210 
rect 36 210 39 213 
rect 36 213 39 216 
rect 36 216 39 219 
rect 36 219 39 222 
rect 36 222 39 225 
rect 36 225 39 228 
rect 36 228 39 231 
rect 36 231 39 234 
rect 36 234 39 237 
rect 36 237 39 240 
rect 36 240 39 243 
rect 36 243 39 246 
rect 36 246 39 249 
rect 36 249 39 252 
rect 36 252 39 255 
rect 36 255 39 258 
rect 36 258 39 261 
rect 36 261 39 264 
rect 36 264 39 267 
rect 36 267 39 270 
rect 36 270 39 273 
rect 36 273 39 276 
rect 36 276 39 279 
rect 36 279 39 282 
rect 36 282 39 285 
rect 36 285 39 288 
rect 36 288 39 291 
rect 36 291 39 294 
rect 36 294 39 297 
rect 36 297 39 300 
rect 36 300 39 303 
rect 36 303 39 306 
rect 36 306 39 309 
rect 36 309 39 312 
rect 36 312 39 315 
rect 36 315 39 318 
rect 36 318 39 321 
rect 36 321 39 324 
rect 36 324 39 327 
rect 36 327 39 330 
rect 36 330 39 333 
rect 36 333 39 336 
rect 36 336 39 339 
rect 36 339 39 342 
rect 36 342 39 345 
rect 36 345 39 348 
rect 36 348 39 351 
rect 36 351 39 354 
rect 36 354 39 357 
rect 36 357 39 360 
rect 36 360 39 363 
rect 36 363 39 366 
rect 36 366 39 369 
rect 36 369 39 372 
rect 36 372 39 375 
rect 36 375 39 378 
rect 36 378 39 381 
rect 36 381 39 384 
rect 36 384 39 387 
rect 36 387 39 390 
rect 36 390 39 393 
rect 36 393 39 396 
rect 36 396 39 399 
rect 36 399 39 402 
rect 36 402 39 405 
rect 36 405 39 408 
rect 36 408 39 411 
rect 36 411 39 414 
rect 36 414 39 417 
rect 36 417 39 420 
rect 36 420 39 423 
rect 36 423 39 426 
rect 36 426 39 429 
rect 36 429 39 432 
rect 36 432 39 435 
rect 36 435 39 438 
rect 36 438 39 441 
rect 36 441 39 444 
rect 36 444 39 447 
rect 36 447 39 450 
rect 36 450 39 453 
rect 36 453 39 456 
rect 36 456 39 459 
rect 36 459 39 462 
rect 36 462 39 465 
rect 36 465 39 468 
rect 36 468 39 471 
rect 36 471 39 474 
rect 36 474 39 477 
rect 36 477 39 480 
rect 36 480 39 483 
rect 36 483 39 486 
rect 36 486 39 489 
rect 36 489 39 492 
rect 36 492 39 495 
rect 36 495 39 498 
rect 36 498 39 501 
rect 36 501 39 504 
rect 36 504 39 507 
rect 36 507 39 510 
rect 39 0 42 3 
rect 39 3 42 6 
rect 39 6 42 9 
rect 39 9 42 12 
rect 39 12 42 15 
rect 39 15 42 18 
rect 39 18 42 21 
rect 39 21 42 24 
rect 39 24 42 27 
rect 39 27 42 30 
rect 39 30 42 33 
rect 39 33 42 36 
rect 39 36 42 39 
rect 39 39 42 42 
rect 39 42 42 45 
rect 39 45 42 48 
rect 39 48 42 51 
rect 39 51 42 54 
rect 39 54 42 57 
rect 39 57 42 60 
rect 39 60 42 63 
rect 39 63 42 66 
rect 39 66 42 69 
rect 39 69 42 72 
rect 39 72 42 75 
rect 39 75 42 78 
rect 39 78 42 81 
rect 39 81 42 84 
rect 39 84 42 87 
rect 39 87 42 90 
rect 39 90 42 93 
rect 39 93 42 96 
rect 39 96 42 99 
rect 39 99 42 102 
rect 39 102 42 105 
rect 39 105 42 108 
rect 39 108 42 111 
rect 39 111 42 114 
rect 39 114 42 117 
rect 39 117 42 120 
rect 39 120 42 123 
rect 39 123 42 126 
rect 39 126 42 129 
rect 39 129 42 132 
rect 39 132 42 135 
rect 39 135 42 138 
rect 39 138 42 141 
rect 39 141 42 144 
rect 39 144 42 147 
rect 39 147 42 150 
rect 39 150 42 153 
rect 39 153 42 156 
rect 39 156 42 159 
rect 39 159 42 162 
rect 39 162 42 165 
rect 39 165 42 168 
rect 39 168 42 171 
rect 39 171 42 174 
rect 39 174 42 177 
rect 39 177 42 180 
rect 39 180 42 183 
rect 39 183 42 186 
rect 39 186 42 189 
rect 39 189 42 192 
rect 39 192 42 195 
rect 39 195 42 198 
rect 39 198 42 201 
rect 39 201 42 204 
rect 39 204 42 207 
rect 39 207 42 210 
rect 39 210 42 213 
rect 39 213 42 216 
rect 39 216 42 219 
rect 39 219 42 222 
rect 39 222 42 225 
rect 39 225 42 228 
rect 39 228 42 231 
rect 39 231 42 234 
rect 39 234 42 237 
rect 39 237 42 240 
rect 39 240 42 243 
rect 39 243 42 246 
rect 39 246 42 249 
rect 39 249 42 252 
rect 39 252 42 255 
rect 39 255 42 258 
rect 39 258 42 261 
rect 39 261 42 264 
rect 39 264 42 267 
rect 39 267 42 270 
rect 39 270 42 273 
rect 39 273 42 276 
rect 39 276 42 279 
rect 39 279 42 282 
rect 39 282 42 285 
rect 39 285 42 288 
rect 39 288 42 291 
rect 39 291 42 294 
rect 39 294 42 297 
rect 39 297 42 300 
rect 39 300 42 303 
rect 39 303 42 306 
rect 39 306 42 309 
rect 39 309 42 312 
rect 39 312 42 315 
rect 39 315 42 318 
rect 39 318 42 321 
rect 39 321 42 324 
rect 39 324 42 327 
rect 39 327 42 330 
rect 39 330 42 333 
rect 39 333 42 336 
rect 39 336 42 339 
rect 39 339 42 342 
rect 39 342 42 345 
rect 39 345 42 348 
rect 39 348 42 351 
rect 39 351 42 354 
rect 39 354 42 357 
rect 39 357 42 360 
rect 39 360 42 363 
rect 39 363 42 366 
rect 39 366 42 369 
rect 39 369 42 372 
rect 39 372 42 375 
rect 39 375 42 378 
rect 39 378 42 381 
rect 39 381 42 384 
rect 39 384 42 387 
rect 39 387 42 390 
rect 39 390 42 393 
rect 39 393 42 396 
rect 39 396 42 399 
rect 39 399 42 402 
rect 39 402 42 405 
rect 39 405 42 408 
rect 39 408 42 411 
rect 39 411 42 414 
rect 39 414 42 417 
rect 39 417 42 420 
rect 39 420 42 423 
rect 39 423 42 426 
rect 39 426 42 429 
rect 39 429 42 432 
rect 39 432 42 435 
rect 39 435 42 438 
rect 39 438 42 441 
rect 39 441 42 444 
rect 39 444 42 447 
rect 39 447 42 450 
rect 39 450 42 453 
rect 39 453 42 456 
rect 39 456 42 459 
rect 39 459 42 462 
rect 39 462 42 465 
rect 39 465 42 468 
rect 39 468 42 471 
rect 39 471 42 474 
rect 39 474 42 477 
rect 39 477 42 480 
rect 39 480 42 483 
rect 39 483 42 486 
rect 39 486 42 489 
rect 39 489 42 492 
rect 39 492 42 495 
rect 39 495 42 498 
rect 39 498 42 501 
rect 39 501 42 504 
rect 39 504 42 507 
rect 39 507 42 510 
rect 42 0 45 3 
rect 42 3 45 6 
rect 42 6 45 9 
rect 42 9 45 12 
rect 42 12 45 15 
rect 42 15 45 18 
rect 42 18 45 21 
rect 42 21 45 24 
rect 42 24 45 27 
rect 42 27 45 30 
rect 42 30 45 33 
rect 42 33 45 36 
rect 42 36 45 39 
rect 42 39 45 42 
rect 42 42 45 45 
rect 42 45 45 48 
rect 42 48 45 51 
rect 42 51 45 54 
rect 42 54 45 57 
rect 42 57 45 60 
rect 42 60 45 63 
rect 42 63 45 66 
rect 42 66 45 69 
rect 42 69 45 72 
rect 42 72 45 75 
rect 42 75 45 78 
rect 42 78 45 81 
rect 42 81 45 84 
rect 42 84 45 87 
rect 42 87 45 90 
rect 42 90 45 93 
rect 42 93 45 96 
rect 42 96 45 99 
rect 42 99 45 102 
rect 42 102 45 105 
rect 42 105 45 108 
rect 42 108 45 111 
rect 42 111 45 114 
rect 42 114 45 117 
rect 42 117 45 120 
rect 42 120 45 123 
rect 42 123 45 126 
rect 42 126 45 129 
rect 42 129 45 132 
rect 42 132 45 135 
rect 42 135 45 138 
rect 42 138 45 141 
rect 42 141 45 144 
rect 42 144 45 147 
rect 42 147 45 150 
rect 42 150 45 153 
rect 42 153 45 156 
rect 42 156 45 159 
rect 42 159 45 162 
rect 42 162 45 165 
rect 42 165 45 168 
rect 42 168 45 171 
rect 42 171 45 174 
rect 42 174 45 177 
rect 42 177 45 180 
rect 42 180 45 183 
rect 42 183 45 186 
rect 42 186 45 189 
rect 42 189 45 192 
rect 42 192 45 195 
rect 42 195 45 198 
rect 42 198 45 201 
rect 42 201 45 204 
rect 42 204 45 207 
rect 42 207 45 210 
rect 42 210 45 213 
rect 42 213 45 216 
rect 42 216 45 219 
rect 42 219 45 222 
rect 42 222 45 225 
rect 42 225 45 228 
rect 42 228 45 231 
rect 42 231 45 234 
rect 42 234 45 237 
rect 42 237 45 240 
rect 42 240 45 243 
rect 42 243 45 246 
rect 42 246 45 249 
rect 42 249 45 252 
rect 42 252 45 255 
rect 42 255 45 258 
rect 42 258 45 261 
rect 42 261 45 264 
rect 42 264 45 267 
rect 42 267 45 270 
rect 42 270 45 273 
rect 42 273 45 276 
rect 42 276 45 279 
rect 42 279 45 282 
rect 42 282 45 285 
rect 42 285 45 288 
rect 42 288 45 291 
rect 42 291 45 294 
rect 42 294 45 297 
rect 42 297 45 300 
rect 42 300 45 303 
rect 42 303 45 306 
rect 42 306 45 309 
rect 42 309 45 312 
rect 42 312 45 315 
rect 42 315 45 318 
rect 42 318 45 321 
rect 42 321 45 324 
rect 42 324 45 327 
rect 42 327 45 330 
rect 42 330 45 333 
rect 42 333 45 336 
rect 42 336 45 339 
rect 42 339 45 342 
rect 42 342 45 345 
rect 42 345 45 348 
rect 42 348 45 351 
rect 42 351 45 354 
rect 42 354 45 357 
rect 42 357 45 360 
rect 42 360 45 363 
rect 42 363 45 366 
rect 42 366 45 369 
rect 42 369 45 372 
rect 42 372 45 375 
rect 42 375 45 378 
rect 42 378 45 381 
rect 42 381 45 384 
rect 42 384 45 387 
rect 42 387 45 390 
rect 42 390 45 393 
rect 42 393 45 396 
rect 42 396 45 399 
rect 42 399 45 402 
rect 42 402 45 405 
rect 42 405 45 408 
rect 42 408 45 411 
rect 42 411 45 414 
rect 42 414 45 417 
rect 42 417 45 420 
rect 42 420 45 423 
rect 42 423 45 426 
rect 42 426 45 429 
rect 42 429 45 432 
rect 42 432 45 435 
rect 42 435 45 438 
rect 42 438 45 441 
rect 42 441 45 444 
rect 42 444 45 447 
rect 42 447 45 450 
rect 42 450 45 453 
rect 42 453 45 456 
rect 42 456 45 459 
rect 42 459 45 462 
rect 42 462 45 465 
rect 42 465 45 468 
rect 42 468 45 471 
rect 42 471 45 474 
rect 42 474 45 477 
rect 42 477 45 480 
rect 42 480 45 483 
rect 42 483 45 486 
rect 42 486 45 489 
rect 42 489 45 492 
rect 42 492 45 495 
rect 42 495 45 498 
rect 42 498 45 501 
rect 42 501 45 504 
rect 42 504 45 507 
rect 42 507 45 510 
rect 45 0 48 3 
rect 45 3 48 6 
rect 45 6 48 9 
rect 45 9 48 12 
rect 45 12 48 15 
rect 45 15 48 18 
rect 45 18 48 21 
rect 45 21 48 24 
rect 45 24 48 27 
rect 45 27 48 30 
rect 45 30 48 33 
rect 45 33 48 36 
rect 45 36 48 39 
rect 45 39 48 42 
rect 45 42 48 45 
rect 45 45 48 48 
rect 45 48 48 51 
rect 45 51 48 54 
rect 45 54 48 57 
rect 45 57 48 60 
rect 45 60 48 63 
rect 45 63 48 66 
rect 45 66 48 69 
rect 45 69 48 72 
rect 45 72 48 75 
rect 45 75 48 78 
rect 45 78 48 81 
rect 45 81 48 84 
rect 45 84 48 87 
rect 45 87 48 90 
rect 45 90 48 93 
rect 45 93 48 96 
rect 45 96 48 99 
rect 45 99 48 102 
rect 45 102 48 105 
rect 45 105 48 108 
rect 45 108 48 111 
rect 45 111 48 114 
rect 45 114 48 117 
rect 45 117 48 120 
rect 45 120 48 123 
rect 45 123 48 126 
rect 45 126 48 129 
rect 45 129 48 132 
rect 45 132 48 135 
rect 45 135 48 138 
rect 45 138 48 141 
rect 45 141 48 144 
rect 45 144 48 147 
rect 45 147 48 150 
rect 45 150 48 153 
rect 45 153 48 156 
rect 45 156 48 159 
rect 45 159 48 162 
rect 45 162 48 165 
rect 45 165 48 168 
rect 45 168 48 171 
rect 45 171 48 174 
rect 45 174 48 177 
rect 45 177 48 180 
rect 45 180 48 183 
rect 45 183 48 186 
rect 45 186 48 189 
rect 45 189 48 192 
rect 45 192 48 195 
rect 45 195 48 198 
rect 45 198 48 201 
rect 45 201 48 204 
rect 45 204 48 207 
rect 45 207 48 210 
rect 45 210 48 213 
rect 45 213 48 216 
rect 45 216 48 219 
rect 45 219 48 222 
rect 45 222 48 225 
rect 45 225 48 228 
rect 45 228 48 231 
rect 45 231 48 234 
rect 45 234 48 237 
rect 45 237 48 240 
rect 45 240 48 243 
rect 45 243 48 246 
rect 45 246 48 249 
rect 45 249 48 252 
rect 45 252 48 255 
rect 45 255 48 258 
rect 45 258 48 261 
rect 45 261 48 264 
rect 45 264 48 267 
rect 45 267 48 270 
rect 45 270 48 273 
rect 45 273 48 276 
rect 45 276 48 279 
rect 45 279 48 282 
rect 45 282 48 285 
rect 45 285 48 288 
rect 45 288 48 291 
rect 45 291 48 294 
rect 45 294 48 297 
rect 45 297 48 300 
rect 45 300 48 303 
rect 45 303 48 306 
rect 45 306 48 309 
rect 45 309 48 312 
rect 45 312 48 315 
rect 45 315 48 318 
rect 45 318 48 321 
rect 45 321 48 324 
rect 45 324 48 327 
rect 45 327 48 330 
rect 45 330 48 333 
rect 45 333 48 336 
rect 45 336 48 339 
rect 45 339 48 342 
rect 45 342 48 345 
rect 45 345 48 348 
rect 45 348 48 351 
rect 45 351 48 354 
rect 45 354 48 357 
rect 45 357 48 360 
rect 45 360 48 363 
rect 45 363 48 366 
rect 45 366 48 369 
rect 45 369 48 372 
rect 45 372 48 375 
rect 45 375 48 378 
rect 45 378 48 381 
rect 45 381 48 384 
rect 45 384 48 387 
rect 45 387 48 390 
rect 45 390 48 393 
rect 45 393 48 396 
rect 45 396 48 399 
rect 45 399 48 402 
rect 45 402 48 405 
rect 45 405 48 408 
rect 45 408 48 411 
rect 45 411 48 414 
rect 45 414 48 417 
rect 45 417 48 420 
rect 45 420 48 423 
rect 45 423 48 426 
rect 45 426 48 429 
rect 45 429 48 432 
rect 45 432 48 435 
rect 45 435 48 438 
rect 45 438 48 441 
rect 45 441 48 444 
rect 45 444 48 447 
rect 45 447 48 450 
rect 45 450 48 453 
rect 45 453 48 456 
rect 45 456 48 459 
rect 45 459 48 462 
rect 45 462 48 465 
rect 45 465 48 468 
rect 45 468 48 471 
rect 45 471 48 474 
rect 45 474 48 477 
rect 45 477 48 480 
rect 45 480 48 483 
rect 45 483 48 486 
rect 45 486 48 489 
rect 45 489 48 492 
rect 45 492 48 495 
rect 45 495 48 498 
rect 45 498 48 501 
rect 45 501 48 504 
rect 45 504 48 507 
rect 45 507 48 510 
rect 48 0 51 3 
rect 48 3 51 6 
rect 48 6 51 9 
rect 48 9 51 12 
rect 48 12 51 15 
rect 48 15 51 18 
rect 48 18 51 21 
rect 48 21 51 24 
rect 48 24 51 27 
rect 48 27 51 30 
rect 48 30 51 33 
rect 48 33 51 36 
rect 48 36 51 39 
rect 48 39 51 42 
rect 48 42 51 45 
rect 48 45 51 48 
rect 48 48 51 51 
rect 48 51 51 54 
rect 48 54 51 57 
rect 48 57 51 60 
rect 48 60 51 63 
rect 48 63 51 66 
rect 48 66 51 69 
rect 48 69 51 72 
rect 48 72 51 75 
rect 48 75 51 78 
rect 48 78 51 81 
rect 48 81 51 84 
rect 48 84 51 87 
rect 48 87 51 90 
rect 48 90 51 93 
rect 48 93 51 96 
rect 48 96 51 99 
rect 48 99 51 102 
rect 48 102 51 105 
rect 48 105 51 108 
rect 48 108 51 111 
rect 48 111 51 114 
rect 48 114 51 117 
rect 48 117 51 120 
rect 48 120 51 123 
rect 48 123 51 126 
rect 48 126 51 129 
rect 48 129 51 132 
rect 48 132 51 135 
rect 48 135 51 138 
rect 48 138 51 141 
rect 48 141 51 144 
rect 48 144 51 147 
rect 48 147 51 150 
rect 48 150 51 153 
rect 48 153 51 156 
rect 48 156 51 159 
rect 48 159 51 162 
rect 48 162 51 165 
rect 48 165 51 168 
rect 48 168 51 171 
rect 48 171 51 174 
rect 48 174 51 177 
rect 48 177 51 180 
rect 48 180 51 183 
rect 48 183 51 186 
rect 48 186 51 189 
rect 48 189 51 192 
rect 48 192 51 195 
rect 48 195 51 198 
rect 48 198 51 201 
rect 48 201 51 204 
rect 48 204 51 207 
rect 48 207 51 210 
rect 48 210 51 213 
rect 48 213 51 216 
rect 48 216 51 219 
rect 48 219 51 222 
rect 48 222 51 225 
rect 48 225 51 228 
rect 48 228 51 231 
rect 48 231 51 234 
rect 48 234 51 237 
rect 48 237 51 240 
rect 48 240 51 243 
rect 48 243 51 246 
rect 48 246 51 249 
rect 48 249 51 252 
rect 48 252 51 255 
rect 48 255 51 258 
rect 48 258 51 261 
rect 48 261 51 264 
rect 48 264 51 267 
rect 48 267 51 270 
rect 48 270 51 273 
rect 48 273 51 276 
rect 48 276 51 279 
rect 48 279 51 282 
rect 48 282 51 285 
rect 48 285 51 288 
rect 48 288 51 291 
rect 48 291 51 294 
rect 48 294 51 297 
rect 48 297 51 300 
rect 48 300 51 303 
rect 48 303 51 306 
rect 48 306 51 309 
rect 48 309 51 312 
rect 48 312 51 315 
rect 48 315 51 318 
rect 48 318 51 321 
rect 48 321 51 324 
rect 48 324 51 327 
rect 48 327 51 330 
rect 48 330 51 333 
rect 48 333 51 336 
rect 48 336 51 339 
rect 48 339 51 342 
rect 48 342 51 345 
rect 48 345 51 348 
rect 48 348 51 351 
rect 48 351 51 354 
rect 48 354 51 357 
rect 48 357 51 360 
rect 48 360 51 363 
rect 48 363 51 366 
rect 48 366 51 369 
rect 48 369 51 372 
rect 48 372 51 375 
rect 48 375 51 378 
rect 48 378 51 381 
rect 48 381 51 384 
rect 48 384 51 387 
rect 48 387 51 390 
rect 48 390 51 393 
rect 48 393 51 396 
rect 48 396 51 399 
rect 48 399 51 402 
rect 48 402 51 405 
rect 48 405 51 408 
rect 48 408 51 411 
rect 48 411 51 414 
rect 48 414 51 417 
rect 48 417 51 420 
rect 48 420 51 423 
rect 48 423 51 426 
rect 48 426 51 429 
rect 48 429 51 432 
rect 48 432 51 435 
rect 48 435 51 438 
rect 48 438 51 441 
rect 48 441 51 444 
rect 48 444 51 447 
rect 48 447 51 450 
rect 48 450 51 453 
rect 48 453 51 456 
rect 48 456 51 459 
rect 48 459 51 462 
rect 48 462 51 465 
rect 48 465 51 468 
rect 48 468 51 471 
rect 48 471 51 474 
rect 48 474 51 477 
rect 48 477 51 480 
rect 48 480 51 483 
rect 48 483 51 486 
rect 48 486 51 489 
rect 48 489 51 492 
rect 48 492 51 495 
rect 48 495 51 498 
rect 48 498 51 501 
rect 48 501 51 504 
rect 48 504 51 507 
rect 48 507 51 510 
rect 51 0 54 3 
rect 51 3 54 6 
rect 51 6 54 9 
rect 51 9 54 12 
rect 51 12 54 15 
rect 51 15 54 18 
rect 51 18 54 21 
rect 51 21 54 24 
rect 51 24 54 27 
rect 51 27 54 30 
rect 51 30 54 33 
rect 51 33 54 36 
rect 51 36 54 39 
rect 51 39 54 42 
rect 51 42 54 45 
rect 51 45 54 48 
rect 51 48 54 51 
rect 51 51 54 54 
rect 51 54 54 57 
rect 51 57 54 60 
rect 51 60 54 63 
rect 51 63 54 66 
rect 51 66 54 69 
rect 51 69 54 72 
rect 51 72 54 75 
rect 51 75 54 78 
rect 51 78 54 81 
rect 51 81 54 84 
rect 51 84 54 87 
rect 51 87 54 90 
rect 51 90 54 93 
rect 51 93 54 96 
rect 51 96 54 99 
rect 51 99 54 102 
rect 51 102 54 105 
rect 51 105 54 108 
rect 51 108 54 111 
rect 51 111 54 114 
rect 51 114 54 117 
rect 51 117 54 120 
rect 51 120 54 123 
rect 51 123 54 126 
rect 51 126 54 129 
rect 51 129 54 132 
rect 51 132 54 135 
rect 51 135 54 138 
rect 51 138 54 141 
rect 51 141 54 144 
rect 51 144 54 147 
rect 51 147 54 150 
rect 51 150 54 153 
rect 51 153 54 156 
rect 51 156 54 159 
rect 51 159 54 162 
rect 51 162 54 165 
rect 51 165 54 168 
rect 51 168 54 171 
rect 51 171 54 174 
rect 51 174 54 177 
rect 51 177 54 180 
rect 51 180 54 183 
rect 51 183 54 186 
rect 51 186 54 189 
rect 51 189 54 192 
rect 51 192 54 195 
rect 51 195 54 198 
rect 51 198 54 201 
rect 51 201 54 204 
rect 51 204 54 207 
rect 51 207 54 210 
rect 51 210 54 213 
rect 51 213 54 216 
rect 51 216 54 219 
rect 51 219 54 222 
rect 51 222 54 225 
rect 51 225 54 228 
rect 51 228 54 231 
rect 51 231 54 234 
rect 51 234 54 237 
rect 51 237 54 240 
rect 51 240 54 243 
rect 51 243 54 246 
rect 51 246 54 249 
rect 51 249 54 252 
rect 51 252 54 255 
rect 51 255 54 258 
rect 51 258 54 261 
rect 51 261 54 264 
rect 51 264 54 267 
rect 51 267 54 270 
rect 51 270 54 273 
rect 51 273 54 276 
rect 51 276 54 279 
rect 51 279 54 282 
rect 51 282 54 285 
rect 51 285 54 288 
rect 51 288 54 291 
rect 51 291 54 294 
rect 51 294 54 297 
rect 51 297 54 300 
rect 51 300 54 303 
rect 51 303 54 306 
rect 51 306 54 309 
rect 51 309 54 312 
rect 51 312 54 315 
rect 51 315 54 318 
rect 51 318 54 321 
rect 51 321 54 324 
rect 51 324 54 327 
rect 51 327 54 330 
rect 51 330 54 333 
rect 51 333 54 336 
rect 51 336 54 339 
rect 51 339 54 342 
rect 51 342 54 345 
rect 51 345 54 348 
rect 51 348 54 351 
rect 51 351 54 354 
rect 51 354 54 357 
rect 51 357 54 360 
rect 51 360 54 363 
rect 51 363 54 366 
rect 51 366 54 369 
rect 51 369 54 372 
rect 51 372 54 375 
rect 51 375 54 378 
rect 51 378 54 381 
rect 51 381 54 384 
rect 51 384 54 387 
rect 51 387 54 390 
rect 51 390 54 393 
rect 51 393 54 396 
rect 51 396 54 399 
rect 51 399 54 402 
rect 51 402 54 405 
rect 51 405 54 408 
rect 51 408 54 411 
rect 51 411 54 414 
rect 51 414 54 417 
rect 51 417 54 420 
rect 51 420 54 423 
rect 51 423 54 426 
rect 51 426 54 429 
rect 51 429 54 432 
rect 51 432 54 435 
rect 51 435 54 438 
rect 51 438 54 441 
rect 51 441 54 444 
rect 51 444 54 447 
rect 51 447 54 450 
rect 51 450 54 453 
rect 51 453 54 456 
rect 51 456 54 459 
rect 51 459 54 462 
rect 51 462 54 465 
rect 51 465 54 468 
rect 51 468 54 471 
rect 51 471 54 474 
rect 51 474 54 477 
rect 51 477 54 480 
rect 51 480 54 483 
rect 51 483 54 486 
rect 51 486 54 489 
rect 51 489 54 492 
rect 51 492 54 495 
rect 51 495 54 498 
rect 51 498 54 501 
rect 51 501 54 504 
rect 51 504 54 507 
rect 51 507 54 510 
rect 54 0 57 3 
rect 54 3 57 6 
rect 54 6 57 9 
rect 54 9 57 12 
rect 54 12 57 15 
rect 54 15 57 18 
rect 54 18 57 21 
rect 54 21 57 24 
rect 54 24 57 27 
rect 54 27 57 30 
rect 54 30 57 33 
rect 54 33 57 36 
rect 54 36 57 39 
rect 54 39 57 42 
rect 54 42 57 45 
rect 54 45 57 48 
rect 54 48 57 51 
rect 54 51 57 54 
rect 54 54 57 57 
rect 54 57 57 60 
rect 54 60 57 63 
rect 54 63 57 66 
rect 54 66 57 69 
rect 54 69 57 72 
rect 54 72 57 75 
rect 54 75 57 78 
rect 54 78 57 81 
rect 54 81 57 84 
rect 54 84 57 87 
rect 54 87 57 90 
rect 54 90 57 93 
rect 54 93 57 96 
rect 54 96 57 99 
rect 54 99 57 102 
rect 54 102 57 105 
rect 54 105 57 108 
rect 54 108 57 111 
rect 54 111 57 114 
rect 54 114 57 117 
rect 54 117 57 120 
rect 54 120 57 123 
rect 54 123 57 126 
rect 54 126 57 129 
rect 54 129 57 132 
rect 54 132 57 135 
rect 54 135 57 138 
rect 54 138 57 141 
rect 54 141 57 144 
rect 54 144 57 147 
rect 54 147 57 150 
rect 54 150 57 153 
rect 54 153 57 156 
rect 54 156 57 159 
rect 54 159 57 162 
rect 54 162 57 165 
rect 54 165 57 168 
rect 54 168 57 171 
rect 54 171 57 174 
rect 54 174 57 177 
rect 54 177 57 180 
rect 54 180 57 183 
rect 54 183 57 186 
rect 54 186 57 189 
rect 54 189 57 192 
rect 54 192 57 195 
rect 54 195 57 198 
rect 54 198 57 201 
rect 54 201 57 204 
rect 54 204 57 207 
rect 54 207 57 210 
rect 54 210 57 213 
rect 54 213 57 216 
rect 54 216 57 219 
rect 54 219 57 222 
rect 54 222 57 225 
rect 54 225 57 228 
rect 54 228 57 231 
rect 54 231 57 234 
rect 54 234 57 237 
rect 54 237 57 240 
rect 54 240 57 243 
rect 54 243 57 246 
rect 54 246 57 249 
rect 54 249 57 252 
rect 54 252 57 255 
rect 54 255 57 258 
rect 54 258 57 261 
rect 54 261 57 264 
rect 54 264 57 267 
rect 54 267 57 270 
rect 54 270 57 273 
rect 54 273 57 276 
rect 54 276 57 279 
rect 54 279 57 282 
rect 54 282 57 285 
rect 54 285 57 288 
rect 54 288 57 291 
rect 54 291 57 294 
rect 54 294 57 297 
rect 54 297 57 300 
rect 54 300 57 303 
rect 54 303 57 306 
rect 54 306 57 309 
rect 54 309 57 312 
rect 54 312 57 315 
rect 54 315 57 318 
rect 54 318 57 321 
rect 54 321 57 324 
rect 54 324 57 327 
rect 54 327 57 330 
rect 54 330 57 333 
rect 54 333 57 336 
rect 54 336 57 339 
rect 54 339 57 342 
rect 54 342 57 345 
rect 54 345 57 348 
rect 54 348 57 351 
rect 54 351 57 354 
rect 54 354 57 357 
rect 54 357 57 360 
rect 54 360 57 363 
rect 54 363 57 366 
rect 54 366 57 369 
rect 54 369 57 372 
rect 54 372 57 375 
rect 54 375 57 378 
rect 54 378 57 381 
rect 54 381 57 384 
rect 54 384 57 387 
rect 54 387 57 390 
rect 54 390 57 393 
rect 54 393 57 396 
rect 54 396 57 399 
rect 54 399 57 402 
rect 54 402 57 405 
rect 54 405 57 408 
rect 54 408 57 411 
rect 54 411 57 414 
rect 54 414 57 417 
rect 54 417 57 420 
rect 54 420 57 423 
rect 54 423 57 426 
rect 54 426 57 429 
rect 54 429 57 432 
rect 54 432 57 435 
rect 54 435 57 438 
rect 54 438 57 441 
rect 54 441 57 444 
rect 54 444 57 447 
rect 54 447 57 450 
rect 54 450 57 453 
rect 54 453 57 456 
rect 54 456 57 459 
rect 54 459 57 462 
rect 54 462 57 465 
rect 54 465 57 468 
rect 54 468 57 471 
rect 54 471 57 474 
rect 54 474 57 477 
rect 54 477 57 480 
rect 54 480 57 483 
rect 54 483 57 486 
rect 54 486 57 489 
rect 54 489 57 492 
rect 54 492 57 495 
rect 54 495 57 498 
rect 54 498 57 501 
rect 54 501 57 504 
rect 54 504 57 507 
rect 54 507 57 510 
rect 57 0 60 3 
rect 57 3 60 6 
rect 57 6 60 9 
rect 57 9 60 12 
rect 57 12 60 15 
rect 57 15 60 18 
rect 57 18 60 21 
rect 57 21 60 24 
rect 57 24 60 27 
rect 57 27 60 30 
rect 57 30 60 33 
rect 57 33 60 36 
rect 57 36 60 39 
rect 57 39 60 42 
rect 57 42 60 45 
rect 57 45 60 48 
rect 57 48 60 51 
rect 57 51 60 54 
rect 57 54 60 57 
rect 57 57 60 60 
rect 57 60 60 63 
rect 57 63 60 66 
rect 57 66 60 69 
rect 57 69 60 72 
rect 57 72 60 75 
rect 57 75 60 78 
rect 57 78 60 81 
rect 57 81 60 84 
rect 57 84 60 87 
rect 57 87 60 90 
rect 57 90 60 93 
rect 57 93 60 96 
rect 57 96 60 99 
rect 57 99 60 102 
rect 57 102 60 105 
rect 57 105 60 108 
rect 57 108 60 111 
rect 57 111 60 114 
rect 57 114 60 117 
rect 57 117 60 120 
rect 57 120 60 123 
rect 57 123 60 126 
rect 57 126 60 129 
rect 57 129 60 132 
rect 57 132 60 135 
rect 57 135 60 138 
rect 57 138 60 141 
rect 57 141 60 144 
rect 57 144 60 147 
rect 57 147 60 150 
rect 57 150 60 153 
rect 57 153 60 156 
rect 57 156 60 159 
rect 57 159 60 162 
rect 57 162 60 165 
rect 57 165 60 168 
rect 57 168 60 171 
rect 57 171 60 174 
rect 57 174 60 177 
rect 57 177 60 180 
rect 57 180 60 183 
rect 57 183 60 186 
rect 57 186 60 189 
rect 57 189 60 192 
rect 57 192 60 195 
rect 57 195 60 198 
rect 57 198 60 201 
rect 57 201 60 204 
rect 57 204 60 207 
rect 57 207 60 210 
rect 57 210 60 213 
rect 57 213 60 216 
rect 57 216 60 219 
rect 57 219 60 222 
rect 57 222 60 225 
rect 57 225 60 228 
rect 57 228 60 231 
rect 57 231 60 234 
rect 57 234 60 237 
rect 57 237 60 240 
rect 57 240 60 243 
rect 57 243 60 246 
rect 57 246 60 249 
rect 57 249 60 252 
rect 57 252 60 255 
rect 57 255 60 258 
rect 57 258 60 261 
rect 57 261 60 264 
rect 57 264 60 267 
rect 57 267 60 270 
rect 57 270 60 273 
rect 57 273 60 276 
rect 57 276 60 279 
rect 57 279 60 282 
rect 57 282 60 285 
rect 57 285 60 288 
rect 57 288 60 291 
rect 57 291 60 294 
rect 57 294 60 297 
rect 57 297 60 300 
rect 57 300 60 303 
rect 57 303 60 306 
rect 57 306 60 309 
rect 57 309 60 312 
rect 57 312 60 315 
rect 57 315 60 318 
rect 57 318 60 321 
rect 57 321 60 324 
rect 57 324 60 327 
rect 57 327 60 330 
rect 57 330 60 333 
rect 57 333 60 336 
rect 57 336 60 339 
rect 57 339 60 342 
rect 57 342 60 345 
rect 57 345 60 348 
rect 57 348 60 351 
rect 57 351 60 354 
rect 57 354 60 357 
rect 57 357 60 360 
rect 57 360 60 363 
rect 57 363 60 366 
rect 57 366 60 369 
rect 57 369 60 372 
rect 57 372 60 375 
rect 57 375 60 378 
rect 57 378 60 381 
rect 57 381 60 384 
rect 57 384 60 387 
rect 57 387 60 390 
rect 57 390 60 393 
rect 57 393 60 396 
rect 57 396 60 399 
rect 57 399 60 402 
rect 57 402 60 405 
rect 57 405 60 408 
rect 57 408 60 411 
rect 57 411 60 414 
rect 57 414 60 417 
rect 57 417 60 420 
rect 57 420 60 423 
rect 57 423 60 426 
rect 57 426 60 429 
rect 57 429 60 432 
rect 57 432 60 435 
rect 57 435 60 438 
rect 57 438 60 441 
rect 57 441 60 444 
rect 57 444 60 447 
rect 57 447 60 450 
rect 57 450 60 453 
rect 57 453 60 456 
rect 57 456 60 459 
rect 57 459 60 462 
rect 57 462 60 465 
rect 57 465 60 468 
rect 57 468 60 471 
rect 57 471 60 474 
rect 57 474 60 477 
rect 57 477 60 480 
rect 57 480 60 483 
rect 57 483 60 486 
rect 57 486 60 489 
rect 57 489 60 492 
rect 57 492 60 495 
rect 57 495 60 498 
rect 57 498 60 501 
rect 57 501 60 504 
rect 57 504 60 507 
rect 57 507 60 510 
rect 60 0 63 3 
rect 60 3 63 6 
rect 60 6 63 9 
rect 60 9 63 12 
rect 60 12 63 15 
rect 60 15 63 18 
rect 60 18 63 21 
rect 60 21 63 24 
rect 60 24 63 27 
rect 60 27 63 30 
rect 60 30 63 33 
rect 60 33 63 36 
rect 60 36 63 39 
rect 60 39 63 42 
rect 60 42 63 45 
rect 60 45 63 48 
rect 60 48 63 51 
rect 60 51 63 54 
rect 60 54 63 57 
rect 60 57 63 60 
rect 60 60 63 63 
rect 60 63 63 66 
rect 60 66 63 69 
rect 60 69 63 72 
rect 60 72 63 75 
rect 60 75 63 78 
rect 60 78 63 81 
rect 60 81 63 84 
rect 60 84 63 87 
rect 60 87 63 90 
rect 60 90 63 93 
rect 60 93 63 96 
rect 60 96 63 99 
rect 60 99 63 102 
rect 60 102 63 105 
rect 60 105 63 108 
rect 60 108 63 111 
rect 60 111 63 114 
rect 60 114 63 117 
rect 60 117 63 120 
rect 60 120 63 123 
rect 60 123 63 126 
rect 60 126 63 129 
rect 60 129 63 132 
rect 60 132 63 135 
rect 60 135 63 138 
rect 60 138 63 141 
rect 60 141 63 144 
rect 60 144 63 147 
rect 60 147 63 150 
rect 60 150 63 153 
rect 60 153 63 156 
rect 60 156 63 159 
rect 60 159 63 162 
rect 60 162 63 165 
rect 60 165 63 168 
rect 60 168 63 171 
rect 60 171 63 174 
rect 60 174 63 177 
rect 60 177 63 180 
rect 60 180 63 183 
rect 60 183 63 186 
rect 60 186 63 189 
rect 60 189 63 192 
rect 60 192 63 195 
rect 60 195 63 198 
rect 60 198 63 201 
rect 60 201 63 204 
rect 60 204 63 207 
rect 60 207 63 210 
rect 60 210 63 213 
rect 60 213 63 216 
rect 60 216 63 219 
rect 60 219 63 222 
rect 60 222 63 225 
rect 60 225 63 228 
rect 60 228 63 231 
rect 60 231 63 234 
rect 60 234 63 237 
rect 60 237 63 240 
rect 60 240 63 243 
rect 60 243 63 246 
rect 60 246 63 249 
rect 60 249 63 252 
rect 60 252 63 255 
rect 60 255 63 258 
rect 60 258 63 261 
rect 60 261 63 264 
rect 60 264 63 267 
rect 60 267 63 270 
rect 60 270 63 273 
rect 60 273 63 276 
rect 60 276 63 279 
rect 60 279 63 282 
rect 60 282 63 285 
rect 60 285 63 288 
rect 60 288 63 291 
rect 60 291 63 294 
rect 60 294 63 297 
rect 60 297 63 300 
rect 60 300 63 303 
rect 60 303 63 306 
rect 60 306 63 309 
rect 60 309 63 312 
rect 60 312 63 315 
rect 60 315 63 318 
rect 60 318 63 321 
rect 60 321 63 324 
rect 60 324 63 327 
rect 60 327 63 330 
rect 60 330 63 333 
rect 60 333 63 336 
rect 60 336 63 339 
rect 60 339 63 342 
rect 60 342 63 345 
rect 60 345 63 348 
rect 60 348 63 351 
rect 60 351 63 354 
rect 60 354 63 357 
rect 60 357 63 360 
rect 60 360 63 363 
rect 60 363 63 366 
rect 60 366 63 369 
rect 60 369 63 372 
rect 60 372 63 375 
rect 60 375 63 378 
rect 60 378 63 381 
rect 60 381 63 384 
rect 60 384 63 387 
rect 60 387 63 390 
rect 60 390 63 393 
rect 60 393 63 396 
rect 60 396 63 399 
rect 60 399 63 402 
rect 60 402 63 405 
rect 60 405 63 408 
rect 60 408 63 411 
rect 60 411 63 414 
rect 60 414 63 417 
rect 60 417 63 420 
rect 60 420 63 423 
rect 60 423 63 426 
rect 60 426 63 429 
rect 60 429 63 432 
rect 60 432 63 435 
rect 60 435 63 438 
rect 60 438 63 441 
rect 60 441 63 444 
rect 60 444 63 447 
rect 60 447 63 450 
rect 60 450 63 453 
rect 60 453 63 456 
rect 60 456 63 459 
rect 60 459 63 462 
rect 60 462 63 465 
rect 60 465 63 468 
rect 60 468 63 471 
rect 60 471 63 474 
rect 60 474 63 477 
rect 60 477 63 480 
rect 60 480 63 483 
rect 60 483 63 486 
rect 60 486 63 489 
rect 60 489 63 492 
rect 60 492 63 495 
rect 60 495 63 498 
rect 60 498 63 501 
rect 60 501 63 504 
rect 60 504 63 507 
rect 60 507 63 510 
rect 63 0 66 3 
rect 63 3 66 6 
rect 63 6 66 9 
rect 63 9 66 12 
rect 63 12 66 15 
rect 63 15 66 18 
rect 63 18 66 21 
rect 63 21 66 24 
rect 63 24 66 27 
rect 63 27 66 30 
rect 63 30 66 33 
rect 63 33 66 36 
rect 63 36 66 39 
rect 63 39 66 42 
rect 63 42 66 45 
rect 63 45 66 48 
rect 63 48 66 51 
rect 63 51 66 54 
rect 63 54 66 57 
rect 63 57 66 60 
rect 63 60 66 63 
rect 63 63 66 66 
rect 63 66 66 69 
rect 63 69 66 72 
rect 63 72 66 75 
rect 63 75 66 78 
rect 63 78 66 81 
rect 63 81 66 84 
rect 63 84 66 87 
rect 63 87 66 90 
rect 63 90 66 93 
rect 63 93 66 96 
rect 63 96 66 99 
rect 63 99 66 102 
rect 63 102 66 105 
rect 63 105 66 108 
rect 63 108 66 111 
rect 63 111 66 114 
rect 63 114 66 117 
rect 63 117 66 120 
rect 63 120 66 123 
rect 63 123 66 126 
rect 63 126 66 129 
rect 63 129 66 132 
rect 63 132 66 135 
rect 63 135 66 138 
rect 63 138 66 141 
rect 63 141 66 144 
rect 63 144 66 147 
rect 63 147 66 150 
rect 63 150 66 153 
rect 63 153 66 156 
rect 63 156 66 159 
rect 63 159 66 162 
rect 63 162 66 165 
rect 63 165 66 168 
rect 63 168 66 171 
rect 63 171 66 174 
rect 63 174 66 177 
rect 63 177 66 180 
rect 63 180 66 183 
rect 63 183 66 186 
rect 63 186 66 189 
rect 63 189 66 192 
rect 63 192 66 195 
rect 63 195 66 198 
rect 63 198 66 201 
rect 63 201 66 204 
rect 63 204 66 207 
rect 63 207 66 210 
rect 63 210 66 213 
rect 63 213 66 216 
rect 63 216 66 219 
rect 63 219 66 222 
rect 63 222 66 225 
rect 63 225 66 228 
rect 63 228 66 231 
rect 63 231 66 234 
rect 63 234 66 237 
rect 63 237 66 240 
rect 63 240 66 243 
rect 63 243 66 246 
rect 63 246 66 249 
rect 63 249 66 252 
rect 63 252 66 255 
rect 63 255 66 258 
rect 63 258 66 261 
rect 63 261 66 264 
rect 63 264 66 267 
rect 63 267 66 270 
rect 63 270 66 273 
rect 63 273 66 276 
rect 63 276 66 279 
rect 63 279 66 282 
rect 63 282 66 285 
rect 63 285 66 288 
rect 63 288 66 291 
rect 63 291 66 294 
rect 63 294 66 297 
rect 63 297 66 300 
rect 63 300 66 303 
rect 63 303 66 306 
rect 63 306 66 309 
rect 63 309 66 312 
rect 63 312 66 315 
rect 63 315 66 318 
rect 63 318 66 321 
rect 63 321 66 324 
rect 63 324 66 327 
rect 63 327 66 330 
rect 63 330 66 333 
rect 63 333 66 336 
rect 63 336 66 339 
rect 63 339 66 342 
rect 63 342 66 345 
rect 63 345 66 348 
rect 63 348 66 351 
rect 63 351 66 354 
rect 63 354 66 357 
rect 63 357 66 360 
rect 63 360 66 363 
rect 63 363 66 366 
rect 63 366 66 369 
rect 63 369 66 372 
rect 63 372 66 375 
rect 63 375 66 378 
rect 63 378 66 381 
rect 63 381 66 384 
rect 63 384 66 387 
rect 63 387 66 390 
rect 63 390 66 393 
rect 63 393 66 396 
rect 63 396 66 399 
rect 63 399 66 402 
rect 63 402 66 405 
rect 63 405 66 408 
rect 63 408 66 411 
rect 63 411 66 414 
rect 63 414 66 417 
rect 63 417 66 420 
rect 63 420 66 423 
rect 63 423 66 426 
rect 63 426 66 429 
rect 63 429 66 432 
rect 63 432 66 435 
rect 63 435 66 438 
rect 63 438 66 441 
rect 63 441 66 444 
rect 63 444 66 447 
rect 63 447 66 450 
rect 63 450 66 453 
rect 63 453 66 456 
rect 63 456 66 459 
rect 63 459 66 462 
rect 63 462 66 465 
rect 63 465 66 468 
rect 63 468 66 471 
rect 63 471 66 474 
rect 63 474 66 477 
rect 63 477 66 480 
rect 63 480 66 483 
rect 63 483 66 486 
rect 63 486 66 489 
rect 63 489 66 492 
rect 63 492 66 495 
rect 63 495 66 498 
rect 63 498 66 501 
rect 63 501 66 504 
rect 63 504 66 507 
rect 63 507 66 510 
rect 66 0 69 3 
rect 66 3 69 6 
rect 66 6 69 9 
rect 66 9 69 12 
rect 66 12 69 15 
rect 66 15 69 18 
rect 66 18 69 21 
rect 66 21 69 24 
rect 66 24 69 27 
rect 66 27 69 30 
rect 66 30 69 33 
rect 66 33 69 36 
rect 66 36 69 39 
rect 66 39 69 42 
rect 66 42 69 45 
rect 66 45 69 48 
rect 66 48 69 51 
rect 66 51 69 54 
rect 66 54 69 57 
rect 66 57 69 60 
rect 66 60 69 63 
rect 66 63 69 66 
rect 66 66 69 69 
rect 66 69 69 72 
rect 66 72 69 75 
rect 66 75 69 78 
rect 66 78 69 81 
rect 66 81 69 84 
rect 66 84 69 87 
rect 66 87 69 90 
rect 66 90 69 93 
rect 66 93 69 96 
rect 66 96 69 99 
rect 66 99 69 102 
rect 66 102 69 105 
rect 66 105 69 108 
rect 66 108 69 111 
rect 66 111 69 114 
rect 66 114 69 117 
rect 66 117 69 120 
rect 66 120 69 123 
rect 66 123 69 126 
rect 66 126 69 129 
rect 66 129 69 132 
rect 66 132 69 135 
rect 66 135 69 138 
rect 66 138 69 141 
rect 66 141 69 144 
rect 66 144 69 147 
rect 66 147 69 150 
rect 66 150 69 153 
rect 66 153 69 156 
rect 66 156 69 159 
rect 66 159 69 162 
rect 66 162 69 165 
rect 66 165 69 168 
rect 66 168 69 171 
rect 66 171 69 174 
rect 66 174 69 177 
rect 66 177 69 180 
rect 66 180 69 183 
rect 66 183 69 186 
rect 66 186 69 189 
rect 66 189 69 192 
rect 66 192 69 195 
rect 66 195 69 198 
rect 66 198 69 201 
rect 66 201 69 204 
rect 66 204 69 207 
rect 66 207 69 210 
rect 66 210 69 213 
rect 66 213 69 216 
rect 66 216 69 219 
rect 66 219 69 222 
rect 66 222 69 225 
rect 66 225 69 228 
rect 66 228 69 231 
rect 66 231 69 234 
rect 66 234 69 237 
rect 66 237 69 240 
rect 66 240 69 243 
rect 66 243 69 246 
rect 66 246 69 249 
rect 66 249 69 252 
rect 66 252 69 255 
rect 66 255 69 258 
rect 66 258 69 261 
rect 66 261 69 264 
rect 66 264 69 267 
rect 66 267 69 270 
rect 66 270 69 273 
rect 66 273 69 276 
rect 66 276 69 279 
rect 66 279 69 282 
rect 66 282 69 285 
rect 66 285 69 288 
rect 66 288 69 291 
rect 66 291 69 294 
rect 66 294 69 297 
rect 66 297 69 300 
rect 66 300 69 303 
rect 66 303 69 306 
rect 66 306 69 309 
rect 66 309 69 312 
rect 66 312 69 315 
rect 66 315 69 318 
rect 66 318 69 321 
rect 66 321 69 324 
rect 66 324 69 327 
rect 66 327 69 330 
rect 66 330 69 333 
rect 66 333 69 336 
rect 66 336 69 339 
rect 66 339 69 342 
rect 66 342 69 345 
rect 66 345 69 348 
rect 66 348 69 351 
rect 66 351 69 354 
rect 66 354 69 357 
rect 66 357 69 360 
rect 66 360 69 363 
rect 66 363 69 366 
rect 66 366 69 369 
rect 66 369 69 372 
rect 66 372 69 375 
rect 66 375 69 378 
rect 66 378 69 381 
rect 66 381 69 384 
rect 66 384 69 387 
rect 66 387 69 390 
rect 66 390 69 393 
rect 66 393 69 396 
rect 66 396 69 399 
rect 66 399 69 402 
rect 66 402 69 405 
rect 66 405 69 408 
rect 66 408 69 411 
rect 66 411 69 414 
rect 66 414 69 417 
rect 66 417 69 420 
rect 66 420 69 423 
rect 66 423 69 426 
rect 66 426 69 429 
rect 66 429 69 432 
rect 66 432 69 435 
rect 66 435 69 438 
rect 66 438 69 441 
rect 66 441 69 444 
rect 66 444 69 447 
rect 66 447 69 450 
rect 66 450 69 453 
rect 66 453 69 456 
rect 66 456 69 459 
rect 66 459 69 462 
rect 66 462 69 465 
rect 66 465 69 468 
rect 66 468 69 471 
rect 66 471 69 474 
rect 66 474 69 477 
rect 66 477 69 480 
rect 66 480 69 483 
rect 66 483 69 486 
rect 66 486 69 489 
rect 66 489 69 492 
rect 66 492 69 495 
rect 66 495 69 498 
rect 66 498 69 501 
rect 66 501 69 504 
rect 66 504 69 507 
rect 66 507 69 510 
rect 69 0 72 3 
rect 69 3 72 6 
rect 69 6 72 9 
rect 69 9 72 12 
rect 69 12 72 15 
rect 69 15 72 18 
rect 69 18 72 21 
rect 69 21 72 24 
rect 69 24 72 27 
rect 69 27 72 30 
rect 69 30 72 33 
rect 69 33 72 36 
rect 69 36 72 39 
rect 69 39 72 42 
rect 69 42 72 45 
rect 69 45 72 48 
rect 69 48 72 51 
rect 69 51 72 54 
rect 69 54 72 57 
rect 69 57 72 60 
rect 69 60 72 63 
rect 69 63 72 66 
rect 69 66 72 69 
rect 69 69 72 72 
rect 69 72 72 75 
rect 69 75 72 78 
rect 69 78 72 81 
rect 69 81 72 84 
rect 69 84 72 87 
rect 69 87 72 90 
rect 69 90 72 93 
rect 69 93 72 96 
rect 69 96 72 99 
rect 69 99 72 102 
rect 69 102 72 105 
rect 69 105 72 108 
rect 69 108 72 111 
rect 69 111 72 114 
rect 69 114 72 117 
rect 69 117 72 120 
rect 69 120 72 123 
rect 69 123 72 126 
rect 69 126 72 129 
rect 69 129 72 132 
rect 69 132 72 135 
rect 69 135 72 138 
rect 69 138 72 141 
rect 69 141 72 144 
rect 69 144 72 147 
rect 69 147 72 150 
rect 69 150 72 153 
rect 69 153 72 156 
rect 69 156 72 159 
rect 69 159 72 162 
rect 69 162 72 165 
rect 69 165 72 168 
rect 69 168 72 171 
rect 69 171 72 174 
rect 69 174 72 177 
rect 69 177 72 180 
rect 69 180 72 183 
rect 69 183 72 186 
rect 69 186 72 189 
rect 69 189 72 192 
rect 69 192 72 195 
rect 69 195 72 198 
rect 69 198 72 201 
rect 69 201 72 204 
rect 69 204 72 207 
rect 69 207 72 210 
rect 69 210 72 213 
rect 69 213 72 216 
rect 69 216 72 219 
rect 69 219 72 222 
rect 69 222 72 225 
rect 69 225 72 228 
rect 69 228 72 231 
rect 69 231 72 234 
rect 69 234 72 237 
rect 69 237 72 240 
rect 69 240 72 243 
rect 69 243 72 246 
rect 69 246 72 249 
rect 69 249 72 252 
rect 69 252 72 255 
rect 69 255 72 258 
rect 69 258 72 261 
rect 69 261 72 264 
rect 69 264 72 267 
rect 69 267 72 270 
rect 69 270 72 273 
rect 69 273 72 276 
rect 69 276 72 279 
rect 69 279 72 282 
rect 69 282 72 285 
rect 69 285 72 288 
rect 69 288 72 291 
rect 69 291 72 294 
rect 69 294 72 297 
rect 69 297 72 300 
rect 69 300 72 303 
rect 69 303 72 306 
rect 69 306 72 309 
rect 69 309 72 312 
rect 69 312 72 315 
rect 69 315 72 318 
rect 69 318 72 321 
rect 69 321 72 324 
rect 69 324 72 327 
rect 69 327 72 330 
rect 69 330 72 333 
rect 69 333 72 336 
rect 69 336 72 339 
rect 69 339 72 342 
rect 69 342 72 345 
rect 69 345 72 348 
rect 69 348 72 351 
rect 69 351 72 354 
rect 69 354 72 357 
rect 69 357 72 360 
rect 69 360 72 363 
rect 69 363 72 366 
rect 69 366 72 369 
rect 69 369 72 372 
rect 69 372 72 375 
rect 69 375 72 378 
rect 69 378 72 381 
rect 69 381 72 384 
rect 69 384 72 387 
rect 69 387 72 390 
rect 69 390 72 393 
rect 69 393 72 396 
rect 69 396 72 399 
rect 69 399 72 402 
rect 69 402 72 405 
rect 69 405 72 408 
rect 69 408 72 411 
rect 69 411 72 414 
rect 69 414 72 417 
rect 69 417 72 420 
rect 69 420 72 423 
rect 69 423 72 426 
rect 69 426 72 429 
rect 69 429 72 432 
rect 69 432 72 435 
rect 69 435 72 438 
rect 69 438 72 441 
rect 69 441 72 444 
rect 69 444 72 447 
rect 69 447 72 450 
rect 69 450 72 453 
rect 69 453 72 456 
rect 69 456 72 459 
rect 69 459 72 462 
rect 69 462 72 465 
rect 69 465 72 468 
rect 69 468 72 471 
rect 69 471 72 474 
rect 69 474 72 477 
rect 69 477 72 480 
rect 69 480 72 483 
rect 69 483 72 486 
rect 69 486 72 489 
rect 69 489 72 492 
rect 69 492 72 495 
rect 69 495 72 498 
rect 69 498 72 501 
rect 69 501 72 504 
rect 69 504 72 507 
rect 69 507 72 510 
rect 72 0 75 3 
rect 72 3 75 6 
rect 72 6 75 9 
rect 72 9 75 12 
rect 72 12 75 15 
rect 72 15 75 18 
rect 72 18 75 21 
rect 72 21 75 24 
rect 72 24 75 27 
rect 72 27 75 30 
rect 72 30 75 33 
rect 72 33 75 36 
rect 72 36 75 39 
rect 72 39 75 42 
rect 72 42 75 45 
rect 72 45 75 48 
rect 72 48 75 51 
rect 72 51 75 54 
rect 72 54 75 57 
rect 72 57 75 60 
rect 72 60 75 63 
rect 72 63 75 66 
rect 72 66 75 69 
rect 72 69 75 72 
rect 72 72 75 75 
rect 72 75 75 78 
rect 72 78 75 81 
rect 72 81 75 84 
rect 72 84 75 87 
rect 72 87 75 90 
rect 72 90 75 93 
rect 72 93 75 96 
rect 72 96 75 99 
rect 72 99 75 102 
rect 72 102 75 105 
rect 72 105 75 108 
rect 72 108 75 111 
rect 72 111 75 114 
rect 72 114 75 117 
rect 72 117 75 120 
rect 72 120 75 123 
rect 72 123 75 126 
rect 72 126 75 129 
rect 72 129 75 132 
rect 72 132 75 135 
rect 72 135 75 138 
rect 72 138 75 141 
rect 72 141 75 144 
rect 72 144 75 147 
rect 72 147 75 150 
rect 72 150 75 153 
rect 72 153 75 156 
rect 72 156 75 159 
rect 72 159 75 162 
rect 72 162 75 165 
rect 72 165 75 168 
rect 72 168 75 171 
rect 72 171 75 174 
rect 72 174 75 177 
rect 72 177 75 180 
rect 72 180 75 183 
rect 72 183 75 186 
rect 72 186 75 189 
rect 72 189 75 192 
rect 72 192 75 195 
rect 72 195 75 198 
rect 72 198 75 201 
rect 72 201 75 204 
rect 72 204 75 207 
rect 72 207 75 210 
rect 72 210 75 213 
rect 72 213 75 216 
rect 72 216 75 219 
rect 72 219 75 222 
rect 72 222 75 225 
rect 72 225 75 228 
rect 72 228 75 231 
rect 72 231 75 234 
rect 72 234 75 237 
rect 72 237 75 240 
rect 72 240 75 243 
rect 72 243 75 246 
rect 72 246 75 249 
rect 72 249 75 252 
rect 72 252 75 255 
rect 72 255 75 258 
rect 72 258 75 261 
rect 72 261 75 264 
rect 72 264 75 267 
rect 72 267 75 270 
rect 72 270 75 273 
rect 72 273 75 276 
rect 72 276 75 279 
rect 72 279 75 282 
rect 72 282 75 285 
rect 72 285 75 288 
rect 72 288 75 291 
rect 72 291 75 294 
rect 72 294 75 297 
rect 72 297 75 300 
rect 72 300 75 303 
rect 72 303 75 306 
rect 72 306 75 309 
rect 72 309 75 312 
rect 72 312 75 315 
rect 72 315 75 318 
rect 72 318 75 321 
rect 72 321 75 324 
rect 72 324 75 327 
rect 72 327 75 330 
rect 72 330 75 333 
rect 72 333 75 336 
rect 72 336 75 339 
rect 72 339 75 342 
rect 72 342 75 345 
rect 72 345 75 348 
rect 72 348 75 351 
rect 72 351 75 354 
rect 72 354 75 357 
rect 72 357 75 360 
rect 72 360 75 363 
rect 72 363 75 366 
rect 72 366 75 369 
rect 72 369 75 372 
rect 72 372 75 375 
rect 72 375 75 378 
rect 72 378 75 381 
rect 72 381 75 384 
rect 72 384 75 387 
rect 72 387 75 390 
rect 72 390 75 393 
rect 72 393 75 396 
rect 72 396 75 399 
rect 72 399 75 402 
rect 72 402 75 405 
rect 72 405 75 408 
rect 72 408 75 411 
rect 72 411 75 414 
rect 72 414 75 417 
rect 72 417 75 420 
rect 72 420 75 423 
rect 72 423 75 426 
rect 72 426 75 429 
rect 72 429 75 432 
rect 72 432 75 435 
rect 72 435 75 438 
rect 72 438 75 441 
rect 72 441 75 444 
rect 72 444 75 447 
rect 72 447 75 450 
rect 72 450 75 453 
rect 72 453 75 456 
rect 72 456 75 459 
rect 72 459 75 462 
rect 72 462 75 465 
rect 72 465 75 468 
rect 72 468 75 471 
rect 72 471 75 474 
rect 72 474 75 477 
rect 72 477 75 480 
rect 72 480 75 483 
rect 72 483 75 486 
rect 72 486 75 489 
rect 72 489 75 492 
rect 72 492 75 495 
rect 72 495 75 498 
rect 72 498 75 501 
rect 72 501 75 504 
rect 72 504 75 507 
rect 72 507 75 510 
rect 75 0 78 3 
rect 75 3 78 6 
rect 75 6 78 9 
rect 75 9 78 12 
rect 75 12 78 15 
rect 75 15 78 18 
rect 75 18 78 21 
rect 75 21 78 24 
rect 75 24 78 27 
rect 75 27 78 30 
rect 75 30 78 33 
rect 75 33 78 36 
rect 75 36 78 39 
rect 75 39 78 42 
rect 75 42 78 45 
rect 75 45 78 48 
rect 75 48 78 51 
rect 75 51 78 54 
rect 75 54 78 57 
rect 75 57 78 60 
rect 75 60 78 63 
rect 75 63 78 66 
rect 75 66 78 69 
rect 75 69 78 72 
rect 75 72 78 75 
rect 75 75 78 78 
rect 75 78 78 81 
rect 75 81 78 84 
rect 75 84 78 87 
rect 75 87 78 90 
rect 75 90 78 93 
rect 75 93 78 96 
rect 75 96 78 99 
rect 75 99 78 102 
rect 75 102 78 105 
rect 75 105 78 108 
rect 75 108 78 111 
rect 75 111 78 114 
rect 75 114 78 117 
rect 75 117 78 120 
rect 75 120 78 123 
rect 75 123 78 126 
rect 75 126 78 129 
rect 75 129 78 132 
rect 75 132 78 135 
rect 75 135 78 138 
rect 75 138 78 141 
rect 75 141 78 144 
rect 75 144 78 147 
rect 75 147 78 150 
rect 75 150 78 153 
rect 75 153 78 156 
rect 75 156 78 159 
rect 75 159 78 162 
rect 75 162 78 165 
rect 75 165 78 168 
rect 75 168 78 171 
rect 75 171 78 174 
rect 75 174 78 177 
rect 75 177 78 180 
rect 75 180 78 183 
rect 75 183 78 186 
rect 75 186 78 189 
rect 75 189 78 192 
rect 75 192 78 195 
rect 75 195 78 198 
rect 75 198 78 201 
rect 75 201 78 204 
rect 75 204 78 207 
rect 75 207 78 210 
rect 75 210 78 213 
rect 75 213 78 216 
rect 75 216 78 219 
rect 75 219 78 222 
rect 75 222 78 225 
rect 75 225 78 228 
rect 75 228 78 231 
rect 75 231 78 234 
rect 75 234 78 237 
rect 75 237 78 240 
rect 75 240 78 243 
rect 75 243 78 246 
rect 75 246 78 249 
rect 75 249 78 252 
rect 75 252 78 255 
rect 75 255 78 258 
rect 75 258 78 261 
rect 75 261 78 264 
rect 75 264 78 267 
rect 75 267 78 270 
rect 75 270 78 273 
rect 75 273 78 276 
rect 75 276 78 279 
rect 75 279 78 282 
rect 75 282 78 285 
rect 75 285 78 288 
rect 75 288 78 291 
rect 75 291 78 294 
rect 75 294 78 297 
rect 75 297 78 300 
rect 75 300 78 303 
rect 75 303 78 306 
rect 75 306 78 309 
rect 75 309 78 312 
rect 75 312 78 315 
rect 75 315 78 318 
rect 75 318 78 321 
rect 75 321 78 324 
rect 75 324 78 327 
rect 75 327 78 330 
rect 75 330 78 333 
rect 75 333 78 336 
rect 75 336 78 339 
rect 75 339 78 342 
rect 75 342 78 345 
rect 75 345 78 348 
rect 75 348 78 351 
rect 75 351 78 354 
rect 75 354 78 357 
rect 75 357 78 360 
rect 75 360 78 363 
rect 75 363 78 366 
rect 75 366 78 369 
rect 75 369 78 372 
rect 75 372 78 375 
rect 75 375 78 378 
rect 75 378 78 381 
rect 75 381 78 384 
rect 75 384 78 387 
rect 75 387 78 390 
rect 75 390 78 393 
rect 75 393 78 396 
rect 75 396 78 399 
rect 75 399 78 402 
rect 75 402 78 405 
rect 75 405 78 408 
rect 75 408 78 411 
rect 75 411 78 414 
rect 75 414 78 417 
rect 75 417 78 420 
rect 75 420 78 423 
rect 75 423 78 426 
rect 75 426 78 429 
rect 75 429 78 432 
rect 75 432 78 435 
rect 75 435 78 438 
rect 75 438 78 441 
rect 75 441 78 444 
rect 75 444 78 447 
rect 75 447 78 450 
rect 75 450 78 453 
rect 75 453 78 456 
rect 75 456 78 459 
rect 75 459 78 462 
rect 75 462 78 465 
rect 75 465 78 468 
rect 75 468 78 471 
rect 75 471 78 474 
rect 75 474 78 477 
rect 75 477 78 480 
rect 75 480 78 483 
rect 75 483 78 486 
rect 75 486 78 489 
rect 75 489 78 492 
rect 75 492 78 495 
rect 75 495 78 498 
rect 75 498 78 501 
rect 75 501 78 504 
rect 75 504 78 507 
rect 75 507 78 510 
rect 78 0 81 3 
rect 78 3 81 6 
rect 78 6 81 9 
rect 78 9 81 12 
rect 78 12 81 15 
rect 78 15 81 18 
rect 78 18 81 21 
rect 78 21 81 24 
rect 78 24 81 27 
rect 78 27 81 30 
rect 78 30 81 33 
rect 78 33 81 36 
rect 78 36 81 39 
rect 78 39 81 42 
rect 78 42 81 45 
rect 78 45 81 48 
rect 78 48 81 51 
rect 78 51 81 54 
rect 78 54 81 57 
rect 78 57 81 60 
rect 78 60 81 63 
rect 78 63 81 66 
rect 78 66 81 69 
rect 78 69 81 72 
rect 78 72 81 75 
rect 78 75 81 78 
rect 78 78 81 81 
rect 78 81 81 84 
rect 78 84 81 87 
rect 78 87 81 90 
rect 78 90 81 93 
rect 78 93 81 96 
rect 78 96 81 99 
rect 78 99 81 102 
rect 78 102 81 105 
rect 78 105 81 108 
rect 78 108 81 111 
rect 78 111 81 114 
rect 78 114 81 117 
rect 78 117 81 120 
rect 78 120 81 123 
rect 78 123 81 126 
rect 78 126 81 129 
rect 78 129 81 132 
rect 78 132 81 135 
rect 78 135 81 138 
rect 78 141 81 144 
rect 78 144 81 147 
rect 78 147 81 150 
rect 78 150 81 153 
rect 78 153 81 156 
rect 78 156 81 159 
rect 78 159 81 162 
rect 78 162 81 165 
rect 78 165 81 168 
rect 78 168 81 171 
rect 78 171 81 174 
rect 78 174 81 177 
rect 78 177 81 180 
rect 78 180 81 183 
rect 78 183 81 186 
rect 78 186 81 189 
rect 78 189 81 192 
rect 78 192 81 195 
rect 78 195 81 198 
rect 78 198 81 201 
rect 78 201 81 204 
rect 78 204 81 207 
rect 78 207 81 210 
rect 78 210 81 213 
rect 78 213 81 216 
rect 78 216 81 219 
rect 78 219 81 222 
rect 78 222 81 225 
rect 78 225 81 228 
rect 78 228 81 231 
rect 78 231 81 234 
rect 78 234 81 237 
rect 78 237 81 240 
rect 78 240 81 243 
rect 78 243 81 246 
rect 78 246 81 249 
rect 78 249 81 252 
rect 78 252 81 255 
rect 78 255 81 258 
rect 78 258 81 261 
rect 78 261 81 264 
rect 78 264 81 267 
rect 78 267 81 270 
rect 78 270 81 273 
rect 78 273 81 276 
rect 78 276 81 279 
rect 78 279 81 282 
rect 78 282 81 285 
rect 78 285 81 288 
rect 78 288 81 291 
rect 78 291 81 294 
rect 78 294 81 297 
rect 78 297 81 300 
rect 78 300 81 303 
rect 78 303 81 306 
rect 78 306 81 309 
rect 78 309 81 312 
rect 78 312 81 315 
rect 78 315 81 318 
rect 78 318 81 321 
rect 78 321 81 324 
rect 78 324 81 327 
rect 78 327 81 330 
rect 78 330 81 333 
rect 78 333 81 336 
rect 78 336 81 339 
rect 78 339 81 342 
rect 78 342 81 345 
rect 78 345 81 348 
rect 78 348 81 351 
rect 78 351 81 354 
rect 78 354 81 357 
rect 78 357 81 360 
rect 78 360 81 363 
rect 78 363 81 366 
rect 78 366 81 369 
rect 78 369 81 372 
rect 78 372 81 375 
rect 78 375 81 378 
rect 78 378 81 381 
rect 78 381 81 384 
rect 78 384 81 387 
rect 78 387 81 390 
rect 78 390 81 393 
rect 78 393 81 396 
rect 78 396 81 399 
rect 78 399 81 402 
rect 78 402 81 405 
rect 78 405 81 408 
rect 78 408 81 411 
rect 78 411 81 414 
rect 78 414 81 417 
rect 78 420 81 423 
rect 78 423 81 426 
rect 78 426 81 429 
rect 78 429 81 432 
rect 78 432 81 435 
rect 78 435 81 438 
rect 78 438 81 441 
rect 78 441 81 444 
rect 78 444 81 447 
rect 78 447 81 450 
rect 78 450 81 453 
rect 78 453 81 456 
rect 78 456 81 459 
rect 78 459 81 462 
rect 78 462 81 465 
rect 78 468 81 471 
rect 78 471 81 474 
rect 78 477 81 480 
rect 78 480 81 483 
rect 78 483 81 486 
rect 78 486 81 489 
rect 78 489 81 492 
rect 78 492 81 495 
rect 78 495 81 498 
rect 78 498 81 501 
rect 78 501 81 504 
rect 78 504 81 507 
rect 78 507 81 510 
rect 81 0 84 3 
rect 81 3 84 6 
rect 81 6 84 9 
rect 81 9 84 12 
rect 81 12 84 15 
rect 81 15 84 18 
rect 81 18 84 21 
rect 81 21 84 24 
rect 81 24 84 27 
rect 81 27 84 30 
rect 81 30 84 33 
rect 81 33 84 36 
rect 81 36 84 39 
rect 81 39 84 42 
rect 81 42 84 45 
rect 81 45 84 48 
rect 81 48 84 51 
rect 81 51 84 54 
rect 81 54 84 57 
rect 81 57 84 60 
rect 81 60 84 63 
rect 81 63 84 66 
rect 81 66 84 69 
rect 81 69 84 72 
rect 81 72 84 75 
rect 81 75 84 78 
rect 81 78 84 81 
rect 81 81 84 84 
rect 81 84 84 87 
rect 81 87 84 90 
rect 81 90 84 93 
rect 81 93 84 96 
rect 81 96 84 99 
rect 81 99 84 102 
rect 81 102 84 105 
rect 81 105 84 108 
rect 81 108 84 111 
rect 81 111 84 114 
rect 81 114 84 117 
rect 81 117 84 120 
rect 81 120 84 123 
rect 81 123 84 126 
rect 81 126 84 129 
rect 81 129 84 132 
rect 81 132 84 135 
rect 81 135 84 138 
rect 81 138 84 141 
rect 81 141 84 144 
rect 81 144 84 147 
rect 81 147 84 150 
rect 81 150 84 153 
rect 81 153 84 156 
rect 81 156 84 159 
rect 81 159 84 162 
rect 81 162 84 165 
rect 81 165 84 168 
rect 81 168 84 171 
rect 81 171 84 174 
rect 81 174 84 177 
rect 81 177 84 180 
rect 81 180 84 183 
rect 81 183 84 186 
rect 81 186 84 189 
rect 81 189 84 192 
rect 81 192 84 195 
rect 81 195 84 198 
rect 81 198 84 201 
rect 81 201 84 204 
rect 81 204 84 207 
rect 81 207 84 210 
rect 81 210 84 213 
rect 81 213 84 216 
rect 81 216 84 219 
rect 81 219 84 222 
rect 81 222 84 225 
rect 81 225 84 228 
rect 81 228 84 231 
rect 81 231 84 234 
rect 81 234 84 237 
rect 81 237 84 240 
rect 81 240 84 243 
rect 81 243 84 246 
rect 81 246 84 249 
rect 81 249 84 252 
rect 81 252 84 255 
rect 81 255 84 258 
rect 81 258 84 261 
rect 81 261 84 264 
rect 81 264 84 267 
rect 81 267 84 270 
rect 81 270 84 273 
rect 81 273 84 276 
rect 81 276 84 279 
rect 81 279 84 282 
rect 81 282 84 285 
rect 81 285 84 288 
rect 81 288 84 291 
rect 81 291 84 294 
rect 81 294 84 297 
rect 81 297 84 300 
rect 81 300 84 303 
rect 81 303 84 306 
rect 81 306 84 309 
rect 81 309 84 312 
rect 81 312 84 315 
rect 81 315 84 318 
rect 81 318 84 321 
rect 81 321 84 324 
rect 81 324 84 327 
rect 81 327 84 330 
rect 81 330 84 333 
rect 81 333 84 336 
rect 81 336 84 339 
rect 81 339 84 342 
rect 81 342 84 345 
rect 81 345 84 348 
rect 81 348 84 351 
rect 81 351 84 354 
rect 81 354 84 357 
rect 81 357 84 360 
rect 81 360 84 363 
rect 81 363 84 366 
rect 81 366 84 369 
rect 81 369 84 372 
rect 81 372 84 375 
rect 81 375 84 378 
rect 81 378 84 381 
rect 81 381 84 384 
rect 81 384 84 387 
rect 81 387 84 390 
rect 81 390 84 393 
rect 81 393 84 396 
rect 81 396 84 399 
rect 81 399 84 402 
rect 81 402 84 405 
rect 81 405 84 408 
rect 81 408 84 411 
rect 81 411 84 414 
rect 81 414 84 417 
rect 81 417 84 420 
rect 81 420 84 423 
rect 81 423 84 426 
rect 81 426 84 429 
rect 81 429 84 432 
rect 81 432 84 435 
rect 81 435 84 438 
rect 81 438 84 441 
rect 81 441 84 444 
rect 81 444 84 447 
rect 81 447 84 450 
rect 81 450 84 453 
rect 81 453 84 456 
rect 81 456 84 459 
rect 81 459 84 462 
rect 81 462 84 465 
rect 81 465 84 468 
rect 81 468 84 471 
rect 81 471 84 474 
rect 81 474 84 477 
rect 81 477 84 480 
rect 81 480 84 483 
rect 81 483 84 486 
rect 81 486 84 489 
rect 81 489 84 492 
rect 81 492 84 495 
rect 81 495 84 498 
rect 81 498 84 501 
rect 81 501 84 504 
rect 81 504 84 507 
rect 81 507 84 510 
rect 84 0 87 3 
rect 84 3 87 6 
rect 84 6 87 9 
rect 84 9 87 12 
rect 84 12 87 15 
rect 84 15 87 18 
rect 84 18 87 21 
rect 84 21 87 24 
rect 84 24 87 27 
rect 84 27 87 30 
rect 84 30 87 33 
rect 84 33 87 36 
rect 84 36 87 39 
rect 84 39 87 42 
rect 84 42 87 45 
rect 84 45 87 48 
rect 84 48 87 51 
rect 84 51 87 54 
rect 84 54 87 57 
rect 84 57 87 60 
rect 84 60 87 63 
rect 84 63 87 66 
rect 84 66 87 69 
rect 84 69 87 72 
rect 84 72 87 75 
rect 84 75 87 78 
rect 84 78 87 81 
rect 84 81 87 84 
rect 84 84 87 87 
rect 84 87 87 90 
rect 84 90 87 93 
rect 84 93 87 96 
rect 84 96 87 99 
rect 84 99 87 102 
rect 84 102 87 105 
rect 84 105 87 108 
rect 84 108 87 111 
rect 84 111 87 114 
rect 84 114 87 117 
rect 84 117 87 120 
rect 84 120 87 123 
rect 84 123 87 126 
rect 84 126 87 129 
rect 84 129 87 132 
rect 84 132 87 135 
rect 84 135 87 138 
rect 84 138 87 141 
rect 84 141 87 144 
rect 84 144 87 147 
rect 84 147 87 150 
rect 84 150 87 153 
rect 84 153 87 156 
rect 84 156 87 159 
rect 84 159 87 162 
rect 84 162 87 165 
rect 84 165 87 168 
rect 84 168 87 171 
rect 84 171 87 174 
rect 84 174 87 177 
rect 84 177 87 180 
rect 84 180 87 183 
rect 84 183 87 186 
rect 84 186 87 189 
rect 84 189 87 192 
rect 84 192 87 195 
rect 84 195 87 198 
rect 84 198 87 201 
rect 84 201 87 204 
rect 84 204 87 207 
rect 84 207 87 210 
rect 84 210 87 213 
rect 84 213 87 216 
rect 84 216 87 219 
rect 84 219 87 222 
rect 84 222 87 225 
rect 84 225 87 228 
rect 84 228 87 231 
rect 84 231 87 234 
rect 84 234 87 237 
rect 84 237 87 240 
rect 84 240 87 243 
rect 84 243 87 246 
rect 84 246 87 249 
rect 84 249 87 252 
rect 84 252 87 255 
rect 84 255 87 258 
rect 84 258 87 261 
rect 84 261 87 264 
rect 84 264 87 267 
rect 84 267 87 270 
rect 84 270 87 273 
rect 84 273 87 276 
rect 84 276 87 279 
rect 84 279 87 282 
rect 84 282 87 285 
rect 84 285 87 288 
rect 84 288 87 291 
rect 84 291 87 294 
rect 84 294 87 297 
rect 84 297 87 300 
rect 84 300 87 303 
rect 84 303 87 306 
rect 84 306 87 309 
rect 84 309 87 312 
rect 84 312 87 315 
rect 84 315 87 318 
rect 84 318 87 321 
rect 84 321 87 324 
rect 84 324 87 327 
rect 84 327 87 330 
rect 84 330 87 333 
rect 84 333 87 336 
rect 84 336 87 339 
rect 84 339 87 342 
rect 84 342 87 345 
rect 84 345 87 348 
rect 84 348 87 351 
rect 84 351 87 354 
rect 84 354 87 357 
rect 84 357 87 360 
rect 84 360 87 363 
rect 84 363 87 366 
rect 84 366 87 369 
rect 84 369 87 372 
rect 84 372 87 375 
rect 84 375 87 378 
rect 84 378 87 381 
rect 84 381 87 384 
rect 84 384 87 387 
rect 84 387 87 390 
rect 84 390 87 393 
rect 84 393 87 396 
rect 84 396 87 399 
rect 84 399 87 402 
rect 84 402 87 405 
rect 84 405 87 408 
rect 84 408 87 411 
rect 84 411 87 414 
rect 84 414 87 417 
rect 84 417 87 420 
rect 84 420 87 423 
rect 84 423 87 426 
rect 84 426 87 429 
rect 84 429 87 432 
rect 84 432 87 435 
rect 84 435 87 438 
rect 84 438 87 441 
rect 84 441 87 444 
rect 84 444 87 447 
rect 84 447 87 450 
rect 84 450 87 453 
rect 84 453 87 456 
rect 84 456 87 459 
rect 84 459 87 462 
rect 84 462 87 465 
rect 84 465 87 468 
rect 84 468 87 471 
rect 84 471 87 474 
rect 84 474 87 477 
rect 84 477 87 480 
rect 84 480 87 483 
rect 84 483 87 486 
rect 84 486 87 489 
rect 84 489 87 492 
rect 84 492 87 495 
rect 84 495 87 498 
rect 84 498 87 501 
rect 84 501 87 504 
rect 84 504 87 507 
rect 84 507 87 510 
rect 87 0 90 3 
rect 87 3 90 6 
rect 87 6 90 9 
rect 87 9 90 12 
rect 87 12 90 15 
rect 87 15 90 18 
rect 87 18 90 21 
rect 87 21 90 24 
rect 87 24 90 27 
rect 87 27 90 30 
rect 87 30 90 33 
rect 87 33 90 36 
rect 87 36 90 39 
rect 87 39 90 42 
rect 87 42 90 45 
rect 87 45 90 48 
rect 87 48 90 51 
rect 87 51 90 54 
rect 87 54 90 57 
rect 87 57 90 60 
rect 87 60 90 63 
rect 87 63 90 66 
rect 87 66 90 69 
rect 87 69 90 72 
rect 87 72 90 75 
rect 87 75 90 78 
rect 87 78 90 81 
rect 87 81 90 84 
rect 87 84 90 87 
rect 87 87 90 90 
rect 87 90 90 93 
rect 87 93 90 96 
rect 87 96 90 99 
rect 87 99 90 102 
rect 87 102 90 105 
rect 87 105 90 108 
rect 87 108 90 111 
rect 87 111 90 114 
rect 87 114 90 117 
rect 87 117 90 120 
rect 87 120 90 123 
rect 87 123 90 126 
rect 87 126 90 129 
rect 87 129 90 132 
rect 87 132 90 135 
rect 87 135 90 138 
rect 87 138 90 141 
rect 87 141 90 144 
rect 87 144 90 147 
rect 87 147 90 150 
rect 87 150 90 153 
rect 87 153 90 156 
rect 87 156 90 159 
rect 87 159 90 162 
rect 87 162 90 165 
rect 87 165 90 168 
rect 87 168 90 171 
rect 87 171 90 174 
rect 87 174 90 177 
rect 87 177 90 180 
rect 87 180 90 183 
rect 87 183 90 186 
rect 87 186 90 189 
rect 87 189 90 192 
rect 87 192 90 195 
rect 87 195 90 198 
rect 87 198 90 201 
rect 87 201 90 204 
rect 87 204 90 207 
rect 87 207 90 210 
rect 87 210 90 213 
rect 87 213 90 216 
rect 87 216 90 219 
rect 87 219 90 222 
rect 87 222 90 225 
rect 87 225 90 228 
rect 87 228 90 231 
rect 87 231 90 234 
rect 87 234 90 237 
rect 87 237 90 240 
rect 87 240 90 243 
rect 87 243 90 246 
rect 87 246 90 249 
rect 87 249 90 252 
rect 87 252 90 255 
rect 87 255 90 258 
rect 87 258 90 261 
rect 87 261 90 264 
rect 87 264 90 267 
rect 87 267 90 270 
rect 87 270 90 273 
rect 87 273 90 276 
rect 87 276 90 279 
rect 87 279 90 282 
rect 87 282 90 285 
rect 87 285 90 288 
rect 87 288 90 291 
rect 87 291 90 294 
rect 87 294 90 297 
rect 87 297 90 300 
rect 87 300 90 303 
rect 87 303 90 306 
rect 87 306 90 309 
rect 87 309 90 312 
rect 87 312 90 315 
rect 87 315 90 318 
rect 87 318 90 321 
rect 87 321 90 324 
rect 87 324 90 327 
rect 87 327 90 330 
rect 87 330 90 333 
rect 87 333 90 336 
rect 87 336 90 339 
rect 87 339 90 342 
rect 87 342 90 345 
rect 87 345 90 348 
rect 87 348 90 351 
rect 87 351 90 354 
rect 87 354 90 357 
rect 87 357 90 360 
rect 87 360 90 363 
rect 87 363 90 366 
rect 87 366 90 369 
rect 87 369 90 372 
rect 87 372 90 375 
rect 87 375 90 378 
rect 87 378 90 381 
rect 87 381 90 384 
rect 87 384 90 387 
rect 87 387 90 390 
rect 87 390 90 393 
rect 87 393 90 396 
rect 87 396 90 399 
rect 87 399 90 402 
rect 87 402 90 405 
rect 87 405 90 408 
rect 87 408 90 411 
rect 87 411 90 414 
rect 87 414 90 417 
rect 87 417 90 420 
rect 87 420 90 423 
rect 87 423 90 426 
rect 87 426 90 429 
rect 87 429 90 432 
rect 87 432 90 435 
rect 87 435 90 438 
rect 87 438 90 441 
rect 87 441 90 444 
rect 87 444 90 447 
rect 87 447 90 450 
rect 87 450 90 453 
rect 87 453 90 456 
rect 87 456 90 459 
rect 87 459 90 462 
rect 87 462 90 465 
rect 87 465 90 468 
rect 87 468 90 471 
rect 87 471 90 474 
rect 87 474 90 477 
rect 87 477 90 480 
rect 87 480 90 483 
rect 87 483 90 486 
rect 87 486 90 489 
rect 87 489 90 492 
rect 87 492 90 495 
rect 87 495 90 498 
rect 87 498 90 501 
rect 87 501 90 504 
rect 87 504 90 507 
rect 87 507 90 510 
rect 90 0 93 3 
rect 90 3 93 6 
rect 90 6 93 9 
rect 90 9 93 12 
rect 90 12 93 15 
rect 90 15 93 18 
rect 90 18 93 21 
rect 90 21 93 24 
rect 90 24 93 27 
rect 90 27 93 30 
rect 90 30 93 33 
rect 90 33 93 36 
rect 90 36 93 39 
rect 90 39 93 42 
rect 90 42 93 45 
rect 90 45 93 48 
rect 90 48 93 51 
rect 90 51 93 54 
rect 90 54 93 57 
rect 90 57 93 60 
rect 90 60 93 63 
rect 90 63 93 66 
rect 90 66 93 69 
rect 90 69 93 72 
rect 90 72 93 75 
rect 90 75 93 78 
rect 90 78 93 81 
rect 90 81 93 84 
rect 90 84 93 87 
rect 90 87 93 90 
rect 90 90 93 93 
rect 90 93 93 96 
rect 90 96 93 99 
rect 90 99 93 102 
rect 90 102 93 105 
rect 90 105 93 108 
rect 90 108 93 111 
rect 90 111 93 114 
rect 90 114 93 117 
rect 90 117 93 120 
rect 90 120 93 123 
rect 90 123 93 126 
rect 90 126 93 129 
rect 90 129 93 132 
rect 90 132 93 135 
rect 90 135 93 138 
rect 90 138 93 141 
rect 90 141 93 144 
rect 90 144 93 147 
rect 90 147 93 150 
rect 90 150 93 153 
rect 90 153 93 156 
rect 90 156 93 159 
rect 90 159 93 162 
rect 90 162 93 165 
rect 90 165 93 168 
rect 90 168 93 171 
rect 90 171 93 174 
rect 90 174 93 177 
rect 90 177 93 180 
rect 90 180 93 183 
rect 90 183 93 186 
rect 90 186 93 189 
rect 90 189 93 192 
rect 90 192 93 195 
rect 90 195 93 198 
rect 90 198 93 201 
rect 90 201 93 204 
rect 90 204 93 207 
rect 90 207 93 210 
rect 90 210 93 213 
rect 90 213 93 216 
rect 90 216 93 219 
rect 90 219 93 222 
rect 90 222 93 225 
rect 90 225 93 228 
rect 90 228 93 231 
rect 90 231 93 234 
rect 90 234 93 237 
rect 90 237 93 240 
rect 90 240 93 243 
rect 90 243 93 246 
rect 90 246 93 249 
rect 90 249 93 252 
rect 90 252 93 255 
rect 90 255 93 258 
rect 90 258 93 261 
rect 90 261 93 264 
rect 90 264 93 267 
rect 90 267 93 270 
rect 90 270 93 273 
rect 90 273 93 276 
rect 90 276 93 279 
rect 90 279 93 282 
rect 90 282 93 285 
rect 90 285 93 288 
rect 90 288 93 291 
rect 90 291 93 294 
rect 90 294 93 297 
rect 90 297 93 300 
rect 90 300 93 303 
rect 90 303 93 306 
rect 90 306 93 309 
rect 90 309 93 312 
rect 90 312 93 315 
rect 90 315 93 318 
rect 90 318 93 321 
rect 90 321 93 324 
rect 90 324 93 327 
rect 90 327 93 330 
rect 90 330 93 333 
rect 90 333 93 336 
rect 90 336 93 339 
rect 90 339 93 342 
rect 90 342 93 345 
rect 90 345 93 348 
rect 90 348 93 351 
rect 90 351 93 354 
rect 90 354 93 357 
rect 90 357 93 360 
rect 90 360 93 363 
rect 90 363 93 366 
rect 90 366 93 369 
rect 90 369 93 372 
rect 90 372 93 375 
rect 90 375 93 378 
rect 90 378 93 381 
rect 90 381 93 384 
rect 90 384 93 387 
rect 90 387 93 390 
rect 90 390 93 393 
rect 90 393 93 396 
rect 90 396 93 399 
rect 90 399 93 402 
rect 90 402 93 405 
rect 90 405 93 408 
rect 90 408 93 411 
rect 90 411 93 414 
rect 90 414 93 417 
rect 90 417 93 420 
rect 90 420 93 423 
rect 90 423 93 426 
rect 90 426 93 429 
rect 90 429 93 432 
rect 90 432 93 435 
rect 90 435 93 438 
rect 90 438 93 441 
rect 90 441 93 444 
rect 90 444 93 447 
rect 90 447 93 450 
rect 90 450 93 453 
rect 90 453 93 456 
rect 90 456 93 459 
rect 90 459 93 462 
rect 90 462 93 465 
rect 90 465 93 468 
rect 90 468 93 471 
rect 90 471 93 474 
rect 90 474 93 477 
rect 90 477 93 480 
rect 90 480 93 483 
rect 90 483 93 486 
rect 90 486 93 489 
rect 90 489 93 492 
rect 90 492 93 495 
rect 90 495 93 498 
rect 90 498 93 501 
rect 90 501 93 504 
rect 90 504 93 507 
rect 90 507 93 510 
rect 93 0 96 3 
rect 93 3 96 6 
rect 93 6 96 9 
rect 93 9 96 12 
rect 93 12 96 15 
rect 93 15 96 18 
rect 93 18 96 21 
rect 93 21 96 24 
rect 93 24 96 27 
rect 93 27 96 30 
rect 93 30 96 33 
rect 93 33 96 36 
rect 93 36 96 39 
rect 93 39 96 42 
rect 93 42 96 45 
rect 93 45 96 48 
rect 93 48 96 51 
rect 93 51 96 54 
rect 93 54 96 57 
rect 93 57 96 60 
rect 93 60 96 63 
rect 93 63 96 66 
rect 93 66 96 69 
rect 93 69 96 72 
rect 93 72 96 75 
rect 93 75 96 78 
rect 93 78 96 81 
rect 93 84 96 87 
rect 93 87 96 90 
rect 93 90 96 93 
rect 93 93 96 96 
rect 93 96 96 99 
rect 93 99 96 102 
rect 93 102 96 105 
rect 93 105 96 108 
rect 93 108 96 111 
rect 93 111 96 114 
rect 93 114 96 117 
rect 93 117 96 120 
rect 93 120 96 123 
rect 93 123 96 126 
rect 93 126 96 129 
rect 93 129 96 132 
rect 93 132 96 135 
rect 93 135 96 138 
rect 93 138 96 141 
rect 93 141 96 144 
rect 93 144 96 147 
rect 93 147 96 150 
rect 93 150 96 153 
rect 93 153 96 156 
rect 93 156 96 159 
rect 93 159 96 162 
rect 93 162 96 165 
rect 93 165 96 168 
rect 93 168 96 171 
rect 93 171 96 174 
rect 93 174 96 177 
rect 93 177 96 180 
rect 93 180 96 183 
rect 93 183 96 186 
rect 93 186 96 189 
rect 93 189 96 192 
rect 93 192 96 195 
rect 93 195 96 198 
rect 93 198 96 201 
rect 93 201 96 204 
rect 93 204 96 207 
rect 93 207 96 210 
rect 93 210 96 213 
rect 93 213 96 216 
rect 93 216 96 219 
rect 93 219 96 222 
rect 93 222 96 225 
rect 93 225 96 228 
rect 93 228 96 231 
rect 93 231 96 234 
rect 93 234 96 237 
rect 93 237 96 240 
rect 93 240 96 243 
rect 93 243 96 246 
rect 93 246 96 249 
rect 93 249 96 252 
rect 93 252 96 255 
rect 93 255 96 258 
rect 93 258 96 261 
rect 93 261 96 264 
rect 93 264 96 267 
rect 93 267 96 270 
rect 93 270 96 273 
rect 93 273 96 276 
rect 93 276 96 279 
rect 93 279 96 282 
rect 93 282 96 285 
rect 93 285 96 288 
rect 93 288 96 291 
rect 93 291 96 294 
rect 93 294 96 297 
rect 93 297 96 300 
rect 93 300 96 303 
rect 93 303 96 306 
rect 93 306 96 309 
rect 93 309 96 312 
rect 93 312 96 315 
rect 93 315 96 318 
rect 93 318 96 321 
rect 93 324 96 327 
rect 93 327 96 330 
rect 93 333 96 336 
rect 93 336 96 339 
rect 93 339 96 342 
rect 93 342 96 345 
rect 93 345 96 348 
rect 93 348 96 351 
rect 93 351 96 354 
rect 93 354 96 357 
rect 93 357 96 360 
rect 93 360 96 363 
rect 93 363 96 366 
rect 93 366 96 369 
rect 93 369 96 372 
rect 93 372 96 375 
rect 93 375 96 378 
rect 93 378 96 381 
rect 93 381 96 384 
rect 93 384 96 387 
rect 93 387 96 390 
rect 93 390 96 393 
rect 93 393 96 396 
rect 93 396 96 399 
rect 93 399 96 402 
rect 93 402 96 405 
rect 93 405 96 408 
rect 93 408 96 411 
rect 93 411 96 414 
rect 93 414 96 417 
rect 93 420 96 423 
rect 93 423 96 426 
rect 93 426 96 429 
rect 93 429 96 432 
rect 93 432 96 435 
rect 93 435 96 438 
rect 93 438 96 441 
rect 93 441 96 444 
rect 93 444 96 447 
rect 93 447 96 450 
rect 93 450 96 453 
rect 93 453 96 456 
rect 93 456 96 459 
rect 93 459 96 462 
rect 93 462 96 465 
rect 93 468 96 471 
rect 93 471 96 474 
rect 93 477 96 480 
rect 93 480 96 483 
rect 93 483 96 486 
rect 93 486 96 489 
rect 93 489 96 492 
rect 93 492 96 495 
rect 93 495 96 498 
rect 93 498 96 501 
rect 93 501 96 504 
rect 93 504 96 507 
rect 93 507 96 510 
rect 96 0 99 3 
rect 96 3 99 6 
rect 96 6 99 9 
rect 96 9 99 12 
rect 96 12 99 15 
rect 96 15 99 18 
rect 96 18 99 21 
rect 96 21 99 24 
rect 96 24 99 27 
rect 96 27 99 30 
rect 96 30 99 33 
rect 96 33 99 36 
rect 96 36 99 39 
rect 96 39 99 42 
rect 96 42 99 45 
rect 96 45 99 48 
rect 96 48 99 51 
rect 96 51 99 54 
rect 96 54 99 57 
rect 96 57 99 60 
rect 96 60 99 63 
rect 96 63 99 66 
rect 96 66 99 69 
rect 96 69 99 72 
rect 96 72 99 75 
rect 96 75 99 78 
rect 96 78 99 81 
rect 96 81 99 84 
rect 96 84 99 87 
rect 96 87 99 90 
rect 96 90 99 93 
rect 96 93 99 96 
rect 96 96 99 99 
rect 96 99 99 102 
rect 96 102 99 105 
rect 96 105 99 108 
rect 96 108 99 111 
rect 96 111 99 114 
rect 96 114 99 117 
rect 96 117 99 120 
rect 96 120 99 123 
rect 96 123 99 126 
rect 96 126 99 129 
rect 96 129 99 132 
rect 96 132 99 135 
rect 96 135 99 138 
rect 96 138 99 141 
rect 96 141 99 144 
rect 96 144 99 147 
rect 96 147 99 150 
rect 96 150 99 153 
rect 96 153 99 156 
rect 96 156 99 159 
rect 96 159 99 162 
rect 96 162 99 165 
rect 96 165 99 168 
rect 96 168 99 171 
rect 96 171 99 174 
rect 96 174 99 177 
rect 96 177 99 180 
rect 96 180 99 183 
rect 96 183 99 186 
rect 96 186 99 189 
rect 96 189 99 192 
rect 96 192 99 195 
rect 96 195 99 198 
rect 96 198 99 201 
rect 96 201 99 204 
rect 96 204 99 207 
rect 96 207 99 210 
rect 96 210 99 213 
rect 96 213 99 216 
rect 96 216 99 219 
rect 96 219 99 222 
rect 96 222 99 225 
rect 96 225 99 228 
rect 96 228 99 231 
rect 96 231 99 234 
rect 96 234 99 237 
rect 96 237 99 240 
rect 96 240 99 243 
rect 96 243 99 246 
rect 96 246 99 249 
rect 96 249 99 252 
rect 96 252 99 255 
rect 96 255 99 258 
rect 96 258 99 261 
rect 96 261 99 264 
rect 96 264 99 267 
rect 96 267 99 270 
rect 96 270 99 273 
rect 96 273 99 276 
rect 96 276 99 279 
rect 96 279 99 282 
rect 96 282 99 285 
rect 96 285 99 288 
rect 96 288 99 291 
rect 96 291 99 294 
rect 96 294 99 297 
rect 96 297 99 300 
rect 96 300 99 303 
rect 96 303 99 306 
rect 96 306 99 309 
rect 96 309 99 312 
rect 96 312 99 315 
rect 96 315 99 318 
rect 96 318 99 321 
rect 96 321 99 324 
rect 96 324 99 327 
rect 96 327 99 330 
rect 96 330 99 333 
rect 96 333 99 336 
rect 96 336 99 339 
rect 96 339 99 342 
rect 96 342 99 345 
rect 96 345 99 348 
rect 96 348 99 351 
rect 96 351 99 354 
rect 96 354 99 357 
rect 96 357 99 360 
rect 96 360 99 363 
rect 96 363 99 366 
rect 96 366 99 369 
rect 96 369 99 372 
rect 96 372 99 375 
rect 96 375 99 378 
rect 96 378 99 381 
rect 96 381 99 384 
rect 96 384 99 387 
rect 96 387 99 390 
rect 96 390 99 393 
rect 96 393 99 396 
rect 96 396 99 399 
rect 96 399 99 402 
rect 96 402 99 405 
rect 96 405 99 408 
rect 96 408 99 411 
rect 96 411 99 414 
rect 96 414 99 417 
rect 96 417 99 420 
rect 96 420 99 423 
rect 96 423 99 426 
rect 96 426 99 429 
rect 96 429 99 432 
rect 96 432 99 435 
rect 96 435 99 438 
rect 96 438 99 441 
rect 96 441 99 444 
rect 96 444 99 447 
rect 96 447 99 450 
rect 96 450 99 453 
rect 96 453 99 456 
rect 96 456 99 459 
rect 96 459 99 462 
rect 96 462 99 465 
rect 96 465 99 468 
rect 96 468 99 471 
rect 96 471 99 474 
rect 96 474 99 477 
rect 96 477 99 480 
rect 96 480 99 483 
rect 96 483 99 486 
rect 96 486 99 489 
rect 96 489 99 492 
rect 96 492 99 495 
rect 96 495 99 498 
rect 96 498 99 501 
rect 96 501 99 504 
rect 96 504 99 507 
rect 96 507 99 510 
rect 99 0 102 3 
rect 99 3 102 6 
rect 99 6 102 9 
rect 99 9 102 12 
rect 99 12 102 15 
rect 99 15 102 18 
rect 99 18 102 21 
rect 99 21 102 24 
rect 99 24 102 27 
rect 99 27 102 30 
rect 99 30 102 33 
rect 99 33 102 36 
rect 99 36 102 39 
rect 99 39 102 42 
rect 99 42 102 45 
rect 99 45 102 48 
rect 99 48 102 51 
rect 99 51 102 54 
rect 99 54 102 57 
rect 99 57 102 60 
rect 99 60 102 63 
rect 99 63 102 66 
rect 99 66 102 69 
rect 99 69 102 72 
rect 99 72 102 75 
rect 99 75 102 78 
rect 99 78 102 81 
rect 99 81 102 84 
rect 99 84 102 87 
rect 99 87 102 90 
rect 99 90 102 93 
rect 99 93 102 96 
rect 99 96 102 99 
rect 99 99 102 102 
rect 99 102 102 105 
rect 99 105 102 108 
rect 99 108 102 111 
rect 99 111 102 114 
rect 99 114 102 117 
rect 99 117 102 120 
rect 99 120 102 123 
rect 99 123 102 126 
rect 99 126 102 129 
rect 99 129 102 132 
rect 99 132 102 135 
rect 99 135 102 138 
rect 99 138 102 141 
rect 99 141 102 144 
rect 99 144 102 147 
rect 99 147 102 150 
rect 99 150 102 153 
rect 99 153 102 156 
rect 99 156 102 159 
rect 99 159 102 162 
rect 99 162 102 165 
rect 99 165 102 168 
rect 99 168 102 171 
rect 99 171 102 174 
rect 99 174 102 177 
rect 99 177 102 180 
rect 99 180 102 183 
rect 99 183 102 186 
rect 99 186 102 189 
rect 99 189 102 192 
rect 99 192 102 195 
rect 99 195 102 198 
rect 99 198 102 201 
rect 99 201 102 204 
rect 99 204 102 207 
rect 99 207 102 210 
rect 99 210 102 213 
rect 99 213 102 216 
rect 99 216 102 219 
rect 99 219 102 222 
rect 99 222 102 225 
rect 99 225 102 228 
rect 99 228 102 231 
rect 99 231 102 234 
rect 99 234 102 237 
rect 99 237 102 240 
rect 99 240 102 243 
rect 99 243 102 246 
rect 99 246 102 249 
rect 99 249 102 252 
rect 99 252 102 255 
rect 99 255 102 258 
rect 99 258 102 261 
rect 99 261 102 264 
rect 99 264 102 267 
rect 99 267 102 270 
rect 99 270 102 273 
rect 99 273 102 276 
rect 99 276 102 279 
rect 99 279 102 282 
rect 99 282 102 285 
rect 99 285 102 288 
rect 99 288 102 291 
rect 99 291 102 294 
rect 99 294 102 297 
rect 99 297 102 300 
rect 99 300 102 303 
rect 99 303 102 306 
rect 99 306 102 309 
rect 99 309 102 312 
rect 99 312 102 315 
rect 99 315 102 318 
rect 99 318 102 321 
rect 99 321 102 324 
rect 99 324 102 327 
rect 99 327 102 330 
rect 99 330 102 333 
rect 99 333 102 336 
rect 99 336 102 339 
rect 99 339 102 342 
rect 99 342 102 345 
rect 99 345 102 348 
rect 99 348 102 351 
rect 99 351 102 354 
rect 99 354 102 357 
rect 99 357 102 360 
rect 99 360 102 363 
rect 99 363 102 366 
rect 99 366 102 369 
rect 99 369 102 372 
rect 99 372 102 375 
rect 99 375 102 378 
rect 99 378 102 381 
rect 99 381 102 384 
rect 99 384 102 387 
rect 99 387 102 390 
rect 99 390 102 393 
rect 99 393 102 396 
rect 99 396 102 399 
rect 99 399 102 402 
rect 99 402 102 405 
rect 99 405 102 408 
rect 99 408 102 411 
rect 99 411 102 414 
rect 99 414 102 417 
rect 99 417 102 420 
rect 99 420 102 423 
rect 99 423 102 426 
rect 99 426 102 429 
rect 99 429 102 432 
rect 99 432 102 435 
rect 99 435 102 438 
rect 99 438 102 441 
rect 99 441 102 444 
rect 99 444 102 447 
rect 99 447 102 450 
rect 99 450 102 453 
rect 99 453 102 456 
rect 99 456 102 459 
rect 99 459 102 462 
rect 99 462 102 465 
rect 99 465 102 468 
rect 99 468 102 471 
rect 99 471 102 474 
rect 99 474 102 477 
rect 99 477 102 480 
rect 99 480 102 483 
rect 99 483 102 486 
rect 99 486 102 489 
rect 99 489 102 492 
rect 99 492 102 495 
rect 99 495 102 498 
rect 99 498 102 501 
rect 99 501 102 504 
rect 99 504 102 507 
rect 99 507 102 510 
rect 102 0 105 3 
rect 102 3 105 6 
rect 102 6 105 9 
rect 102 9 105 12 
rect 102 12 105 15 
rect 102 15 105 18 
rect 102 18 105 21 
rect 102 21 105 24 
rect 102 24 105 27 
rect 102 27 105 30 
rect 102 30 105 33 
rect 102 33 105 36 
rect 102 36 105 39 
rect 102 39 105 42 
rect 102 42 105 45 
rect 102 45 105 48 
rect 102 48 105 51 
rect 102 51 105 54 
rect 102 54 105 57 
rect 102 57 105 60 
rect 102 60 105 63 
rect 102 63 105 66 
rect 102 66 105 69 
rect 102 69 105 72 
rect 102 72 105 75 
rect 102 75 105 78 
rect 102 78 105 81 
rect 102 81 105 84 
rect 102 84 105 87 
rect 102 87 105 90 
rect 102 90 105 93 
rect 102 93 105 96 
rect 102 96 105 99 
rect 102 99 105 102 
rect 102 102 105 105 
rect 102 105 105 108 
rect 102 108 105 111 
rect 102 111 105 114 
rect 102 114 105 117 
rect 102 117 105 120 
rect 102 120 105 123 
rect 102 123 105 126 
rect 102 126 105 129 
rect 102 129 105 132 
rect 102 132 105 135 
rect 102 135 105 138 
rect 102 138 105 141 
rect 102 141 105 144 
rect 102 144 105 147 
rect 102 147 105 150 
rect 102 150 105 153 
rect 102 153 105 156 
rect 102 156 105 159 
rect 102 159 105 162 
rect 102 162 105 165 
rect 102 165 105 168 
rect 102 168 105 171 
rect 102 171 105 174 
rect 102 174 105 177 
rect 102 177 105 180 
rect 102 180 105 183 
rect 102 183 105 186 
rect 102 186 105 189 
rect 102 189 105 192 
rect 102 192 105 195 
rect 102 195 105 198 
rect 102 198 105 201 
rect 102 201 105 204 
rect 102 204 105 207 
rect 102 207 105 210 
rect 102 210 105 213 
rect 102 213 105 216 
rect 102 216 105 219 
rect 102 219 105 222 
rect 102 222 105 225 
rect 102 225 105 228 
rect 102 228 105 231 
rect 102 231 105 234 
rect 102 234 105 237 
rect 102 237 105 240 
rect 102 240 105 243 
rect 102 243 105 246 
rect 102 246 105 249 
rect 102 249 105 252 
rect 102 252 105 255 
rect 102 255 105 258 
rect 102 258 105 261 
rect 102 261 105 264 
rect 102 264 105 267 
rect 102 267 105 270 
rect 102 270 105 273 
rect 102 273 105 276 
rect 102 276 105 279 
rect 102 279 105 282 
rect 102 282 105 285 
rect 102 285 105 288 
rect 102 288 105 291 
rect 102 291 105 294 
rect 102 294 105 297 
rect 102 297 105 300 
rect 102 300 105 303 
rect 102 303 105 306 
rect 102 306 105 309 
rect 102 309 105 312 
rect 102 312 105 315 
rect 102 315 105 318 
rect 102 318 105 321 
rect 102 321 105 324 
rect 102 324 105 327 
rect 102 327 105 330 
rect 102 330 105 333 
rect 102 333 105 336 
rect 102 336 105 339 
rect 102 339 105 342 
rect 102 342 105 345 
rect 102 345 105 348 
rect 102 348 105 351 
rect 102 351 105 354 
rect 102 354 105 357 
rect 102 357 105 360 
rect 102 360 105 363 
rect 102 363 105 366 
rect 102 366 105 369 
rect 102 369 105 372 
rect 102 372 105 375 
rect 102 375 105 378 
rect 102 378 105 381 
rect 102 381 105 384 
rect 102 384 105 387 
rect 102 387 105 390 
rect 102 390 105 393 
rect 102 393 105 396 
rect 102 396 105 399 
rect 102 399 105 402 
rect 102 402 105 405 
rect 102 405 105 408 
rect 102 408 105 411 
rect 102 411 105 414 
rect 102 414 105 417 
rect 102 417 105 420 
rect 102 420 105 423 
rect 102 423 105 426 
rect 102 426 105 429 
rect 102 429 105 432 
rect 102 432 105 435 
rect 102 435 105 438 
rect 102 438 105 441 
rect 102 441 105 444 
rect 102 444 105 447 
rect 102 447 105 450 
rect 102 450 105 453 
rect 102 453 105 456 
rect 102 456 105 459 
rect 102 459 105 462 
rect 102 462 105 465 
rect 102 465 105 468 
rect 102 468 105 471 
rect 102 471 105 474 
rect 102 474 105 477 
rect 102 477 105 480 
rect 102 480 105 483 
rect 102 483 105 486 
rect 102 486 105 489 
rect 102 489 105 492 
rect 102 492 105 495 
rect 102 495 105 498 
rect 102 498 105 501 
rect 102 501 105 504 
rect 102 504 105 507 
rect 102 507 105 510 
rect 105 0 108 3 
rect 105 3 108 6 
rect 105 6 108 9 
rect 105 9 108 12 
rect 105 12 108 15 
rect 105 15 108 18 
rect 105 18 108 21 
rect 105 21 108 24 
rect 105 24 108 27 
rect 105 27 108 30 
rect 105 30 108 33 
rect 105 33 108 36 
rect 105 36 108 39 
rect 105 39 108 42 
rect 105 42 108 45 
rect 105 45 108 48 
rect 105 48 108 51 
rect 105 51 108 54 
rect 105 54 108 57 
rect 105 57 108 60 
rect 105 60 108 63 
rect 105 63 108 66 
rect 105 66 108 69 
rect 105 69 108 72 
rect 105 72 108 75 
rect 105 75 108 78 
rect 105 78 108 81 
rect 105 81 108 84 
rect 105 84 108 87 
rect 105 87 108 90 
rect 105 90 108 93 
rect 105 93 108 96 
rect 105 96 108 99 
rect 105 99 108 102 
rect 105 102 108 105 
rect 105 105 108 108 
rect 105 108 108 111 
rect 105 111 108 114 
rect 105 114 108 117 
rect 105 117 108 120 
rect 105 120 108 123 
rect 105 123 108 126 
rect 105 126 108 129 
rect 105 129 108 132 
rect 105 132 108 135 
rect 105 135 108 138 
rect 105 138 108 141 
rect 105 141 108 144 
rect 105 144 108 147 
rect 105 147 108 150 
rect 105 150 108 153 
rect 105 153 108 156 
rect 105 156 108 159 
rect 105 159 108 162 
rect 105 162 108 165 
rect 105 165 108 168 
rect 105 168 108 171 
rect 105 171 108 174 
rect 105 174 108 177 
rect 105 177 108 180 
rect 105 180 108 183 
rect 105 183 108 186 
rect 105 186 108 189 
rect 105 189 108 192 
rect 105 192 108 195 
rect 105 195 108 198 
rect 105 198 108 201 
rect 105 201 108 204 
rect 105 204 108 207 
rect 105 207 108 210 
rect 105 210 108 213 
rect 105 213 108 216 
rect 105 216 108 219 
rect 105 219 108 222 
rect 105 222 108 225 
rect 105 225 108 228 
rect 105 228 108 231 
rect 105 231 108 234 
rect 105 234 108 237 
rect 105 237 108 240 
rect 105 240 108 243 
rect 105 243 108 246 
rect 105 246 108 249 
rect 105 249 108 252 
rect 105 252 108 255 
rect 105 255 108 258 
rect 105 258 108 261 
rect 105 261 108 264 
rect 105 264 108 267 
rect 105 267 108 270 
rect 105 270 108 273 
rect 105 273 108 276 
rect 105 276 108 279 
rect 105 279 108 282 
rect 105 282 108 285 
rect 105 285 108 288 
rect 105 288 108 291 
rect 105 291 108 294 
rect 105 294 108 297 
rect 105 297 108 300 
rect 105 300 108 303 
rect 105 303 108 306 
rect 105 306 108 309 
rect 105 309 108 312 
rect 105 312 108 315 
rect 105 315 108 318 
rect 105 318 108 321 
rect 105 321 108 324 
rect 105 324 108 327 
rect 105 327 108 330 
rect 105 330 108 333 
rect 105 333 108 336 
rect 105 336 108 339 
rect 105 339 108 342 
rect 105 342 108 345 
rect 105 345 108 348 
rect 105 348 108 351 
rect 105 351 108 354 
rect 105 354 108 357 
rect 105 357 108 360 
rect 105 360 108 363 
rect 105 363 108 366 
rect 105 366 108 369 
rect 105 369 108 372 
rect 105 372 108 375 
rect 105 375 108 378 
rect 105 378 108 381 
rect 105 381 108 384 
rect 105 384 108 387 
rect 105 387 108 390 
rect 105 390 108 393 
rect 105 393 108 396 
rect 105 396 108 399 
rect 105 399 108 402 
rect 105 402 108 405 
rect 105 405 108 408 
rect 105 408 108 411 
rect 105 411 108 414 
rect 105 414 108 417 
rect 105 417 108 420 
rect 105 420 108 423 
rect 105 423 108 426 
rect 105 426 108 429 
rect 105 429 108 432 
rect 105 432 108 435 
rect 105 435 108 438 
rect 105 438 108 441 
rect 105 441 108 444 
rect 105 444 108 447 
rect 105 447 108 450 
rect 105 450 108 453 
rect 105 453 108 456 
rect 105 456 108 459 
rect 105 459 108 462 
rect 105 462 108 465 
rect 105 465 108 468 
rect 105 468 108 471 
rect 105 471 108 474 
rect 105 474 108 477 
rect 105 477 108 480 
rect 105 480 108 483 
rect 105 483 108 486 
rect 105 486 108 489 
rect 105 489 108 492 
rect 105 492 108 495 
rect 105 495 108 498 
rect 105 498 108 501 
rect 105 501 108 504 
rect 105 504 108 507 
rect 105 507 108 510 
rect 108 0 111 3 
rect 108 3 111 6 
rect 108 6 111 9 
rect 108 9 111 12 
rect 108 12 111 15 
rect 108 15 111 18 
rect 108 18 111 21 
rect 108 21 111 24 
rect 108 24 111 27 
rect 108 27 111 30 
rect 108 30 111 33 
rect 108 33 111 36 
rect 108 36 111 39 
rect 108 39 111 42 
rect 108 42 111 45 
rect 108 45 111 48 
rect 108 48 111 51 
rect 108 51 111 54 
rect 108 54 111 57 
rect 108 57 111 60 
rect 108 60 111 63 
rect 108 63 111 66 
rect 108 66 111 69 
rect 108 69 111 72 
rect 108 72 111 75 
rect 108 75 111 78 
rect 108 78 111 81 
rect 108 81 111 84 
rect 108 84 111 87 
rect 108 87 111 90 
rect 108 90 111 93 
rect 108 93 111 96 
rect 108 96 111 99 
rect 108 99 111 102 
rect 108 102 111 105 
rect 108 105 111 108 
rect 108 108 111 111 
rect 108 111 111 114 
rect 108 114 111 117 
rect 108 117 111 120 
rect 108 120 111 123 
rect 108 123 111 126 
rect 108 126 111 129 
rect 108 129 111 132 
rect 108 132 111 135 
rect 108 135 111 138 
rect 108 138 111 141 
rect 108 141 111 144 
rect 108 144 111 147 
rect 108 147 111 150 
rect 108 150 111 153 
rect 108 153 111 156 
rect 108 156 111 159 
rect 108 159 111 162 
rect 108 162 111 165 
rect 108 165 111 168 
rect 108 168 111 171 
rect 108 171 111 174 
rect 108 174 111 177 
rect 108 177 111 180 
rect 108 180 111 183 
rect 108 183 111 186 
rect 108 186 111 189 
rect 108 189 111 192 
rect 108 192 111 195 
rect 108 195 111 198 
rect 108 198 111 201 
rect 108 201 111 204 
rect 108 204 111 207 
rect 108 207 111 210 
rect 108 210 111 213 
rect 108 213 111 216 
rect 108 216 111 219 
rect 108 219 111 222 
rect 108 222 111 225 
rect 108 225 111 228 
rect 108 228 111 231 
rect 108 231 111 234 
rect 108 234 111 237 
rect 108 237 111 240 
rect 108 240 111 243 
rect 108 243 111 246 
rect 108 246 111 249 
rect 108 249 111 252 
rect 108 252 111 255 
rect 108 255 111 258 
rect 108 258 111 261 
rect 108 261 111 264 
rect 108 264 111 267 
rect 108 267 111 270 
rect 108 270 111 273 
rect 108 273 111 276 
rect 108 276 111 279 
rect 108 279 111 282 
rect 108 282 111 285 
rect 108 285 111 288 
rect 108 288 111 291 
rect 108 291 111 294 
rect 108 294 111 297 
rect 108 297 111 300 
rect 108 300 111 303 
rect 108 303 111 306 
rect 108 306 111 309 
rect 108 309 111 312 
rect 108 312 111 315 
rect 108 315 111 318 
rect 108 318 111 321 
rect 108 321 111 324 
rect 108 324 111 327 
rect 108 327 111 330 
rect 108 330 111 333 
rect 108 333 111 336 
rect 108 336 111 339 
rect 108 339 111 342 
rect 108 342 111 345 
rect 108 345 111 348 
rect 108 348 111 351 
rect 108 351 111 354 
rect 108 354 111 357 
rect 108 357 111 360 
rect 108 360 111 363 
rect 108 363 111 366 
rect 108 366 111 369 
rect 108 369 111 372 
rect 108 372 111 375 
rect 108 375 111 378 
rect 108 378 111 381 
rect 108 381 111 384 
rect 108 384 111 387 
rect 108 387 111 390 
rect 108 390 111 393 
rect 108 393 111 396 
rect 108 396 111 399 
rect 108 399 111 402 
rect 108 402 111 405 
rect 108 405 111 408 
rect 108 408 111 411 
rect 108 411 111 414 
rect 108 414 111 417 
rect 108 417 111 420 
rect 108 420 111 423 
rect 108 423 111 426 
rect 108 426 111 429 
rect 108 429 111 432 
rect 108 432 111 435 
rect 108 435 111 438 
rect 108 438 111 441 
rect 108 441 111 444 
rect 108 444 111 447 
rect 108 447 111 450 
rect 108 450 111 453 
rect 108 453 111 456 
rect 108 456 111 459 
rect 108 459 111 462 
rect 108 462 111 465 
rect 108 465 111 468 
rect 108 468 111 471 
rect 108 471 111 474 
rect 108 474 111 477 
rect 108 477 111 480 
rect 108 480 111 483 
rect 108 483 111 486 
rect 108 486 111 489 
rect 108 489 111 492 
rect 108 492 111 495 
rect 108 495 111 498 
rect 108 498 111 501 
rect 108 501 111 504 
rect 108 504 111 507 
rect 108 507 111 510 
rect 111 0 114 3 
rect 111 3 114 6 
rect 111 6 114 9 
rect 111 9 114 12 
rect 111 12 114 15 
rect 111 15 114 18 
rect 111 18 114 21 
rect 111 21 114 24 
rect 111 24 114 27 
rect 111 27 114 30 
rect 111 30 114 33 
rect 111 33 114 36 
rect 111 36 114 39 
rect 111 39 114 42 
rect 111 42 114 45 
rect 111 45 114 48 
rect 111 48 114 51 
rect 111 51 114 54 
rect 111 54 114 57 
rect 111 57 114 60 
rect 111 60 114 63 
rect 111 63 114 66 
rect 111 66 114 69 
rect 111 69 114 72 
rect 111 72 114 75 
rect 111 75 114 78 
rect 111 78 114 81 
rect 111 81 114 84 
rect 111 84 114 87 
rect 111 87 114 90 
rect 111 90 114 93 
rect 111 93 114 96 
rect 111 96 114 99 
rect 111 99 114 102 
rect 111 102 114 105 
rect 111 105 114 108 
rect 111 108 114 111 
rect 111 111 114 114 
rect 111 114 114 117 
rect 111 117 114 120 
rect 111 120 114 123 
rect 111 123 114 126 
rect 111 126 114 129 
rect 111 129 114 132 
rect 111 132 114 135 
rect 111 135 114 138 
rect 111 138 114 141 
rect 111 141 114 144 
rect 111 144 114 147 
rect 111 147 114 150 
rect 111 150 114 153 
rect 111 153 114 156 
rect 111 156 114 159 
rect 111 159 114 162 
rect 111 162 114 165 
rect 111 165 114 168 
rect 111 168 114 171 
rect 111 171 114 174 
rect 111 174 114 177 
rect 111 177 114 180 
rect 111 180 114 183 
rect 111 183 114 186 
rect 111 186 114 189 
rect 111 189 114 192 
rect 111 192 114 195 
rect 111 195 114 198 
rect 111 198 114 201 
rect 111 201 114 204 
rect 111 204 114 207 
rect 111 207 114 210 
rect 111 210 114 213 
rect 111 213 114 216 
rect 111 216 114 219 
rect 111 219 114 222 
rect 111 222 114 225 
rect 111 225 114 228 
rect 111 228 114 231 
rect 111 231 114 234 
rect 111 234 114 237 
rect 111 237 114 240 
rect 111 240 114 243 
rect 111 243 114 246 
rect 111 246 114 249 
rect 111 249 114 252 
rect 111 252 114 255 
rect 111 255 114 258 
rect 111 258 114 261 
rect 111 261 114 264 
rect 111 264 114 267 
rect 111 267 114 270 
rect 111 270 114 273 
rect 111 273 114 276 
rect 111 276 114 279 
rect 111 279 114 282 
rect 111 282 114 285 
rect 111 285 114 288 
rect 111 288 114 291 
rect 111 291 114 294 
rect 111 294 114 297 
rect 111 297 114 300 
rect 111 300 114 303 
rect 111 303 114 306 
rect 111 306 114 309 
rect 111 309 114 312 
rect 111 312 114 315 
rect 111 315 114 318 
rect 111 318 114 321 
rect 111 321 114 324 
rect 111 324 114 327 
rect 111 327 114 330 
rect 111 330 114 333 
rect 111 333 114 336 
rect 111 336 114 339 
rect 111 339 114 342 
rect 111 342 114 345 
rect 111 345 114 348 
rect 111 348 114 351 
rect 111 351 114 354 
rect 111 354 114 357 
rect 111 357 114 360 
rect 111 360 114 363 
rect 111 363 114 366 
rect 111 366 114 369 
rect 111 369 114 372 
rect 111 372 114 375 
rect 111 375 114 378 
rect 111 378 114 381 
rect 111 381 114 384 
rect 111 384 114 387 
rect 111 387 114 390 
rect 111 390 114 393 
rect 111 393 114 396 
rect 111 396 114 399 
rect 111 399 114 402 
rect 111 402 114 405 
rect 111 405 114 408 
rect 111 408 114 411 
rect 111 411 114 414 
rect 111 414 114 417 
rect 111 417 114 420 
rect 111 420 114 423 
rect 111 423 114 426 
rect 111 426 114 429 
rect 111 429 114 432 
rect 111 432 114 435 
rect 111 435 114 438 
rect 111 438 114 441 
rect 111 441 114 444 
rect 111 444 114 447 
rect 111 447 114 450 
rect 111 450 114 453 
rect 111 453 114 456 
rect 111 456 114 459 
rect 111 459 114 462 
rect 111 462 114 465 
rect 111 465 114 468 
rect 111 468 114 471 
rect 111 471 114 474 
rect 111 474 114 477 
rect 111 477 114 480 
rect 111 480 114 483 
rect 111 483 114 486 
rect 111 486 114 489 
rect 111 489 114 492 
rect 111 492 114 495 
rect 111 495 114 498 
rect 111 498 114 501 
rect 111 501 114 504 
rect 111 504 114 507 
rect 111 507 114 510 
rect 114 0 117 3 
rect 114 3 117 6 
rect 114 6 117 9 
rect 114 9 117 12 
rect 114 12 117 15 
rect 114 15 117 18 
rect 114 18 117 21 
rect 114 21 117 24 
rect 114 24 117 27 
rect 114 27 117 30 
rect 114 30 117 33 
rect 114 33 117 36 
rect 114 36 117 39 
rect 114 39 117 42 
rect 114 42 117 45 
rect 114 45 117 48 
rect 114 48 117 51 
rect 114 51 117 54 
rect 114 54 117 57 
rect 114 57 117 60 
rect 114 60 117 63 
rect 114 63 117 66 
rect 114 66 117 69 
rect 114 69 117 72 
rect 114 72 117 75 
rect 114 75 117 78 
rect 114 78 117 81 
rect 114 81 117 84 
rect 114 84 117 87 
rect 114 87 117 90 
rect 114 90 117 93 
rect 114 93 117 96 
rect 114 96 117 99 
rect 114 99 117 102 
rect 114 102 117 105 
rect 114 105 117 108 
rect 114 108 117 111 
rect 114 111 117 114 
rect 114 114 117 117 
rect 114 117 117 120 
rect 114 120 117 123 
rect 114 123 117 126 
rect 114 126 117 129 
rect 114 129 117 132 
rect 114 132 117 135 
rect 114 135 117 138 
rect 114 138 117 141 
rect 114 141 117 144 
rect 114 144 117 147 
rect 114 147 117 150 
rect 114 150 117 153 
rect 114 153 117 156 
rect 114 156 117 159 
rect 114 159 117 162 
rect 114 162 117 165 
rect 114 165 117 168 
rect 114 168 117 171 
rect 114 171 117 174 
rect 114 174 117 177 
rect 114 177 117 180 
rect 114 180 117 183 
rect 114 183 117 186 
rect 114 186 117 189 
rect 114 189 117 192 
rect 114 192 117 195 
rect 114 195 117 198 
rect 114 198 117 201 
rect 114 201 117 204 
rect 114 204 117 207 
rect 114 207 117 210 
rect 114 210 117 213 
rect 114 213 117 216 
rect 114 216 117 219 
rect 114 219 117 222 
rect 114 222 117 225 
rect 114 225 117 228 
rect 114 228 117 231 
rect 114 231 117 234 
rect 114 234 117 237 
rect 114 237 117 240 
rect 114 240 117 243 
rect 114 243 117 246 
rect 114 246 117 249 
rect 114 249 117 252 
rect 114 252 117 255 
rect 114 255 117 258 
rect 114 258 117 261 
rect 114 261 117 264 
rect 114 264 117 267 
rect 114 267 117 270 
rect 114 270 117 273 
rect 114 273 117 276 
rect 114 276 117 279 
rect 114 279 117 282 
rect 114 282 117 285 
rect 114 285 117 288 
rect 114 288 117 291 
rect 114 291 117 294 
rect 114 294 117 297 
rect 114 297 117 300 
rect 114 300 117 303 
rect 114 303 117 306 
rect 114 306 117 309 
rect 114 309 117 312 
rect 114 312 117 315 
rect 114 315 117 318 
rect 114 318 117 321 
rect 114 321 117 324 
rect 114 324 117 327 
rect 114 327 117 330 
rect 114 330 117 333 
rect 114 333 117 336 
rect 114 336 117 339 
rect 114 339 117 342 
rect 114 342 117 345 
rect 114 345 117 348 
rect 114 348 117 351 
rect 114 351 117 354 
rect 114 354 117 357 
rect 114 357 117 360 
rect 114 360 117 363 
rect 114 363 117 366 
rect 114 366 117 369 
rect 114 369 117 372 
rect 114 372 117 375 
rect 114 375 117 378 
rect 114 378 117 381 
rect 114 381 117 384 
rect 114 384 117 387 
rect 114 387 117 390 
rect 114 390 117 393 
rect 114 393 117 396 
rect 114 396 117 399 
rect 114 399 117 402 
rect 114 402 117 405 
rect 114 405 117 408 
rect 114 408 117 411 
rect 114 411 117 414 
rect 114 414 117 417 
rect 114 417 117 420 
rect 114 420 117 423 
rect 114 423 117 426 
rect 114 426 117 429 
rect 114 429 117 432 
rect 114 432 117 435 
rect 114 435 117 438 
rect 114 438 117 441 
rect 114 441 117 444 
rect 114 444 117 447 
rect 114 447 117 450 
rect 114 450 117 453 
rect 114 453 117 456 
rect 114 456 117 459 
rect 114 459 117 462 
rect 114 462 117 465 
rect 114 465 117 468 
rect 114 468 117 471 
rect 114 471 117 474 
rect 114 474 117 477 
rect 114 477 117 480 
rect 114 480 117 483 
rect 114 483 117 486 
rect 114 486 117 489 
rect 114 489 117 492 
rect 114 492 117 495 
rect 114 495 117 498 
rect 114 498 117 501 
rect 114 501 117 504 
rect 114 504 117 507 
rect 114 507 117 510 
rect 117 0 120 3 
rect 117 3 120 6 
rect 117 6 120 9 
rect 117 9 120 12 
rect 117 12 120 15 
rect 117 15 120 18 
rect 117 18 120 21 
rect 117 21 120 24 
rect 117 24 120 27 
rect 117 27 120 30 
rect 117 30 120 33 
rect 117 33 120 36 
rect 117 36 120 39 
rect 117 39 120 42 
rect 117 42 120 45 
rect 117 45 120 48 
rect 117 48 120 51 
rect 117 51 120 54 
rect 117 54 120 57 
rect 117 57 120 60 
rect 117 60 120 63 
rect 117 63 120 66 
rect 117 66 120 69 
rect 117 69 120 72 
rect 117 72 120 75 
rect 117 75 120 78 
rect 117 78 120 81 
rect 117 81 120 84 
rect 117 84 120 87 
rect 117 87 120 90 
rect 117 90 120 93 
rect 117 93 120 96 
rect 117 96 120 99 
rect 117 99 120 102 
rect 117 102 120 105 
rect 117 105 120 108 
rect 117 108 120 111 
rect 117 111 120 114 
rect 117 114 120 117 
rect 117 117 120 120 
rect 117 120 120 123 
rect 117 123 120 126 
rect 117 126 120 129 
rect 117 129 120 132 
rect 117 132 120 135 
rect 117 135 120 138 
rect 117 138 120 141 
rect 117 141 120 144 
rect 117 144 120 147 
rect 117 147 120 150 
rect 117 150 120 153 
rect 117 153 120 156 
rect 117 156 120 159 
rect 117 159 120 162 
rect 117 162 120 165 
rect 117 165 120 168 
rect 117 168 120 171 
rect 117 171 120 174 
rect 117 174 120 177 
rect 117 177 120 180 
rect 117 180 120 183 
rect 117 183 120 186 
rect 117 186 120 189 
rect 117 189 120 192 
rect 117 192 120 195 
rect 117 195 120 198 
rect 117 198 120 201 
rect 117 201 120 204 
rect 117 204 120 207 
rect 117 207 120 210 
rect 117 210 120 213 
rect 117 213 120 216 
rect 117 216 120 219 
rect 117 219 120 222 
rect 117 222 120 225 
rect 117 225 120 228 
rect 117 228 120 231 
rect 117 231 120 234 
rect 117 234 120 237 
rect 117 237 120 240 
rect 117 240 120 243 
rect 117 243 120 246 
rect 117 246 120 249 
rect 117 249 120 252 
rect 117 252 120 255 
rect 117 255 120 258 
rect 117 258 120 261 
rect 117 261 120 264 
rect 117 264 120 267 
rect 117 267 120 270 
rect 117 270 120 273 
rect 117 273 120 276 
rect 117 276 120 279 
rect 117 279 120 282 
rect 117 282 120 285 
rect 117 285 120 288 
rect 117 288 120 291 
rect 117 291 120 294 
rect 117 294 120 297 
rect 117 297 120 300 
rect 117 300 120 303 
rect 117 303 120 306 
rect 117 306 120 309 
rect 117 309 120 312 
rect 117 312 120 315 
rect 117 315 120 318 
rect 117 318 120 321 
rect 117 321 120 324 
rect 117 324 120 327 
rect 117 327 120 330 
rect 117 330 120 333 
rect 117 333 120 336 
rect 117 336 120 339 
rect 117 339 120 342 
rect 117 342 120 345 
rect 117 345 120 348 
rect 117 348 120 351 
rect 117 351 120 354 
rect 117 354 120 357 
rect 117 357 120 360 
rect 117 360 120 363 
rect 117 363 120 366 
rect 117 366 120 369 
rect 117 369 120 372 
rect 117 372 120 375 
rect 117 375 120 378 
rect 117 378 120 381 
rect 117 381 120 384 
rect 117 384 120 387 
rect 117 387 120 390 
rect 117 390 120 393 
rect 117 393 120 396 
rect 117 396 120 399 
rect 117 399 120 402 
rect 117 402 120 405 
rect 117 405 120 408 
rect 117 408 120 411 
rect 117 411 120 414 
rect 117 414 120 417 
rect 117 417 120 420 
rect 117 420 120 423 
rect 117 423 120 426 
rect 117 426 120 429 
rect 117 429 120 432 
rect 117 432 120 435 
rect 117 435 120 438 
rect 117 438 120 441 
rect 117 441 120 444 
rect 117 444 120 447 
rect 117 447 120 450 
rect 117 450 120 453 
rect 117 453 120 456 
rect 117 456 120 459 
rect 117 459 120 462 
rect 117 462 120 465 
rect 117 465 120 468 
rect 117 468 120 471 
rect 117 471 120 474 
rect 117 474 120 477 
rect 117 477 120 480 
rect 117 480 120 483 
rect 117 483 120 486 
rect 117 486 120 489 
rect 117 489 120 492 
rect 117 492 120 495 
rect 117 495 120 498 
rect 117 498 120 501 
rect 117 501 120 504 
rect 117 504 120 507 
rect 117 507 120 510 
rect 120 0 123 3 
rect 120 3 123 6 
rect 120 6 123 9 
rect 120 9 123 12 
rect 120 12 123 15 
rect 120 15 123 18 
rect 120 18 123 21 
rect 120 21 123 24 
rect 120 24 123 27 
rect 120 27 123 30 
rect 120 30 123 33 
rect 120 33 123 36 
rect 120 36 123 39 
rect 120 39 123 42 
rect 120 42 123 45 
rect 120 45 123 48 
rect 120 48 123 51 
rect 120 51 123 54 
rect 120 54 123 57 
rect 120 57 123 60 
rect 120 60 123 63 
rect 120 63 123 66 
rect 120 66 123 69 
rect 120 69 123 72 
rect 120 72 123 75 
rect 120 75 123 78 
rect 120 78 123 81 
rect 120 81 123 84 
rect 120 84 123 87 
rect 120 87 123 90 
rect 120 90 123 93 
rect 120 93 123 96 
rect 120 96 123 99 
rect 120 99 123 102 
rect 120 102 123 105 
rect 120 105 123 108 
rect 120 108 123 111 
rect 120 111 123 114 
rect 120 114 123 117 
rect 120 117 123 120 
rect 120 120 123 123 
rect 120 123 123 126 
rect 120 126 123 129 
rect 120 129 123 132 
rect 120 132 123 135 
rect 120 135 123 138 
rect 120 138 123 141 
rect 120 141 123 144 
rect 120 144 123 147 
rect 120 147 123 150 
rect 120 150 123 153 
rect 120 153 123 156 
rect 120 156 123 159 
rect 120 159 123 162 
rect 120 162 123 165 
rect 120 165 123 168 
rect 120 168 123 171 
rect 120 171 123 174 
rect 120 174 123 177 
rect 120 177 123 180 
rect 120 180 123 183 
rect 120 183 123 186 
rect 120 186 123 189 
rect 120 189 123 192 
rect 120 192 123 195 
rect 120 195 123 198 
rect 120 198 123 201 
rect 120 201 123 204 
rect 120 204 123 207 
rect 120 207 123 210 
rect 120 210 123 213 
rect 120 213 123 216 
rect 120 216 123 219 
rect 120 219 123 222 
rect 120 222 123 225 
rect 120 225 123 228 
rect 120 228 123 231 
rect 120 231 123 234 
rect 120 234 123 237 
rect 120 237 123 240 
rect 120 240 123 243 
rect 120 243 123 246 
rect 120 246 123 249 
rect 120 249 123 252 
rect 120 252 123 255 
rect 120 255 123 258 
rect 120 258 123 261 
rect 120 261 123 264 
rect 120 264 123 267 
rect 120 267 123 270 
rect 120 270 123 273 
rect 120 273 123 276 
rect 120 276 123 279 
rect 120 279 123 282 
rect 120 282 123 285 
rect 120 285 123 288 
rect 120 288 123 291 
rect 120 291 123 294 
rect 120 294 123 297 
rect 120 297 123 300 
rect 120 300 123 303 
rect 120 303 123 306 
rect 120 306 123 309 
rect 120 309 123 312 
rect 120 312 123 315 
rect 120 315 123 318 
rect 120 318 123 321 
rect 120 321 123 324 
rect 120 324 123 327 
rect 120 327 123 330 
rect 120 330 123 333 
rect 120 333 123 336 
rect 120 336 123 339 
rect 120 339 123 342 
rect 120 342 123 345 
rect 120 345 123 348 
rect 120 348 123 351 
rect 120 351 123 354 
rect 120 354 123 357 
rect 120 357 123 360 
rect 120 360 123 363 
rect 120 363 123 366 
rect 120 366 123 369 
rect 120 369 123 372 
rect 120 372 123 375 
rect 120 375 123 378 
rect 120 378 123 381 
rect 120 381 123 384 
rect 120 384 123 387 
rect 120 387 123 390 
rect 120 390 123 393 
rect 120 393 123 396 
rect 120 396 123 399 
rect 120 399 123 402 
rect 120 402 123 405 
rect 120 405 123 408 
rect 120 408 123 411 
rect 120 411 123 414 
rect 120 414 123 417 
rect 120 417 123 420 
rect 120 420 123 423 
rect 120 423 123 426 
rect 120 426 123 429 
rect 120 429 123 432 
rect 120 432 123 435 
rect 120 435 123 438 
rect 120 438 123 441 
rect 120 441 123 444 
rect 120 444 123 447 
rect 120 447 123 450 
rect 120 450 123 453 
rect 120 453 123 456 
rect 120 456 123 459 
rect 120 459 123 462 
rect 120 462 123 465 
rect 120 465 123 468 
rect 120 468 123 471 
rect 120 471 123 474 
rect 120 474 123 477 
rect 120 477 123 480 
rect 120 480 123 483 
rect 120 483 123 486 
rect 120 486 123 489 
rect 120 489 123 492 
rect 120 492 123 495 
rect 120 495 123 498 
rect 120 498 123 501 
rect 120 501 123 504 
rect 120 504 123 507 
rect 120 507 123 510 
rect 123 0 126 3 
rect 123 3 126 6 
rect 123 6 126 9 
rect 123 9 126 12 
rect 123 12 126 15 
rect 123 15 126 18 
rect 123 18 126 21 
rect 123 21 126 24 
rect 123 24 126 27 
rect 123 27 126 30 
rect 123 30 126 33 
rect 123 33 126 36 
rect 123 36 126 39 
rect 123 39 126 42 
rect 123 42 126 45 
rect 123 45 126 48 
rect 123 48 126 51 
rect 123 51 126 54 
rect 123 54 126 57 
rect 123 57 126 60 
rect 123 60 126 63 
rect 123 63 126 66 
rect 123 66 126 69 
rect 123 69 126 72 
rect 123 72 126 75 
rect 123 75 126 78 
rect 123 78 126 81 
rect 123 81 126 84 
rect 123 84 126 87 
rect 123 87 126 90 
rect 123 90 126 93 
rect 123 93 126 96 
rect 123 96 126 99 
rect 123 99 126 102 
rect 123 102 126 105 
rect 123 105 126 108 
rect 123 108 126 111 
rect 123 111 126 114 
rect 123 114 126 117 
rect 123 117 126 120 
rect 123 120 126 123 
rect 123 123 126 126 
rect 123 126 126 129 
rect 123 129 126 132 
rect 123 132 126 135 
rect 123 135 126 138 
rect 123 138 126 141 
rect 123 141 126 144 
rect 123 144 126 147 
rect 123 147 126 150 
rect 123 150 126 153 
rect 123 153 126 156 
rect 123 156 126 159 
rect 123 159 126 162 
rect 123 162 126 165 
rect 123 165 126 168 
rect 123 168 126 171 
rect 123 171 126 174 
rect 123 174 126 177 
rect 123 177 126 180 
rect 123 180 126 183 
rect 123 183 126 186 
rect 123 186 126 189 
rect 123 189 126 192 
rect 123 192 126 195 
rect 123 195 126 198 
rect 123 198 126 201 
rect 123 201 126 204 
rect 123 204 126 207 
rect 123 207 126 210 
rect 123 210 126 213 
rect 123 213 126 216 
rect 123 216 126 219 
rect 123 219 126 222 
rect 123 222 126 225 
rect 123 225 126 228 
rect 123 228 126 231 
rect 123 231 126 234 
rect 123 234 126 237 
rect 123 237 126 240 
rect 123 240 126 243 
rect 123 243 126 246 
rect 123 246 126 249 
rect 123 249 126 252 
rect 123 252 126 255 
rect 123 255 126 258 
rect 123 258 126 261 
rect 123 261 126 264 
rect 123 264 126 267 
rect 123 267 126 270 
rect 123 270 126 273 
rect 123 273 126 276 
rect 123 276 126 279 
rect 123 279 126 282 
rect 123 282 126 285 
rect 123 285 126 288 
rect 123 288 126 291 
rect 123 291 126 294 
rect 123 294 126 297 
rect 123 297 126 300 
rect 123 300 126 303 
rect 123 303 126 306 
rect 123 306 126 309 
rect 123 309 126 312 
rect 123 312 126 315 
rect 123 315 126 318 
rect 123 318 126 321 
rect 123 321 126 324 
rect 123 324 126 327 
rect 123 327 126 330 
rect 123 330 126 333 
rect 123 333 126 336 
rect 123 336 126 339 
rect 123 339 126 342 
rect 123 342 126 345 
rect 123 345 126 348 
rect 123 348 126 351 
rect 123 351 126 354 
rect 123 354 126 357 
rect 123 357 126 360 
rect 123 360 126 363 
rect 123 363 126 366 
rect 123 366 126 369 
rect 123 369 126 372 
rect 123 372 126 375 
rect 123 375 126 378 
rect 123 378 126 381 
rect 123 381 126 384 
rect 123 384 126 387 
rect 123 387 126 390 
rect 123 390 126 393 
rect 123 393 126 396 
rect 123 396 126 399 
rect 123 399 126 402 
rect 123 402 126 405 
rect 123 405 126 408 
rect 123 408 126 411 
rect 123 411 126 414 
rect 123 414 126 417 
rect 123 417 126 420 
rect 123 420 126 423 
rect 123 423 126 426 
rect 123 426 126 429 
rect 123 429 126 432 
rect 123 432 126 435 
rect 123 435 126 438 
rect 123 438 126 441 
rect 123 441 126 444 
rect 123 444 126 447 
rect 123 447 126 450 
rect 123 450 126 453 
rect 123 453 126 456 
rect 123 456 126 459 
rect 123 459 126 462 
rect 123 462 126 465 
rect 123 465 126 468 
rect 123 468 126 471 
rect 123 471 126 474 
rect 123 474 126 477 
rect 123 477 126 480 
rect 123 480 126 483 
rect 123 483 126 486 
rect 123 486 126 489 
rect 123 489 126 492 
rect 123 492 126 495 
rect 123 495 126 498 
rect 123 498 126 501 
rect 123 501 126 504 
rect 123 504 126 507 
rect 123 507 126 510 
rect 126 0 129 3 
rect 126 3 129 6 
rect 126 6 129 9 
rect 126 9 129 12 
rect 126 12 129 15 
rect 126 15 129 18 
rect 126 18 129 21 
rect 126 21 129 24 
rect 126 24 129 27 
rect 126 27 129 30 
rect 126 30 129 33 
rect 126 33 129 36 
rect 126 36 129 39 
rect 126 39 129 42 
rect 126 42 129 45 
rect 126 45 129 48 
rect 126 48 129 51 
rect 126 51 129 54 
rect 126 54 129 57 
rect 126 57 129 60 
rect 126 60 129 63 
rect 126 63 129 66 
rect 126 66 129 69 
rect 126 69 129 72 
rect 126 72 129 75 
rect 126 75 129 78 
rect 126 78 129 81 
rect 126 84 129 87 
rect 126 87 129 90 
rect 126 90 129 93 
rect 126 93 129 96 
rect 126 96 129 99 
rect 126 99 129 102 
rect 126 102 129 105 
rect 126 105 129 108 
rect 126 108 129 111 
rect 126 111 129 114 
rect 126 114 129 117 
rect 126 117 129 120 
rect 126 120 129 123 
rect 126 123 129 126 
rect 126 126 129 129 
rect 126 129 129 132 
rect 126 132 129 135 
rect 126 135 129 138 
rect 126 138 129 141 
rect 126 141 129 144 
rect 126 144 129 147 
rect 126 147 129 150 
rect 126 150 129 153 
rect 126 153 129 156 
rect 126 156 129 159 
rect 126 159 129 162 
rect 126 162 129 165 
rect 126 165 129 168 
rect 126 168 129 171 
rect 126 171 129 174 
rect 126 174 129 177 
rect 126 177 129 180 
rect 126 180 129 183 
rect 126 183 129 186 
rect 126 186 129 189 
rect 126 189 129 192 
rect 126 192 129 195 
rect 126 195 129 198 
rect 126 198 129 201 
rect 126 201 129 204 
rect 126 204 129 207 
rect 126 207 129 210 
rect 126 210 129 213 
rect 126 213 129 216 
rect 126 216 129 219 
rect 126 219 129 222 
rect 126 222 129 225 
rect 126 225 129 228 
rect 126 228 129 231 
rect 126 231 129 234 
rect 126 234 129 237 
rect 126 237 129 240 
rect 126 240 129 243 
rect 126 243 129 246 
rect 126 246 129 249 
rect 126 249 129 252 
rect 126 252 129 255 
rect 126 255 129 258 
rect 126 258 129 261 
rect 126 261 129 264 
rect 126 264 129 267 
rect 126 267 129 270 
rect 126 270 129 273 
rect 126 273 129 276 
rect 126 276 129 279 
rect 126 279 129 282 
rect 126 282 129 285 
rect 126 285 129 288 
rect 126 288 129 291 
rect 126 291 129 294 
rect 126 294 129 297 
rect 126 297 129 300 
rect 126 300 129 303 
rect 126 303 129 306 
rect 126 306 129 309 
rect 126 309 129 312 
rect 126 312 129 315 
rect 126 315 129 318 
rect 126 318 129 321 
rect 126 321 129 324 
rect 126 324 129 327 
rect 126 327 129 330 
rect 126 330 129 333 
rect 126 333 129 336 
rect 126 336 129 339 
rect 126 339 129 342 
rect 126 342 129 345 
rect 126 345 129 348 
rect 126 348 129 351 
rect 126 351 129 354 
rect 126 354 129 357 
rect 126 357 129 360 
rect 126 360 129 363 
rect 126 363 129 366 
rect 126 366 129 369 
rect 126 369 129 372 
rect 126 372 129 375 
rect 126 375 129 378 
rect 126 378 129 381 
rect 126 381 129 384 
rect 126 384 129 387 
rect 126 387 129 390 
rect 126 390 129 393 
rect 126 393 129 396 
rect 126 396 129 399 
rect 126 399 129 402 
rect 126 402 129 405 
rect 126 405 129 408 
rect 126 408 129 411 
rect 126 411 129 414 
rect 126 414 129 417 
rect 126 420 129 423 
rect 126 423 129 426 
rect 126 429 129 432 
rect 126 432 129 435 
rect 126 435 129 438 
rect 126 438 129 441 
rect 126 441 129 444 
rect 126 444 129 447 
rect 126 447 129 450 
rect 126 450 129 453 
rect 126 453 129 456 
rect 126 456 129 459 
rect 126 459 129 462 
rect 126 462 129 465 
rect 126 465 129 468 
rect 126 468 129 471 
rect 126 471 129 474 
rect 126 474 129 477 
rect 126 477 129 480 
rect 126 480 129 483 
rect 126 483 129 486 
rect 126 486 129 489 
rect 126 489 129 492 
rect 126 492 129 495 
rect 126 495 129 498 
rect 126 498 129 501 
rect 126 501 129 504 
rect 126 504 129 507 
rect 126 507 129 510 
rect 129 0 132 3 
rect 129 3 132 6 
rect 129 6 132 9 
rect 129 9 132 12 
rect 129 12 132 15 
rect 129 15 132 18 
rect 129 18 132 21 
rect 129 21 132 24 
rect 129 24 132 27 
rect 129 27 132 30 
rect 129 30 132 33 
rect 129 33 132 36 
rect 129 36 132 39 
rect 129 39 132 42 
rect 129 42 132 45 
rect 129 45 132 48 
rect 129 48 132 51 
rect 129 51 132 54 
rect 129 54 132 57 
rect 129 57 132 60 
rect 129 60 132 63 
rect 129 63 132 66 
rect 129 66 132 69 
rect 129 69 132 72 
rect 129 72 132 75 
rect 129 75 132 78 
rect 129 78 132 81 
rect 129 81 132 84 
rect 129 84 132 87 
rect 129 87 132 90 
rect 129 90 132 93 
rect 129 93 132 96 
rect 129 96 132 99 
rect 129 99 132 102 
rect 129 102 132 105 
rect 129 105 132 108 
rect 129 108 132 111 
rect 129 111 132 114 
rect 129 114 132 117 
rect 129 117 132 120 
rect 129 120 132 123 
rect 129 123 132 126 
rect 129 126 132 129 
rect 129 129 132 132 
rect 129 132 132 135 
rect 129 135 132 138 
rect 129 138 132 141 
rect 129 141 132 144 
rect 129 144 132 147 
rect 129 147 132 150 
rect 129 150 132 153 
rect 129 153 132 156 
rect 129 156 132 159 
rect 129 159 132 162 
rect 129 162 132 165 
rect 129 165 132 168 
rect 129 168 132 171 
rect 129 171 132 174 
rect 129 174 132 177 
rect 129 177 132 180 
rect 129 180 132 183 
rect 129 183 132 186 
rect 129 186 132 189 
rect 129 189 132 192 
rect 129 192 132 195 
rect 129 195 132 198 
rect 129 198 132 201 
rect 129 201 132 204 
rect 129 204 132 207 
rect 129 207 132 210 
rect 129 210 132 213 
rect 129 213 132 216 
rect 129 216 132 219 
rect 129 219 132 222 
rect 129 222 132 225 
rect 129 225 132 228 
rect 129 228 132 231 
rect 129 231 132 234 
rect 129 234 132 237 
rect 129 237 132 240 
rect 129 240 132 243 
rect 129 243 132 246 
rect 129 246 132 249 
rect 129 249 132 252 
rect 129 252 132 255 
rect 129 255 132 258 
rect 129 258 132 261 
rect 129 261 132 264 
rect 129 264 132 267 
rect 129 267 132 270 
rect 129 270 132 273 
rect 129 273 132 276 
rect 129 276 132 279 
rect 129 279 132 282 
rect 129 282 132 285 
rect 129 285 132 288 
rect 129 288 132 291 
rect 129 291 132 294 
rect 129 294 132 297 
rect 129 297 132 300 
rect 129 300 132 303 
rect 129 303 132 306 
rect 129 306 132 309 
rect 129 309 132 312 
rect 129 312 132 315 
rect 129 315 132 318 
rect 129 318 132 321 
rect 129 321 132 324 
rect 129 324 132 327 
rect 129 327 132 330 
rect 129 330 132 333 
rect 129 333 132 336 
rect 129 336 132 339 
rect 129 339 132 342 
rect 129 342 132 345 
rect 129 345 132 348 
rect 129 348 132 351 
rect 129 351 132 354 
rect 129 354 132 357 
rect 129 357 132 360 
rect 129 360 132 363 
rect 129 363 132 366 
rect 129 366 132 369 
rect 129 369 132 372 
rect 129 372 132 375 
rect 129 375 132 378 
rect 129 378 132 381 
rect 129 381 132 384 
rect 129 384 132 387 
rect 129 387 132 390 
rect 129 390 132 393 
rect 129 393 132 396 
rect 129 396 132 399 
rect 129 399 132 402 
rect 129 402 132 405 
rect 129 405 132 408 
rect 129 408 132 411 
rect 129 411 132 414 
rect 129 414 132 417 
rect 129 417 132 420 
rect 129 420 132 423 
rect 129 423 132 426 
rect 129 426 132 429 
rect 129 429 132 432 
rect 129 432 132 435 
rect 129 435 132 438 
rect 129 438 132 441 
rect 129 441 132 444 
rect 129 444 132 447 
rect 129 447 132 450 
rect 129 450 132 453 
rect 129 453 132 456 
rect 129 456 132 459 
rect 129 459 132 462 
rect 129 462 132 465 
rect 129 465 132 468 
rect 129 468 132 471 
rect 129 471 132 474 
rect 129 474 132 477 
rect 129 477 132 480 
rect 129 480 132 483 
rect 129 483 132 486 
rect 129 486 132 489 
rect 129 489 132 492 
rect 129 492 132 495 
rect 129 495 132 498 
rect 129 498 132 501 
rect 129 501 132 504 
rect 129 504 132 507 
rect 129 507 132 510 
rect 132 0 135 3 
rect 132 3 135 6 
rect 132 6 135 9 
rect 132 9 135 12 
rect 132 12 135 15 
rect 132 15 135 18 
rect 132 18 135 21 
rect 132 21 135 24 
rect 132 24 135 27 
rect 132 27 135 30 
rect 132 30 135 33 
rect 132 33 135 36 
rect 132 36 135 39 
rect 132 39 135 42 
rect 132 42 135 45 
rect 132 45 135 48 
rect 132 48 135 51 
rect 132 51 135 54 
rect 132 54 135 57 
rect 132 57 135 60 
rect 132 60 135 63 
rect 132 63 135 66 
rect 132 66 135 69 
rect 132 69 135 72 
rect 132 72 135 75 
rect 132 75 135 78 
rect 132 78 135 81 
rect 132 81 135 84 
rect 132 84 135 87 
rect 132 87 135 90 
rect 132 90 135 93 
rect 132 93 135 96 
rect 132 96 135 99 
rect 132 99 135 102 
rect 132 102 135 105 
rect 132 105 135 108 
rect 132 108 135 111 
rect 132 111 135 114 
rect 132 114 135 117 
rect 132 117 135 120 
rect 132 120 135 123 
rect 132 123 135 126 
rect 132 126 135 129 
rect 132 129 135 132 
rect 132 132 135 135 
rect 132 135 135 138 
rect 132 138 135 141 
rect 132 141 135 144 
rect 132 144 135 147 
rect 132 147 135 150 
rect 132 150 135 153 
rect 132 153 135 156 
rect 132 156 135 159 
rect 132 159 135 162 
rect 132 162 135 165 
rect 132 165 135 168 
rect 132 168 135 171 
rect 132 171 135 174 
rect 132 174 135 177 
rect 132 177 135 180 
rect 132 180 135 183 
rect 132 183 135 186 
rect 132 186 135 189 
rect 132 189 135 192 
rect 132 192 135 195 
rect 132 195 135 198 
rect 132 198 135 201 
rect 132 201 135 204 
rect 132 204 135 207 
rect 132 207 135 210 
rect 132 210 135 213 
rect 132 213 135 216 
rect 132 216 135 219 
rect 132 219 135 222 
rect 132 222 135 225 
rect 132 225 135 228 
rect 132 228 135 231 
rect 132 231 135 234 
rect 132 234 135 237 
rect 132 237 135 240 
rect 132 240 135 243 
rect 132 243 135 246 
rect 132 246 135 249 
rect 132 249 135 252 
rect 132 252 135 255 
rect 132 255 135 258 
rect 132 258 135 261 
rect 132 261 135 264 
rect 132 264 135 267 
rect 132 267 135 270 
rect 132 270 135 273 
rect 132 273 135 276 
rect 132 276 135 279 
rect 132 279 135 282 
rect 132 282 135 285 
rect 132 285 135 288 
rect 132 288 135 291 
rect 132 291 135 294 
rect 132 294 135 297 
rect 132 297 135 300 
rect 132 300 135 303 
rect 132 303 135 306 
rect 132 306 135 309 
rect 132 309 135 312 
rect 132 312 135 315 
rect 132 315 135 318 
rect 132 318 135 321 
rect 132 321 135 324 
rect 132 324 135 327 
rect 132 327 135 330 
rect 132 330 135 333 
rect 132 333 135 336 
rect 132 336 135 339 
rect 132 339 135 342 
rect 132 342 135 345 
rect 132 345 135 348 
rect 132 348 135 351 
rect 132 351 135 354 
rect 132 354 135 357 
rect 132 357 135 360 
rect 132 360 135 363 
rect 132 363 135 366 
rect 132 366 135 369 
rect 132 369 135 372 
rect 132 372 135 375 
rect 132 375 135 378 
rect 132 378 135 381 
rect 132 381 135 384 
rect 132 384 135 387 
rect 132 387 135 390 
rect 132 390 135 393 
rect 132 393 135 396 
rect 132 396 135 399 
rect 132 399 135 402 
rect 132 402 135 405 
rect 132 405 135 408 
rect 132 408 135 411 
rect 132 411 135 414 
rect 132 414 135 417 
rect 132 417 135 420 
rect 132 420 135 423 
rect 132 423 135 426 
rect 132 426 135 429 
rect 132 429 135 432 
rect 132 432 135 435 
rect 132 435 135 438 
rect 132 438 135 441 
rect 132 441 135 444 
rect 132 444 135 447 
rect 132 447 135 450 
rect 132 450 135 453 
rect 132 453 135 456 
rect 132 456 135 459 
rect 132 459 135 462 
rect 132 462 135 465 
rect 132 465 135 468 
rect 132 468 135 471 
rect 132 471 135 474 
rect 132 474 135 477 
rect 132 477 135 480 
rect 132 480 135 483 
rect 132 483 135 486 
rect 132 486 135 489 
rect 132 489 135 492 
rect 132 492 135 495 
rect 132 495 135 498 
rect 132 498 135 501 
rect 132 501 135 504 
rect 132 504 135 507 
rect 132 507 135 510 
rect 135 0 138 3 
rect 135 3 138 6 
rect 135 6 138 9 
rect 135 9 138 12 
rect 135 12 138 15 
rect 135 15 138 18 
rect 135 18 138 21 
rect 135 21 138 24 
rect 135 24 138 27 
rect 135 27 138 30 
rect 135 30 138 33 
rect 135 33 138 36 
rect 135 36 138 39 
rect 135 39 138 42 
rect 135 42 138 45 
rect 135 45 138 48 
rect 135 48 138 51 
rect 135 51 138 54 
rect 135 54 138 57 
rect 135 57 138 60 
rect 135 60 138 63 
rect 135 63 138 66 
rect 135 66 138 69 
rect 135 69 138 72 
rect 135 72 138 75 
rect 135 75 138 78 
rect 135 78 138 81 
rect 135 81 138 84 
rect 135 84 138 87 
rect 135 87 138 90 
rect 135 90 138 93 
rect 135 93 138 96 
rect 135 96 138 99 
rect 135 99 138 102 
rect 135 102 138 105 
rect 135 105 138 108 
rect 135 108 138 111 
rect 135 111 138 114 
rect 135 114 138 117 
rect 135 117 138 120 
rect 135 120 138 123 
rect 135 123 138 126 
rect 135 126 138 129 
rect 135 129 138 132 
rect 135 132 138 135 
rect 135 135 138 138 
rect 135 138 138 141 
rect 135 141 138 144 
rect 135 144 138 147 
rect 135 147 138 150 
rect 135 150 138 153 
rect 135 153 138 156 
rect 135 156 138 159 
rect 135 159 138 162 
rect 135 162 138 165 
rect 135 165 138 168 
rect 135 168 138 171 
rect 135 171 138 174 
rect 135 174 138 177 
rect 135 177 138 180 
rect 135 180 138 183 
rect 135 183 138 186 
rect 135 186 138 189 
rect 135 189 138 192 
rect 135 192 138 195 
rect 135 195 138 198 
rect 135 198 138 201 
rect 135 201 138 204 
rect 135 204 138 207 
rect 135 207 138 210 
rect 135 210 138 213 
rect 135 213 138 216 
rect 135 216 138 219 
rect 135 219 138 222 
rect 135 222 138 225 
rect 135 225 138 228 
rect 135 228 138 231 
rect 135 231 138 234 
rect 135 234 138 237 
rect 135 237 138 240 
rect 135 240 138 243 
rect 135 243 138 246 
rect 135 246 138 249 
rect 135 249 138 252 
rect 135 252 138 255 
rect 135 255 138 258 
rect 135 258 138 261 
rect 135 261 138 264 
rect 135 264 138 267 
rect 135 267 138 270 
rect 135 270 138 273 
rect 135 273 138 276 
rect 135 276 138 279 
rect 135 279 138 282 
rect 135 282 138 285 
rect 135 285 138 288 
rect 135 288 138 291 
rect 135 291 138 294 
rect 135 294 138 297 
rect 135 297 138 300 
rect 135 300 138 303 
rect 135 303 138 306 
rect 135 306 138 309 
rect 135 309 138 312 
rect 135 312 138 315 
rect 135 315 138 318 
rect 135 318 138 321 
rect 135 321 138 324 
rect 135 324 138 327 
rect 135 327 138 330 
rect 135 330 138 333 
rect 135 333 138 336 
rect 135 336 138 339 
rect 135 339 138 342 
rect 135 342 138 345 
rect 135 345 138 348 
rect 135 348 138 351 
rect 135 351 138 354 
rect 135 354 138 357 
rect 135 357 138 360 
rect 135 360 138 363 
rect 135 363 138 366 
rect 135 366 138 369 
rect 135 369 138 372 
rect 135 372 138 375 
rect 135 375 138 378 
rect 135 378 138 381 
rect 135 381 138 384 
rect 135 384 138 387 
rect 135 387 138 390 
rect 135 390 138 393 
rect 135 393 138 396 
rect 135 396 138 399 
rect 135 399 138 402 
rect 135 402 138 405 
rect 135 405 138 408 
rect 135 408 138 411 
rect 135 411 138 414 
rect 135 414 138 417 
rect 135 417 138 420 
rect 135 420 138 423 
rect 135 423 138 426 
rect 135 426 138 429 
rect 135 429 138 432 
rect 135 432 138 435 
rect 135 435 138 438 
rect 135 438 138 441 
rect 135 441 138 444 
rect 135 444 138 447 
rect 135 447 138 450 
rect 135 450 138 453 
rect 135 453 138 456 
rect 135 456 138 459 
rect 135 459 138 462 
rect 135 462 138 465 
rect 135 465 138 468 
rect 135 468 138 471 
rect 135 471 138 474 
rect 135 474 138 477 
rect 135 477 138 480 
rect 135 480 138 483 
rect 135 483 138 486 
rect 135 486 138 489 
rect 135 489 138 492 
rect 135 492 138 495 
rect 135 495 138 498 
rect 135 498 138 501 
rect 135 501 138 504 
rect 135 504 138 507 
rect 135 507 138 510 
rect 138 0 141 3 
rect 138 3 141 6 
rect 138 6 141 9 
rect 138 9 141 12 
rect 138 12 141 15 
rect 138 15 141 18 
rect 138 18 141 21 
rect 138 21 141 24 
rect 138 24 141 27 
rect 138 27 141 30 
rect 138 30 141 33 
rect 138 33 141 36 
rect 138 36 141 39 
rect 138 39 141 42 
rect 138 42 141 45 
rect 138 45 141 48 
rect 138 48 141 51 
rect 138 51 141 54 
rect 138 54 141 57 
rect 138 57 141 60 
rect 138 60 141 63 
rect 138 63 141 66 
rect 138 66 141 69 
rect 138 69 141 72 
rect 138 72 141 75 
rect 138 75 141 78 
rect 138 78 141 81 
rect 138 81 141 84 
rect 138 84 141 87 
rect 138 87 141 90 
rect 138 90 141 93 
rect 138 93 141 96 
rect 138 96 141 99 
rect 138 99 141 102 
rect 138 102 141 105 
rect 138 105 141 108 
rect 138 108 141 111 
rect 138 111 141 114 
rect 138 114 141 117 
rect 138 117 141 120 
rect 138 120 141 123 
rect 138 123 141 126 
rect 138 126 141 129 
rect 138 129 141 132 
rect 138 132 141 135 
rect 138 135 141 138 
rect 138 138 141 141 
rect 138 141 141 144 
rect 138 144 141 147 
rect 138 147 141 150 
rect 138 150 141 153 
rect 138 153 141 156 
rect 138 156 141 159 
rect 138 159 141 162 
rect 138 162 141 165 
rect 138 165 141 168 
rect 138 168 141 171 
rect 138 171 141 174 
rect 138 174 141 177 
rect 138 177 141 180 
rect 138 180 141 183 
rect 138 183 141 186 
rect 138 186 141 189 
rect 138 189 141 192 
rect 138 192 141 195 
rect 138 195 141 198 
rect 138 198 141 201 
rect 138 201 141 204 
rect 138 204 141 207 
rect 138 207 141 210 
rect 138 210 141 213 
rect 138 213 141 216 
rect 138 216 141 219 
rect 138 219 141 222 
rect 138 222 141 225 
rect 138 225 141 228 
rect 138 228 141 231 
rect 138 231 141 234 
rect 138 234 141 237 
rect 138 237 141 240 
rect 138 240 141 243 
rect 138 243 141 246 
rect 138 246 141 249 
rect 138 249 141 252 
rect 138 252 141 255 
rect 138 255 141 258 
rect 138 258 141 261 
rect 138 261 141 264 
rect 138 264 141 267 
rect 138 267 141 270 
rect 138 270 141 273 
rect 138 273 141 276 
rect 138 276 141 279 
rect 138 279 141 282 
rect 138 282 141 285 
rect 138 285 141 288 
rect 138 288 141 291 
rect 138 291 141 294 
rect 138 294 141 297 
rect 138 297 141 300 
rect 138 300 141 303 
rect 138 303 141 306 
rect 138 306 141 309 
rect 138 309 141 312 
rect 138 312 141 315 
rect 138 315 141 318 
rect 138 318 141 321 
rect 138 321 141 324 
rect 138 324 141 327 
rect 138 327 141 330 
rect 138 330 141 333 
rect 138 333 141 336 
rect 138 336 141 339 
rect 138 339 141 342 
rect 138 342 141 345 
rect 138 345 141 348 
rect 138 348 141 351 
rect 138 351 141 354 
rect 138 354 141 357 
rect 138 357 141 360 
rect 138 360 141 363 
rect 138 363 141 366 
rect 138 366 141 369 
rect 138 369 141 372 
rect 138 372 141 375 
rect 138 375 141 378 
rect 138 378 141 381 
rect 138 381 141 384 
rect 138 384 141 387 
rect 138 387 141 390 
rect 138 390 141 393 
rect 138 393 141 396 
rect 138 396 141 399 
rect 138 399 141 402 
rect 138 402 141 405 
rect 138 405 141 408 
rect 138 408 141 411 
rect 138 411 141 414 
rect 138 414 141 417 
rect 138 417 141 420 
rect 138 420 141 423 
rect 138 423 141 426 
rect 138 426 141 429 
rect 138 429 141 432 
rect 138 432 141 435 
rect 138 435 141 438 
rect 138 438 141 441 
rect 138 441 141 444 
rect 138 444 141 447 
rect 138 447 141 450 
rect 138 450 141 453 
rect 138 453 141 456 
rect 138 456 141 459 
rect 138 459 141 462 
rect 138 462 141 465 
rect 138 465 141 468 
rect 138 468 141 471 
rect 138 471 141 474 
rect 138 474 141 477 
rect 138 477 141 480 
rect 138 480 141 483 
rect 138 483 141 486 
rect 138 486 141 489 
rect 138 489 141 492 
rect 138 492 141 495 
rect 138 495 141 498 
rect 138 498 141 501 
rect 138 501 141 504 
rect 138 504 141 507 
rect 138 507 141 510 
rect 141 0 144 3 
rect 141 3 144 6 
rect 141 6 144 9 
rect 141 9 144 12 
rect 141 12 144 15 
rect 141 15 144 18 
rect 141 18 144 21 
rect 141 21 144 24 
rect 141 24 144 27 
rect 141 27 144 30 
rect 141 30 144 33 
rect 141 33 144 36 
rect 141 36 144 39 
rect 141 39 144 42 
rect 141 42 144 45 
rect 141 45 144 48 
rect 141 48 144 51 
rect 141 51 144 54 
rect 141 54 144 57 
rect 141 57 144 60 
rect 141 60 144 63 
rect 141 63 144 66 
rect 141 66 144 69 
rect 141 69 144 72 
rect 141 72 144 75 
rect 141 75 144 78 
rect 141 78 144 81 
rect 141 84 144 87 
rect 141 87 144 90 
rect 141 90 144 93 
rect 141 93 144 96 
rect 141 96 144 99 
rect 141 99 144 102 
rect 141 102 144 105 
rect 141 105 144 108 
rect 141 108 144 111 
rect 141 111 144 114 
rect 141 114 144 117 
rect 141 117 144 120 
rect 141 120 144 123 
rect 141 123 144 126 
rect 141 126 144 129 
rect 141 129 144 132 
rect 141 132 144 135 
rect 141 135 144 138 
rect 141 138 144 141 
rect 141 141 144 144 
rect 141 144 144 147 
rect 141 147 144 150 
rect 141 150 144 153 
rect 141 153 144 156 
rect 141 156 144 159 
rect 141 159 144 162 
rect 141 162 144 165 
rect 141 165 144 168 
rect 141 168 144 171 
rect 141 171 144 174 
rect 141 174 144 177 
rect 141 177 144 180 
rect 141 180 144 183 
rect 141 183 144 186 
rect 141 186 144 189 
rect 141 189 144 192 
rect 141 192 144 195 
rect 141 195 144 198 
rect 141 198 144 201 
rect 141 201 144 204 
rect 141 204 144 207 
rect 141 207 144 210 
rect 141 210 144 213 
rect 141 213 144 216 
rect 141 216 144 219 
rect 141 219 144 222 
rect 141 222 144 225 
rect 141 228 144 231 
rect 141 231 144 234 
rect 141 237 144 240 
rect 141 240 144 243 
rect 141 243 144 246 
rect 141 246 144 249 
rect 141 249 144 252 
rect 141 252 144 255 
rect 141 255 144 258 
rect 141 258 144 261 
rect 141 261 144 264 
rect 141 264 144 267 
rect 141 267 144 270 
rect 141 270 144 273 
rect 141 273 144 276 
rect 141 276 144 279 
rect 141 279 144 282 
rect 141 282 144 285 
rect 141 285 144 288 
rect 141 288 144 291 
rect 141 291 144 294 
rect 141 294 144 297 
rect 141 297 144 300 
rect 141 300 144 303 
rect 141 303 144 306 
rect 141 306 144 309 
rect 141 309 144 312 
rect 141 312 144 315 
rect 141 315 144 318 
rect 141 318 144 321 
rect 141 324 144 327 
rect 141 327 144 330 
rect 141 333 144 336 
rect 141 336 144 339 
rect 141 339 144 342 
rect 141 342 144 345 
rect 141 345 144 348 
rect 141 348 144 351 
rect 141 351 144 354 
rect 141 354 144 357 
rect 141 357 144 360 
rect 141 360 144 363 
rect 141 363 144 366 
rect 141 366 144 369 
rect 141 369 144 372 
rect 141 372 144 375 
rect 141 375 144 378 
rect 141 378 144 381 
rect 141 381 144 384 
rect 141 384 144 387 
rect 141 387 144 390 
rect 141 390 144 393 
rect 141 393 144 396 
rect 141 396 144 399 
rect 141 399 144 402 
rect 141 402 144 405 
rect 141 405 144 408 
rect 141 408 144 411 
rect 141 411 144 414 
rect 141 414 144 417 
rect 141 420 144 423 
rect 141 423 144 426 
rect 141 429 144 432 
rect 141 432 144 435 
rect 141 435 144 438 
rect 141 438 144 441 
rect 141 441 144 444 
rect 141 444 144 447 
rect 141 447 144 450 
rect 141 450 144 453 
rect 141 453 144 456 
rect 141 456 144 459 
rect 141 459 144 462 
rect 141 462 144 465 
rect 141 465 144 468 
rect 141 468 144 471 
rect 141 471 144 474 
rect 141 474 144 477 
rect 141 477 144 480 
rect 141 480 144 483 
rect 141 483 144 486 
rect 141 486 144 489 
rect 141 489 144 492 
rect 141 492 144 495 
rect 141 495 144 498 
rect 141 498 144 501 
rect 141 501 144 504 
rect 141 504 144 507 
rect 141 507 144 510 
rect 144 0 147 3 
rect 144 3 147 6 
rect 144 6 147 9 
rect 144 9 147 12 
rect 144 12 147 15 
rect 144 15 147 18 
rect 144 18 147 21 
rect 144 21 147 24 
rect 144 24 147 27 
rect 144 27 147 30 
rect 144 30 147 33 
rect 144 33 147 36 
rect 144 36 147 39 
rect 144 39 147 42 
rect 144 42 147 45 
rect 144 45 147 48 
rect 144 48 147 51 
rect 144 51 147 54 
rect 144 54 147 57 
rect 144 57 147 60 
rect 144 60 147 63 
rect 144 63 147 66 
rect 144 66 147 69 
rect 144 69 147 72 
rect 144 72 147 75 
rect 144 75 147 78 
rect 144 78 147 81 
rect 144 81 147 84 
rect 144 84 147 87 
rect 144 87 147 90 
rect 144 90 147 93 
rect 144 93 147 96 
rect 144 96 147 99 
rect 144 99 147 102 
rect 144 102 147 105 
rect 144 105 147 108 
rect 144 108 147 111 
rect 144 111 147 114 
rect 144 114 147 117 
rect 144 117 147 120 
rect 144 120 147 123 
rect 144 123 147 126 
rect 144 126 147 129 
rect 144 129 147 132 
rect 144 132 147 135 
rect 144 135 147 138 
rect 144 138 147 141 
rect 144 141 147 144 
rect 144 144 147 147 
rect 144 147 147 150 
rect 144 150 147 153 
rect 144 153 147 156 
rect 144 156 147 159 
rect 144 159 147 162 
rect 144 162 147 165 
rect 144 165 147 168 
rect 144 168 147 171 
rect 144 171 147 174 
rect 144 174 147 177 
rect 144 177 147 180 
rect 144 180 147 183 
rect 144 183 147 186 
rect 144 186 147 189 
rect 144 189 147 192 
rect 144 192 147 195 
rect 144 195 147 198 
rect 144 198 147 201 
rect 144 201 147 204 
rect 144 204 147 207 
rect 144 207 147 210 
rect 144 210 147 213 
rect 144 213 147 216 
rect 144 216 147 219 
rect 144 219 147 222 
rect 144 222 147 225 
rect 144 225 147 228 
rect 144 228 147 231 
rect 144 231 147 234 
rect 144 234 147 237 
rect 144 237 147 240 
rect 144 240 147 243 
rect 144 243 147 246 
rect 144 246 147 249 
rect 144 249 147 252 
rect 144 252 147 255 
rect 144 255 147 258 
rect 144 258 147 261 
rect 144 261 147 264 
rect 144 264 147 267 
rect 144 267 147 270 
rect 144 270 147 273 
rect 144 273 147 276 
rect 144 276 147 279 
rect 144 279 147 282 
rect 144 282 147 285 
rect 144 285 147 288 
rect 144 288 147 291 
rect 144 291 147 294 
rect 144 294 147 297 
rect 144 297 147 300 
rect 144 300 147 303 
rect 144 303 147 306 
rect 144 306 147 309 
rect 144 309 147 312 
rect 144 312 147 315 
rect 144 315 147 318 
rect 144 318 147 321 
rect 144 321 147 324 
rect 144 324 147 327 
rect 144 327 147 330 
rect 144 330 147 333 
rect 144 333 147 336 
rect 144 336 147 339 
rect 144 339 147 342 
rect 144 342 147 345 
rect 144 345 147 348 
rect 144 348 147 351 
rect 144 351 147 354 
rect 144 354 147 357 
rect 144 357 147 360 
rect 144 360 147 363 
rect 144 363 147 366 
rect 144 366 147 369 
rect 144 369 147 372 
rect 144 372 147 375 
rect 144 375 147 378 
rect 144 378 147 381 
rect 144 381 147 384 
rect 144 384 147 387 
rect 144 387 147 390 
rect 144 390 147 393 
rect 144 393 147 396 
rect 144 396 147 399 
rect 144 399 147 402 
rect 144 402 147 405 
rect 144 405 147 408 
rect 144 408 147 411 
rect 144 411 147 414 
rect 144 414 147 417 
rect 144 417 147 420 
rect 144 420 147 423 
rect 144 423 147 426 
rect 144 426 147 429 
rect 144 429 147 432 
rect 144 432 147 435 
rect 144 435 147 438 
rect 144 438 147 441 
rect 144 441 147 444 
rect 144 444 147 447 
rect 144 447 147 450 
rect 144 450 147 453 
rect 144 453 147 456 
rect 144 456 147 459 
rect 144 459 147 462 
rect 144 462 147 465 
rect 144 465 147 468 
rect 144 468 147 471 
rect 144 471 147 474 
rect 144 474 147 477 
rect 144 477 147 480 
rect 144 480 147 483 
rect 144 483 147 486 
rect 144 486 147 489 
rect 144 489 147 492 
rect 144 492 147 495 
rect 144 495 147 498 
rect 144 498 147 501 
rect 144 501 147 504 
rect 144 504 147 507 
rect 144 507 147 510 
rect 147 0 150 3 
rect 147 3 150 6 
rect 147 6 150 9 
rect 147 9 150 12 
rect 147 12 150 15 
rect 147 15 150 18 
rect 147 18 150 21 
rect 147 21 150 24 
rect 147 24 150 27 
rect 147 27 150 30 
rect 147 30 150 33 
rect 147 33 150 36 
rect 147 36 150 39 
rect 147 39 150 42 
rect 147 42 150 45 
rect 147 45 150 48 
rect 147 48 150 51 
rect 147 51 150 54 
rect 147 54 150 57 
rect 147 57 150 60 
rect 147 60 150 63 
rect 147 63 150 66 
rect 147 66 150 69 
rect 147 69 150 72 
rect 147 72 150 75 
rect 147 75 150 78 
rect 147 78 150 81 
rect 147 81 150 84 
rect 147 84 150 87 
rect 147 87 150 90 
rect 147 90 150 93 
rect 147 93 150 96 
rect 147 96 150 99 
rect 147 99 150 102 
rect 147 102 150 105 
rect 147 105 150 108 
rect 147 108 150 111 
rect 147 111 150 114 
rect 147 114 150 117 
rect 147 117 150 120 
rect 147 120 150 123 
rect 147 123 150 126 
rect 147 126 150 129 
rect 147 129 150 132 
rect 147 132 150 135 
rect 147 135 150 138 
rect 147 138 150 141 
rect 147 141 150 144 
rect 147 144 150 147 
rect 147 147 150 150 
rect 147 150 150 153 
rect 147 153 150 156 
rect 147 156 150 159 
rect 147 159 150 162 
rect 147 162 150 165 
rect 147 165 150 168 
rect 147 168 150 171 
rect 147 171 150 174 
rect 147 174 150 177 
rect 147 177 150 180 
rect 147 180 150 183 
rect 147 183 150 186 
rect 147 186 150 189 
rect 147 189 150 192 
rect 147 192 150 195 
rect 147 195 150 198 
rect 147 198 150 201 
rect 147 201 150 204 
rect 147 204 150 207 
rect 147 207 150 210 
rect 147 210 150 213 
rect 147 213 150 216 
rect 147 216 150 219 
rect 147 219 150 222 
rect 147 222 150 225 
rect 147 225 150 228 
rect 147 228 150 231 
rect 147 231 150 234 
rect 147 234 150 237 
rect 147 237 150 240 
rect 147 240 150 243 
rect 147 243 150 246 
rect 147 246 150 249 
rect 147 249 150 252 
rect 147 252 150 255 
rect 147 255 150 258 
rect 147 258 150 261 
rect 147 261 150 264 
rect 147 264 150 267 
rect 147 267 150 270 
rect 147 270 150 273 
rect 147 273 150 276 
rect 147 276 150 279 
rect 147 279 150 282 
rect 147 282 150 285 
rect 147 285 150 288 
rect 147 288 150 291 
rect 147 291 150 294 
rect 147 294 150 297 
rect 147 297 150 300 
rect 147 300 150 303 
rect 147 303 150 306 
rect 147 306 150 309 
rect 147 309 150 312 
rect 147 312 150 315 
rect 147 315 150 318 
rect 147 318 150 321 
rect 147 321 150 324 
rect 147 324 150 327 
rect 147 327 150 330 
rect 147 330 150 333 
rect 147 333 150 336 
rect 147 336 150 339 
rect 147 339 150 342 
rect 147 342 150 345 
rect 147 345 150 348 
rect 147 348 150 351 
rect 147 351 150 354 
rect 147 354 150 357 
rect 147 357 150 360 
rect 147 360 150 363 
rect 147 363 150 366 
rect 147 366 150 369 
rect 147 369 150 372 
rect 147 372 150 375 
rect 147 375 150 378 
rect 147 378 150 381 
rect 147 381 150 384 
rect 147 384 150 387 
rect 147 387 150 390 
rect 147 390 150 393 
rect 147 393 150 396 
rect 147 396 150 399 
rect 147 399 150 402 
rect 147 402 150 405 
rect 147 405 150 408 
rect 147 408 150 411 
rect 147 411 150 414 
rect 147 414 150 417 
rect 147 417 150 420 
rect 147 420 150 423 
rect 147 423 150 426 
rect 147 426 150 429 
rect 147 429 150 432 
rect 147 432 150 435 
rect 147 435 150 438 
rect 147 438 150 441 
rect 147 441 150 444 
rect 147 444 150 447 
rect 147 447 150 450 
rect 147 450 150 453 
rect 147 453 150 456 
rect 147 456 150 459 
rect 147 459 150 462 
rect 147 462 150 465 
rect 147 465 150 468 
rect 147 468 150 471 
rect 147 471 150 474 
rect 147 474 150 477 
rect 147 477 150 480 
rect 147 480 150 483 
rect 147 483 150 486 
rect 147 486 150 489 
rect 147 489 150 492 
rect 147 492 150 495 
rect 147 495 150 498 
rect 147 498 150 501 
rect 147 501 150 504 
rect 147 504 150 507 
rect 147 507 150 510 
rect 150 0 153 3 
rect 150 3 153 6 
rect 150 6 153 9 
rect 150 9 153 12 
rect 150 12 153 15 
rect 150 15 153 18 
rect 150 18 153 21 
rect 150 21 153 24 
rect 150 24 153 27 
rect 150 27 153 30 
rect 150 30 153 33 
rect 150 33 153 36 
rect 150 36 153 39 
rect 150 39 153 42 
rect 150 42 153 45 
rect 150 45 153 48 
rect 150 48 153 51 
rect 150 51 153 54 
rect 150 54 153 57 
rect 150 57 153 60 
rect 150 60 153 63 
rect 150 63 153 66 
rect 150 66 153 69 
rect 150 69 153 72 
rect 150 72 153 75 
rect 150 75 153 78 
rect 150 78 153 81 
rect 150 81 153 84 
rect 150 84 153 87 
rect 150 87 153 90 
rect 150 90 153 93 
rect 150 93 153 96 
rect 150 96 153 99 
rect 150 99 153 102 
rect 150 102 153 105 
rect 150 105 153 108 
rect 150 108 153 111 
rect 150 111 153 114 
rect 150 114 153 117 
rect 150 117 153 120 
rect 150 120 153 123 
rect 150 123 153 126 
rect 150 126 153 129 
rect 150 129 153 132 
rect 150 132 153 135 
rect 150 135 153 138 
rect 150 138 153 141 
rect 150 141 153 144 
rect 150 144 153 147 
rect 150 147 153 150 
rect 150 150 153 153 
rect 150 153 153 156 
rect 150 156 153 159 
rect 150 159 153 162 
rect 150 162 153 165 
rect 150 165 153 168 
rect 150 168 153 171 
rect 150 171 153 174 
rect 150 174 153 177 
rect 150 177 153 180 
rect 150 180 153 183 
rect 150 183 153 186 
rect 150 186 153 189 
rect 150 189 153 192 
rect 150 192 153 195 
rect 150 195 153 198 
rect 150 198 153 201 
rect 150 201 153 204 
rect 150 204 153 207 
rect 150 207 153 210 
rect 150 210 153 213 
rect 150 213 153 216 
rect 150 216 153 219 
rect 150 219 153 222 
rect 150 222 153 225 
rect 150 225 153 228 
rect 150 228 153 231 
rect 150 231 153 234 
rect 150 234 153 237 
rect 150 237 153 240 
rect 150 240 153 243 
rect 150 243 153 246 
rect 150 246 153 249 
rect 150 249 153 252 
rect 150 252 153 255 
rect 150 255 153 258 
rect 150 258 153 261 
rect 150 261 153 264 
rect 150 264 153 267 
rect 150 267 153 270 
rect 150 270 153 273 
rect 150 273 153 276 
rect 150 276 153 279 
rect 150 279 153 282 
rect 150 282 153 285 
rect 150 285 153 288 
rect 150 288 153 291 
rect 150 291 153 294 
rect 150 294 153 297 
rect 150 297 153 300 
rect 150 300 153 303 
rect 150 303 153 306 
rect 150 306 153 309 
rect 150 309 153 312 
rect 150 312 153 315 
rect 150 315 153 318 
rect 150 318 153 321 
rect 150 321 153 324 
rect 150 324 153 327 
rect 150 327 153 330 
rect 150 330 153 333 
rect 150 333 153 336 
rect 150 336 153 339 
rect 150 339 153 342 
rect 150 342 153 345 
rect 150 345 153 348 
rect 150 348 153 351 
rect 150 351 153 354 
rect 150 354 153 357 
rect 150 357 153 360 
rect 150 360 153 363 
rect 150 363 153 366 
rect 150 366 153 369 
rect 150 369 153 372 
rect 150 372 153 375 
rect 150 375 153 378 
rect 150 378 153 381 
rect 150 381 153 384 
rect 150 384 153 387 
rect 150 387 153 390 
rect 150 390 153 393 
rect 150 393 153 396 
rect 150 396 153 399 
rect 150 399 153 402 
rect 150 402 153 405 
rect 150 405 153 408 
rect 150 408 153 411 
rect 150 411 153 414 
rect 150 414 153 417 
rect 150 417 153 420 
rect 150 420 153 423 
rect 150 423 153 426 
rect 150 426 153 429 
rect 150 429 153 432 
rect 150 432 153 435 
rect 150 435 153 438 
rect 150 438 153 441 
rect 150 441 153 444 
rect 150 444 153 447 
rect 150 447 153 450 
rect 150 450 153 453 
rect 150 453 153 456 
rect 150 456 153 459 
rect 150 459 153 462 
rect 150 462 153 465 
rect 150 465 153 468 
rect 150 468 153 471 
rect 150 471 153 474 
rect 150 474 153 477 
rect 150 477 153 480 
rect 150 480 153 483 
rect 150 483 153 486 
rect 150 486 153 489 
rect 150 489 153 492 
rect 150 492 153 495 
rect 150 495 153 498 
rect 150 498 153 501 
rect 150 501 153 504 
rect 150 504 153 507 
rect 150 507 153 510 
rect 153 0 156 3 
rect 153 3 156 6 
rect 153 6 156 9 
rect 153 9 156 12 
rect 153 12 156 15 
rect 153 15 156 18 
rect 153 18 156 21 
rect 153 21 156 24 
rect 153 24 156 27 
rect 153 27 156 30 
rect 153 30 156 33 
rect 153 33 156 36 
rect 153 36 156 39 
rect 153 39 156 42 
rect 153 42 156 45 
rect 153 45 156 48 
rect 153 48 156 51 
rect 153 51 156 54 
rect 153 54 156 57 
rect 153 57 156 60 
rect 153 60 156 63 
rect 153 63 156 66 
rect 153 66 156 69 
rect 153 69 156 72 
rect 153 72 156 75 
rect 153 75 156 78 
rect 153 78 156 81 
rect 153 81 156 84 
rect 153 84 156 87 
rect 153 87 156 90 
rect 153 90 156 93 
rect 153 93 156 96 
rect 153 96 156 99 
rect 153 99 156 102 
rect 153 102 156 105 
rect 153 105 156 108 
rect 153 108 156 111 
rect 153 111 156 114 
rect 153 114 156 117 
rect 153 117 156 120 
rect 153 120 156 123 
rect 153 123 156 126 
rect 153 126 156 129 
rect 153 129 156 132 
rect 153 132 156 135 
rect 153 135 156 138 
rect 153 138 156 141 
rect 153 141 156 144 
rect 153 144 156 147 
rect 153 147 156 150 
rect 153 150 156 153 
rect 153 153 156 156 
rect 153 156 156 159 
rect 153 159 156 162 
rect 153 162 156 165 
rect 153 165 156 168 
rect 153 168 156 171 
rect 153 171 156 174 
rect 153 174 156 177 
rect 153 177 156 180 
rect 153 180 156 183 
rect 153 183 156 186 
rect 153 186 156 189 
rect 153 189 156 192 
rect 153 192 156 195 
rect 153 195 156 198 
rect 153 198 156 201 
rect 153 201 156 204 
rect 153 204 156 207 
rect 153 207 156 210 
rect 153 210 156 213 
rect 153 213 156 216 
rect 153 216 156 219 
rect 153 219 156 222 
rect 153 222 156 225 
rect 153 225 156 228 
rect 153 228 156 231 
rect 153 231 156 234 
rect 153 234 156 237 
rect 153 237 156 240 
rect 153 240 156 243 
rect 153 243 156 246 
rect 153 246 156 249 
rect 153 249 156 252 
rect 153 252 156 255 
rect 153 255 156 258 
rect 153 258 156 261 
rect 153 261 156 264 
rect 153 264 156 267 
rect 153 267 156 270 
rect 153 270 156 273 
rect 153 273 156 276 
rect 153 276 156 279 
rect 153 279 156 282 
rect 153 282 156 285 
rect 153 285 156 288 
rect 153 288 156 291 
rect 153 291 156 294 
rect 153 294 156 297 
rect 153 297 156 300 
rect 153 300 156 303 
rect 153 303 156 306 
rect 153 306 156 309 
rect 153 309 156 312 
rect 153 312 156 315 
rect 153 315 156 318 
rect 153 318 156 321 
rect 153 321 156 324 
rect 153 324 156 327 
rect 153 327 156 330 
rect 153 330 156 333 
rect 153 333 156 336 
rect 153 336 156 339 
rect 153 339 156 342 
rect 153 342 156 345 
rect 153 345 156 348 
rect 153 348 156 351 
rect 153 351 156 354 
rect 153 354 156 357 
rect 153 357 156 360 
rect 153 360 156 363 
rect 153 363 156 366 
rect 153 366 156 369 
rect 153 369 156 372 
rect 153 372 156 375 
rect 153 375 156 378 
rect 153 378 156 381 
rect 153 381 156 384 
rect 153 384 156 387 
rect 153 387 156 390 
rect 153 390 156 393 
rect 153 393 156 396 
rect 153 396 156 399 
rect 153 399 156 402 
rect 153 402 156 405 
rect 153 405 156 408 
rect 153 408 156 411 
rect 153 411 156 414 
rect 153 414 156 417 
rect 153 417 156 420 
rect 153 420 156 423 
rect 153 423 156 426 
rect 153 426 156 429 
rect 153 429 156 432 
rect 153 432 156 435 
rect 153 435 156 438 
rect 153 438 156 441 
rect 153 441 156 444 
rect 153 444 156 447 
rect 153 447 156 450 
rect 153 450 156 453 
rect 153 453 156 456 
rect 153 456 156 459 
rect 153 459 156 462 
rect 153 462 156 465 
rect 153 465 156 468 
rect 153 468 156 471 
rect 153 471 156 474 
rect 153 474 156 477 
rect 153 477 156 480 
rect 153 480 156 483 
rect 153 483 156 486 
rect 153 486 156 489 
rect 153 489 156 492 
rect 153 492 156 495 
rect 153 495 156 498 
rect 153 498 156 501 
rect 153 501 156 504 
rect 153 504 156 507 
rect 153 507 156 510 
rect 156 0 159 3 
rect 156 3 159 6 
rect 156 6 159 9 
rect 156 9 159 12 
rect 156 12 159 15 
rect 156 15 159 18 
rect 156 18 159 21 
rect 156 21 159 24 
rect 156 24 159 27 
rect 156 27 159 30 
rect 156 30 159 33 
rect 156 33 159 36 
rect 156 36 159 39 
rect 156 39 159 42 
rect 156 42 159 45 
rect 156 45 159 48 
rect 156 48 159 51 
rect 156 51 159 54 
rect 156 54 159 57 
rect 156 57 159 60 
rect 156 60 159 63 
rect 156 63 159 66 
rect 156 66 159 69 
rect 156 69 159 72 
rect 156 72 159 75 
rect 156 75 159 78 
rect 156 78 159 81 
rect 156 81 159 84 
rect 156 84 159 87 
rect 156 87 159 90 
rect 156 90 159 93 
rect 156 93 159 96 
rect 156 96 159 99 
rect 156 99 159 102 
rect 156 102 159 105 
rect 156 105 159 108 
rect 156 108 159 111 
rect 156 111 159 114 
rect 156 114 159 117 
rect 156 117 159 120 
rect 156 120 159 123 
rect 156 123 159 126 
rect 156 126 159 129 
rect 156 129 159 132 
rect 156 132 159 135 
rect 156 135 159 138 
rect 156 138 159 141 
rect 156 141 159 144 
rect 156 144 159 147 
rect 156 147 159 150 
rect 156 150 159 153 
rect 156 153 159 156 
rect 156 156 159 159 
rect 156 159 159 162 
rect 156 162 159 165 
rect 156 165 159 168 
rect 156 168 159 171 
rect 156 171 159 174 
rect 156 174 159 177 
rect 156 177 159 180 
rect 156 180 159 183 
rect 156 183 159 186 
rect 156 186 159 189 
rect 156 189 159 192 
rect 156 192 159 195 
rect 156 195 159 198 
rect 156 198 159 201 
rect 156 201 159 204 
rect 156 204 159 207 
rect 156 207 159 210 
rect 156 210 159 213 
rect 156 213 159 216 
rect 156 216 159 219 
rect 156 219 159 222 
rect 156 222 159 225 
rect 156 225 159 228 
rect 156 228 159 231 
rect 156 231 159 234 
rect 156 234 159 237 
rect 156 237 159 240 
rect 156 240 159 243 
rect 156 243 159 246 
rect 156 246 159 249 
rect 156 249 159 252 
rect 156 252 159 255 
rect 156 255 159 258 
rect 156 258 159 261 
rect 156 261 159 264 
rect 156 264 159 267 
rect 156 267 159 270 
rect 156 270 159 273 
rect 156 273 159 276 
rect 156 276 159 279 
rect 156 279 159 282 
rect 156 282 159 285 
rect 156 285 159 288 
rect 156 288 159 291 
rect 156 291 159 294 
rect 156 294 159 297 
rect 156 297 159 300 
rect 156 300 159 303 
rect 156 303 159 306 
rect 156 306 159 309 
rect 156 309 159 312 
rect 156 312 159 315 
rect 156 315 159 318 
rect 156 318 159 321 
rect 156 321 159 324 
rect 156 324 159 327 
rect 156 327 159 330 
rect 156 330 159 333 
rect 156 333 159 336 
rect 156 336 159 339 
rect 156 339 159 342 
rect 156 342 159 345 
rect 156 345 159 348 
rect 156 348 159 351 
rect 156 351 159 354 
rect 156 354 159 357 
rect 156 357 159 360 
rect 156 360 159 363 
rect 156 363 159 366 
rect 156 366 159 369 
rect 156 369 159 372 
rect 156 372 159 375 
rect 156 375 159 378 
rect 156 378 159 381 
rect 156 381 159 384 
rect 156 384 159 387 
rect 156 387 159 390 
rect 156 390 159 393 
rect 156 393 159 396 
rect 156 396 159 399 
rect 156 399 159 402 
rect 156 402 159 405 
rect 156 405 159 408 
rect 156 408 159 411 
rect 156 411 159 414 
rect 156 414 159 417 
rect 156 417 159 420 
rect 156 420 159 423 
rect 156 423 159 426 
rect 156 426 159 429 
rect 156 429 159 432 
rect 156 432 159 435 
rect 156 435 159 438 
rect 156 438 159 441 
rect 156 441 159 444 
rect 156 444 159 447 
rect 156 447 159 450 
rect 156 450 159 453 
rect 156 453 159 456 
rect 156 456 159 459 
rect 156 459 159 462 
rect 156 462 159 465 
rect 156 465 159 468 
rect 156 468 159 471 
rect 156 471 159 474 
rect 156 474 159 477 
rect 156 477 159 480 
rect 156 480 159 483 
rect 156 483 159 486 
rect 156 486 159 489 
rect 156 489 159 492 
rect 156 492 159 495 
rect 156 495 159 498 
rect 156 498 159 501 
rect 156 501 159 504 
rect 156 504 159 507 
rect 156 507 159 510 
rect 159 0 162 3 
rect 159 3 162 6 
rect 159 6 162 9 
rect 159 9 162 12 
rect 159 12 162 15 
rect 159 15 162 18 
rect 159 18 162 21 
rect 159 21 162 24 
rect 159 24 162 27 
rect 159 27 162 30 
rect 159 30 162 33 
rect 159 33 162 36 
rect 159 36 162 39 
rect 159 39 162 42 
rect 159 42 162 45 
rect 159 45 162 48 
rect 159 48 162 51 
rect 159 51 162 54 
rect 159 54 162 57 
rect 159 57 162 60 
rect 159 60 162 63 
rect 159 63 162 66 
rect 159 66 162 69 
rect 159 69 162 72 
rect 159 72 162 75 
rect 159 75 162 78 
rect 159 78 162 81 
rect 159 81 162 84 
rect 159 84 162 87 
rect 159 87 162 90 
rect 159 90 162 93 
rect 159 93 162 96 
rect 159 96 162 99 
rect 159 99 162 102 
rect 159 102 162 105 
rect 159 105 162 108 
rect 159 108 162 111 
rect 159 111 162 114 
rect 159 114 162 117 
rect 159 117 162 120 
rect 159 120 162 123 
rect 159 123 162 126 
rect 159 126 162 129 
rect 159 129 162 132 
rect 159 132 162 135 
rect 159 135 162 138 
rect 159 138 162 141 
rect 159 141 162 144 
rect 159 144 162 147 
rect 159 147 162 150 
rect 159 150 162 153 
rect 159 153 162 156 
rect 159 156 162 159 
rect 159 159 162 162 
rect 159 162 162 165 
rect 159 165 162 168 
rect 159 168 162 171 
rect 159 171 162 174 
rect 159 174 162 177 
rect 159 177 162 180 
rect 159 180 162 183 
rect 159 183 162 186 
rect 159 186 162 189 
rect 159 189 162 192 
rect 159 192 162 195 
rect 159 195 162 198 
rect 159 198 162 201 
rect 159 201 162 204 
rect 159 204 162 207 
rect 159 207 162 210 
rect 159 210 162 213 
rect 159 213 162 216 
rect 159 216 162 219 
rect 159 219 162 222 
rect 159 222 162 225 
rect 159 225 162 228 
rect 159 228 162 231 
rect 159 231 162 234 
rect 159 234 162 237 
rect 159 237 162 240 
rect 159 240 162 243 
rect 159 243 162 246 
rect 159 246 162 249 
rect 159 249 162 252 
rect 159 252 162 255 
rect 159 255 162 258 
rect 159 258 162 261 
rect 159 261 162 264 
rect 159 264 162 267 
rect 159 267 162 270 
rect 159 270 162 273 
rect 159 273 162 276 
rect 159 276 162 279 
rect 159 279 162 282 
rect 159 282 162 285 
rect 159 285 162 288 
rect 159 288 162 291 
rect 159 291 162 294 
rect 159 294 162 297 
rect 159 297 162 300 
rect 159 300 162 303 
rect 159 303 162 306 
rect 159 306 162 309 
rect 159 309 162 312 
rect 159 312 162 315 
rect 159 315 162 318 
rect 159 318 162 321 
rect 159 321 162 324 
rect 159 324 162 327 
rect 159 327 162 330 
rect 159 330 162 333 
rect 159 333 162 336 
rect 159 336 162 339 
rect 159 339 162 342 
rect 159 342 162 345 
rect 159 345 162 348 
rect 159 348 162 351 
rect 159 351 162 354 
rect 159 354 162 357 
rect 159 357 162 360 
rect 159 360 162 363 
rect 159 363 162 366 
rect 159 366 162 369 
rect 159 369 162 372 
rect 159 372 162 375 
rect 159 375 162 378 
rect 159 378 162 381 
rect 159 381 162 384 
rect 159 384 162 387 
rect 159 387 162 390 
rect 159 390 162 393 
rect 159 393 162 396 
rect 159 396 162 399 
rect 159 399 162 402 
rect 159 402 162 405 
rect 159 405 162 408 
rect 159 408 162 411 
rect 159 411 162 414 
rect 159 414 162 417 
rect 159 417 162 420 
rect 159 420 162 423 
rect 159 423 162 426 
rect 159 426 162 429 
rect 159 429 162 432 
rect 159 432 162 435 
rect 159 435 162 438 
rect 159 438 162 441 
rect 159 441 162 444 
rect 159 444 162 447 
rect 159 447 162 450 
rect 159 450 162 453 
rect 159 453 162 456 
rect 159 456 162 459 
rect 159 459 162 462 
rect 159 462 162 465 
rect 159 465 162 468 
rect 159 468 162 471 
rect 159 471 162 474 
rect 159 474 162 477 
rect 159 477 162 480 
rect 159 480 162 483 
rect 159 483 162 486 
rect 159 486 162 489 
rect 159 489 162 492 
rect 159 492 162 495 
rect 159 495 162 498 
rect 159 498 162 501 
rect 159 501 162 504 
rect 159 504 162 507 
rect 159 507 162 510 
rect 162 0 165 3 
rect 162 3 165 6 
rect 162 6 165 9 
rect 162 9 165 12 
rect 162 12 165 15 
rect 162 15 165 18 
rect 162 18 165 21 
rect 162 21 165 24 
rect 162 24 165 27 
rect 162 27 165 30 
rect 162 30 165 33 
rect 162 33 165 36 
rect 162 36 165 39 
rect 162 39 165 42 
rect 162 42 165 45 
rect 162 45 165 48 
rect 162 48 165 51 
rect 162 51 165 54 
rect 162 54 165 57 
rect 162 57 165 60 
rect 162 60 165 63 
rect 162 63 165 66 
rect 162 66 165 69 
rect 162 69 165 72 
rect 162 72 165 75 
rect 162 75 165 78 
rect 162 78 165 81 
rect 162 81 165 84 
rect 162 84 165 87 
rect 162 87 165 90 
rect 162 90 165 93 
rect 162 93 165 96 
rect 162 96 165 99 
rect 162 99 165 102 
rect 162 102 165 105 
rect 162 105 165 108 
rect 162 108 165 111 
rect 162 111 165 114 
rect 162 114 165 117 
rect 162 117 165 120 
rect 162 120 165 123 
rect 162 123 165 126 
rect 162 126 165 129 
rect 162 129 165 132 
rect 162 132 165 135 
rect 162 135 165 138 
rect 162 138 165 141 
rect 162 141 165 144 
rect 162 144 165 147 
rect 162 147 165 150 
rect 162 150 165 153 
rect 162 153 165 156 
rect 162 156 165 159 
rect 162 159 165 162 
rect 162 162 165 165 
rect 162 165 165 168 
rect 162 168 165 171 
rect 162 171 165 174 
rect 162 174 165 177 
rect 162 177 165 180 
rect 162 180 165 183 
rect 162 183 165 186 
rect 162 186 165 189 
rect 162 189 165 192 
rect 162 192 165 195 
rect 162 195 165 198 
rect 162 198 165 201 
rect 162 201 165 204 
rect 162 204 165 207 
rect 162 207 165 210 
rect 162 210 165 213 
rect 162 213 165 216 
rect 162 216 165 219 
rect 162 219 165 222 
rect 162 222 165 225 
rect 162 225 165 228 
rect 162 228 165 231 
rect 162 231 165 234 
rect 162 234 165 237 
rect 162 237 165 240 
rect 162 240 165 243 
rect 162 243 165 246 
rect 162 246 165 249 
rect 162 249 165 252 
rect 162 252 165 255 
rect 162 255 165 258 
rect 162 258 165 261 
rect 162 261 165 264 
rect 162 264 165 267 
rect 162 267 165 270 
rect 162 270 165 273 
rect 162 273 165 276 
rect 162 276 165 279 
rect 162 279 165 282 
rect 162 282 165 285 
rect 162 285 165 288 
rect 162 288 165 291 
rect 162 291 165 294 
rect 162 294 165 297 
rect 162 297 165 300 
rect 162 300 165 303 
rect 162 303 165 306 
rect 162 306 165 309 
rect 162 309 165 312 
rect 162 312 165 315 
rect 162 315 165 318 
rect 162 318 165 321 
rect 162 321 165 324 
rect 162 324 165 327 
rect 162 327 165 330 
rect 162 330 165 333 
rect 162 333 165 336 
rect 162 336 165 339 
rect 162 339 165 342 
rect 162 342 165 345 
rect 162 345 165 348 
rect 162 348 165 351 
rect 162 351 165 354 
rect 162 354 165 357 
rect 162 357 165 360 
rect 162 360 165 363 
rect 162 363 165 366 
rect 162 366 165 369 
rect 162 369 165 372 
rect 162 372 165 375 
rect 162 375 165 378 
rect 162 378 165 381 
rect 162 381 165 384 
rect 162 384 165 387 
rect 162 387 165 390 
rect 162 390 165 393 
rect 162 393 165 396 
rect 162 396 165 399 
rect 162 399 165 402 
rect 162 402 165 405 
rect 162 405 165 408 
rect 162 408 165 411 
rect 162 411 165 414 
rect 162 414 165 417 
rect 162 417 165 420 
rect 162 420 165 423 
rect 162 423 165 426 
rect 162 426 165 429 
rect 162 429 165 432 
rect 162 432 165 435 
rect 162 435 165 438 
rect 162 438 165 441 
rect 162 441 165 444 
rect 162 444 165 447 
rect 162 447 165 450 
rect 162 450 165 453 
rect 162 453 165 456 
rect 162 456 165 459 
rect 162 459 165 462 
rect 162 462 165 465 
rect 162 465 165 468 
rect 162 468 165 471 
rect 162 471 165 474 
rect 162 474 165 477 
rect 162 477 165 480 
rect 162 480 165 483 
rect 162 483 165 486 
rect 162 486 165 489 
rect 162 489 165 492 
rect 162 492 165 495 
rect 162 495 165 498 
rect 162 498 165 501 
rect 162 501 165 504 
rect 162 504 165 507 
rect 162 507 165 510 
rect 165 0 168 3 
rect 165 3 168 6 
rect 165 6 168 9 
rect 165 9 168 12 
rect 165 12 168 15 
rect 165 15 168 18 
rect 165 18 168 21 
rect 165 21 168 24 
rect 165 24 168 27 
rect 165 27 168 30 
rect 165 30 168 33 
rect 165 33 168 36 
rect 165 36 168 39 
rect 165 39 168 42 
rect 165 42 168 45 
rect 165 45 168 48 
rect 165 48 168 51 
rect 165 51 168 54 
rect 165 54 168 57 
rect 165 57 168 60 
rect 165 60 168 63 
rect 165 63 168 66 
rect 165 66 168 69 
rect 165 69 168 72 
rect 165 72 168 75 
rect 165 75 168 78 
rect 165 78 168 81 
rect 165 81 168 84 
rect 165 84 168 87 
rect 165 87 168 90 
rect 165 90 168 93 
rect 165 93 168 96 
rect 165 96 168 99 
rect 165 99 168 102 
rect 165 102 168 105 
rect 165 105 168 108 
rect 165 108 168 111 
rect 165 111 168 114 
rect 165 114 168 117 
rect 165 117 168 120 
rect 165 120 168 123 
rect 165 123 168 126 
rect 165 126 168 129 
rect 165 129 168 132 
rect 165 132 168 135 
rect 165 135 168 138 
rect 165 138 168 141 
rect 165 141 168 144 
rect 165 144 168 147 
rect 165 147 168 150 
rect 165 150 168 153 
rect 165 153 168 156 
rect 165 156 168 159 
rect 165 159 168 162 
rect 165 162 168 165 
rect 165 165 168 168 
rect 165 168 168 171 
rect 165 171 168 174 
rect 165 174 168 177 
rect 165 177 168 180 
rect 165 180 168 183 
rect 165 183 168 186 
rect 165 186 168 189 
rect 165 189 168 192 
rect 165 192 168 195 
rect 165 195 168 198 
rect 165 198 168 201 
rect 165 201 168 204 
rect 165 204 168 207 
rect 165 207 168 210 
rect 165 210 168 213 
rect 165 213 168 216 
rect 165 216 168 219 
rect 165 219 168 222 
rect 165 222 168 225 
rect 165 225 168 228 
rect 165 228 168 231 
rect 165 231 168 234 
rect 165 234 168 237 
rect 165 237 168 240 
rect 165 240 168 243 
rect 165 243 168 246 
rect 165 246 168 249 
rect 165 249 168 252 
rect 165 252 168 255 
rect 165 255 168 258 
rect 165 258 168 261 
rect 165 261 168 264 
rect 165 264 168 267 
rect 165 267 168 270 
rect 165 270 168 273 
rect 165 273 168 276 
rect 165 276 168 279 
rect 165 279 168 282 
rect 165 282 168 285 
rect 165 285 168 288 
rect 165 288 168 291 
rect 165 291 168 294 
rect 165 294 168 297 
rect 165 297 168 300 
rect 165 300 168 303 
rect 165 303 168 306 
rect 165 306 168 309 
rect 165 309 168 312 
rect 165 312 168 315 
rect 165 315 168 318 
rect 165 318 168 321 
rect 165 321 168 324 
rect 165 324 168 327 
rect 165 327 168 330 
rect 165 330 168 333 
rect 165 333 168 336 
rect 165 336 168 339 
rect 165 339 168 342 
rect 165 342 168 345 
rect 165 345 168 348 
rect 165 348 168 351 
rect 165 351 168 354 
rect 165 354 168 357 
rect 165 357 168 360 
rect 165 360 168 363 
rect 165 363 168 366 
rect 165 366 168 369 
rect 165 369 168 372 
rect 165 372 168 375 
rect 165 375 168 378 
rect 165 378 168 381 
rect 165 381 168 384 
rect 165 384 168 387 
rect 165 387 168 390 
rect 165 390 168 393 
rect 165 393 168 396 
rect 165 396 168 399 
rect 165 399 168 402 
rect 165 402 168 405 
rect 165 405 168 408 
rect 165 408 168 411 
rect 165 411 168 414 
rect 165 414 168 417 
rect 165 417 168 420 
rect 165 420 168 423 
rect 165 423 168 426 
rect 165 426 168 429 
rect 165 429 168 432 
rect 165 432 168 435 
rect 165 435 168 438 
rect 165 438 168 441 
rect 165 441 168 444 
rect 165 444 168 447 
rect 165 447 168 450 
rect 165 450 168 453 
rect 165 453 168 456 
rect 165 456 168 459 
rect 165 459 168 462 
rect 165 462 168 465 
rect 165 465 168 468 
rect 165 468 168 471 
rect 165 471 168 474 
rect 165 474 168 477 
rect 165 477 168 480 
rect 165 480 168 483 
rect 165 483 168 486 
rect 165 486 168 489 
rect 165 489 168 492 
rect 165 492 168 495 
rect 165 495 168 498 
rect 165 498 168 501 
rect 165 501 168 504 
rect 165 504 168 507 
rect 165 507 168 510 
rect 168 0 171 3 
rect 168 3 171 6 
rect 168 6 171 9 
rect 168 9 171 12 
rect 168 12 171 15 
rect 168 15 171 18 
rect 168 18 171 21 
rect 168 21 171 24 
rect 168 24 171 27 
rect 168 27 171 30 
rect 168 30 171 33 
rect 168 33 171 36 
rect 168 36 171 39 
rect 168 39 171 42 
rect 168 42 171 45 
rect 168 45 171 48 
rect 168 48 171 51 
rect 168 51 171 54 
rect 168 54 171 57 
rect 168 57 171 60 
rect 168 60 171 63 
rect 168 63 171 66 
rect 168 66 171 69 
rect 168 69 171 72 
rect 168 72 171 75 
rect 168 75 171 78 
rect 168 78 171 81 
rect 168 81 171 84 
rect 168 84 171 87 
rect 168 87 171 90 
rect 168 90 171 93 
rect 168 93 171 96 
rect 168 96 171 99 
rect 168 99 171 102 
rect 168 102 171 105 
rect 168 105 171 108 
rect 168 108 171 111 
rect 168 111 171 114 
rect 168 114 171 117 
rect 168 117 171 120 
rect 168 120 171 123 
rect 168 123 171 126 
rect 168 126 171 129 
rect 168 129 171 132 
rect 168 132 171 135 
rect 168 135 171 138 
rect 168 138 171 141 
rect 168 141 171 144 
rect 168 144 171 147 
rect 168 147 171 150 
rect 168 150 171 153 
rect 168 153 171 156 
rect 168 156 171 159 
rect 168 159 171 162 
rect 168 162 171 165 
rect 168 165 171 168 
rect 168 168 171 171 
rect 168 171 171 174 
rect 168 174 171 177 
rect 168 177 171 180 
rect 168 180 171 183 
rect 168 183 171 186 
rect 168 186 171 189 
rect 168 189 171 192 
rect 168 192 171 195 
rect 168 195 171 198 
rect 168 198 171 201 
rect 168 201 171 204 
rect 168 204 171 207 
rect 168 207 171 210 
rect 168 210 171 213 
rect 168 213 171 216 
rect 168 216 171 219 
rect 168 219 171 222 
rect 168 222 171 225 
rect 168 225 171 228 
rect 168 228 171 231 
rect 168 231 171 234 
rect 168 234 171 237 
rect 168 237 171 240 
rect 168 240 171 243 
rect 168 243 171 246 
rect 168 246 171 249 
rect 168 249 171 252 
rect 168 252 171 255 
rect 168 255 171 258 
rect 168 258 171 261 
rect 168 261 171 264 
rect 168 264 171 267 
rect 168 267 171 270 
rect 168 270 171 273 
rect 168 273 171 276 
rect 168 276 171 279 
rect 168 279 171 282 
rect 168 282 171 285 
rect 168 285 171 288 
rect 168 288 171 291 
rect 168 291 171 294 
rect 168 294 171 297 
rect 168 297 171 300 
rect 168 300 171 303 
rect 168 303 171 306 
rect 168 306 171 309 
rect 168 309 171 312 
rect 168 312 171 315 
rect 168 315 171 318 
rect 168 318 171 321 
rect 168 321 171 324 
rect 168 324 171 327 
rect 168 327 171 330 
rect 168 330 171 333 
rect 168 333 171 336 
rect 168 336 171 339 
rect 168 339 171 342 
rect 168 342 171 345 
rect 168 345 171 348 
rect 168 348 171 351 
rect 168 351 171 354 
rect 168 354 171 357 
rect 168 357 171 360 
rect 168 360 171 363 
rect 168 363 171 366 
rect 168 366 171 369 
rect 168 369 171 372 
rect 168 372 171 375 
rect 168 375 171 378 
rect 168 378 171 381 
rect 168 381 171 384 
rect 168 384 171 387 
rect 168 387 171 390 
rect 168 390 171 393 
rect 168 393 171 396 
rect 168 396 171 399 
rect 168 399 171 402 
rect 168 402 171 405 
rect 168 405 171 408 
rect 168 408 171 411 
rect 168 411 171 414 
rect 168 414 171 417 
rect 168 417 171 420 
rect 168 420 171 423 
rect 168 423 171 426 
rect 168 426 171 429 
rect 168 429 171 432 
rect 168 432 171 435 
rect 168 435 171 438 
rect 168 438 171 441 
rect 168 441 171 444 
rect 168 444 171 447 
rect 168 447 171 450 
rect 168 450 171 453 
rect 168 453 171 456 
rect 168 456 171 459 
rect 168 459 171 462 
rect 168 462 171 465 
rect 168 465 171 468 
rect 168 468 171 471 
rect 168 471 171 474 
rect 168 474 171 477 
rect 168 477 171 480 
rect 168 480 171 483 
rect 168 483 171 486 
rect 168 486 171 489 
rect 168 489 171 492 
rect 168 492 171 495 
rect 168 495 171 498 
rect 168 498 171 501 
rect 168 501 171 504 
rect 168 504 171 507 
rect 168 507 171 510 
rect 171 0 174 3 
rect 171 3 174 6 
rect 171 6 174 9 
rect 171 9 174 12 
rect 171 12 174 15 
rect 171 15 174 18 
rect 171 18 174 21 
rect 171 21 174 24 
rect 171 24 174 27 
rect 171 27 174 30 
rect 171 30 174 33 
rect 171 33 174 36 
rect 171 36 174 39 
rect 171 39 174 42 
rect 171 42 174 45 
rect 171 45 174 48 
rect 171 48 174 51 
rect 171 51 174 54 
rect 171 54 174 57 
rect 171 57 174 60 
rect 171 60 174 63 
rect 171 63 174 66 
rect 171 66 174 69 
rect 171 69 174 72 
rect 171 72 174 75 
rect 171 75 174 78 
rect 171 78 174 81 
rect 171 81 174 84 
rect 171 84 174 87 
rect 171 87 174 90 
rect 171 90 174 93 
rect 171 93 174 96 
rect 171 96 174 99 
rect 171 99 174 102 
rect 171 102 174 105 
rect 171 105 174 108 
rect 171 108 174 111 
rect 171 111 174 114 
rect 171 114 174 117 
rect 171 117 174 120 
rect 171 120 174 123 
rect 171 123 174 126 
rect 171 126 174 129 
rect 171 129 174 132 
rect 171 132 174 135 
rect 171 135 174 138 
rect 171 138 174 141 
rect 171 141 174 144 
rect 171 144 174 147 
rect 171 147 174 150 
rect 171 150 174 153 
rect 171 153 174 156 
rect 171 156 174 159 
rect 171 159 174 162 
rect 171 162 174 165 
rect 171 165 174 168 
rect 171 168 174 171 
rect 171 171 174 174 
rect 171 174 174 177 
rect 171 177 174 180 
rect 171 180 174 183 
rect 171 183 174 186 
rect 171 186 174 189 
rect 171 189 174 192 
rect 171 192 174 195 
rect 171 195 174 198 
rect 171 198 174 201 
rect 171 201 174 204 
rect 171 204 174 207 
rect 171 207 174 210 
rect 171 210 174 213 
rect 171 213 174 216 
rect 171 216 174 219 
rect 171 219 174 222 
rect 171 222 174 225 
rect 171 225 174 228 
rect 171 228 174 231 
rect 171 231 174 234 
rect 171 234 174 237 
rect 171 237 174 240 
rect 171 240 174 243 
rect 171 243 174 246 
rect 171 246 174 249 
rect 171 249 174 252 
rect 171 252 174 255 
rect 171 255 174 258 
rect 171 258 174 261 
rect 171 261 174 264 
rect 171 264 174 267 
rect 171 267 174 270 
rect 171 270 174 273 
rect 171 273 174 276 
rect 171 276 174 279 
rect 171 279 174 282 
rect 171 282 174 285 
rect 171 285 174 288 
rect 171 288 174 291 
rect 171 291 174 294 
rect 171 294 174 297 
rect 171 297 174 300 
rect 171 300 174 303 
rect 171 303 174 306 
rect 171 306 174 309 
rect 171 309 174 312 
rect 171 312 174 315 
rect 171 315 174 318 
rect 171 318 174 321 
rect 171 321 174 324 
rect 171 324 174 327 
rect 171 327 174 330 
rect 171 330 174 333 
rect 171 333 174 336 
rect 171 336 174 339 
rect 171 339 174 342 
rect 171 342 174 345 
rect 171 345 174 348 
rect 171 348 174 351 
rect 171 351 174 354 
rect 171 354 174 357 
rect 171 357 174 360 
rect 171 360 174 363 
rect 171 363 174 366 
rect 171 366 174 369 
rect 171 369 174 372 
rect 171 372 174 375 
rect 171 375 174 378 
rect 171 378 174 381 
rect 171 381 174 384 
rect 171 384 174 387 
rect 171 387 174 390 
rect 171 390 174 393 
rect 171 393 174 396 
rect 171 396 174 399 
rect 171 399 174 402 
rect 171 402 174 405 
rect 171 405 174 408 
rect 171 408 174 411 
rect 171 411 174 414 
rect 171 414 174 417 
rect 171 417 174 420 
rect 171 420 174 423 
rect 171 423 174 426 
rect 171 426 174 429 
rect 171 429 174 432 
rect 171 432 174 435 
rect 171 435 174 438 
rect 171 438 174 441 
rect 171 441 174 444 
rect 171 444 174 447 
rect 171 447 174 450 
rect 171 450 174 453 
rect 171 453 174 456 
rect 171 456 174 459 
rect 171 459 174 462 
rect 171 462 174 465 
rect 171 465 174 468 
rect 171 468 174 471 
rect 171 471 174 474 
rect 171 474 174 477 
rect 171 477 174 480 
rect 171 480 174 483 
rect 171 483 174 486 
rect 171 486 174 489 
rect 171 489 174 492 
rect 171 492 174 495 
rect 171 495 174 498 
rect 171 498 174 501 
rect 171 501 174 504 
rect 171 504 174 507 
rect 171 507 174 510 
rect 174 0 177 3 
rect 174 3 177 6 
rect 174 6 177 9 
rect 174 9 177 12 
rect 174 12 177 15 
rect 174 15 177 18 
rect 174 18 177 21 
rect 174 21 177 24 
rect 174 24 177 27 
rect 174 27 177 30 
rect 174 30 177 33 
rect 174 33 177 36 
rect 174 36 177 39 
rect 174 39 177 42 
rect 174 42 177 45 
rect 174 45 177 48 
rect 174 48 177 51 
rect 174 51 177 54 
rect 174 54 177 57 
rect 174 57 177 60 
rect 174 60 177 63 
rect 174 63 177 66 
rect 174 66 177 69 
rect 174 69 177 72 
rect 174 72 177 75 
rect 174 75 177 78 
rect 174 78 177 81 
rect 174 81 177 84 
rect 174 84 177 87 
rect 174 87 177 90 
rect 174 90 177 93 
rect 174 93 177 96 
rect 174 96 177 99 
rect 174 99 177 102 
rect 174 102 177 105 
rect 174 105 177 108 
rect 174 108 177 111 
rect 174 111 177 114 
rect 174 114 177 117 
rect 174 117 177 120 
rect 174 120 177 123 
rect 174 123 177 126 
rect 174 126 177 129 
rect 174 132 177 135 
rect 174 135 177 138 
rect 174 138 177 141 
rect 174 141 177 144 
rect 174 144 177 147 
rect 174 147 177 150 
rect 174 150 177 153 
rect 174 153 177 156 
rect 174 156 177 159 
rect 174 159 177 162 
rect 174 162 177 165 
rect 174 165 177 168 
rect 174 168 177 171 
rect 174 171 177 174 
rect 174 174 177 177 
rect 174 177 177 180 
rect 174 180 177 183 
rect 174 183 177 186 
rect 174 186 177 189 
rect 174 189 177 192 
rect 174 192 177 195 
rect 174 195 177 198 
rect 174 198 177 201 
rect 174 201 177 204 
rect 174 204 177 207 
rect 174 207 177 210 
rect 174 210 177 213 
rect 174 213 177 216 
rect 174 216 177 219 
rect 174 219 177 222 
rect 174 222 177 225 
rect 174 225 177 228 
rect 174 228 177 231 
rect 174 231 177 234 
rect 174 234 177 237 
rect 174 237 177 240 
rect 174 240 177 243 
rect 174 243 177 246 
rect 174 246 177 249 
rect 174 249 177 252 
rect 174 252 177 255 
rect 174 255 177 258 
rect 174 258 177 261 
rect 174 261 177 264 
rect 174 264 177 267 
rect 174 267 177 270 
rect 174 270 177 273 
rect 174 273 177 276 
rect 174 276 177 279 
rect 174 279 177 282 
rect 174 282 177 285 
rect 174 285 177 288 
rect 174 288 177 291 
rect 174 291 177 294 
rect 174 294 177 297 
rect 174 297 177 300 
rect 174 300 177 303 
rect 174 303 177 306 
rect 174 306 177 309 
rect 174 309 177 312 
rect 174 312 177 315 
rect 174 315 177 318 
rect 174 318 177 321 
rect 174 321 177 324 
rect 174 324 177 327 
rect 174 327 177 330 
rect 174 330 177 333 
rect 174 333 177 336 
rect 174 336 177 339 
rect 174 339 177 342 
rect 174 342 177 345 
rect 174 345 177 348 
rect 174 348 177 351 
rect 174 351 177 354 
rect 174 354 177 357 
rect 174 357 177 360 
rect 174 360 177 363 
rect 174 363 177 366 
rect 174 366 177 369 
rect 174 369 177 372 
rect 174 372 177 375 
rect 174 375 177 378 
rect 174 378 177 381 
rect 174 381 177 384 
rect 174 384 177 387 
rect 174 387 177 390 
rect 174 390 177 393 
rect 174 393 177 396 
rect 174 396 177 399 
rect 174 399 177 402 
rect 174 402 177 405 
rect 174 405 177 408 
rect 174 408 177 411 
rect 174 411 177 414 
rect 174 414 177 417 
rect 174 417 177 420 
rect 174 420 177 423 
rect 174 423 177 426 
rect 174 426 177 429 
rect 174 429 177 432 
rect 174 432 177 435 
rect 174 435 177 438 
rect 174 438 177 441 
rect 174 441 177 444 
rect 174 444 177 447 
rect 174 447 177 450 
rect 174 450 177 453 
rect 174 453 177 456 
rect 174 456 177 459 
rect 174 459 177 462 
rect 174 462 177 465 
rect 174 468 177 471 
rect 174 471 177 474 
rect 174 474 177 477 
rect 174 477 177 480 
rect 174 480 177 483 
rect 174 483 177 486 
rect 174 486 177 489 
rect 174 489 177 492 
rect 174 492 177 495 
rect 174 495 177 498 
rect 174 498 177 501 
rect 174 501 177 504 
rect 174 504 177 507 
rect 174 507 177 510 
rect 177 0 180 3 
rect 177 3 180 6 
rect 177 6 180 9 
rect 177 9 180 12 
rect 177 12 180 15 
rect 177 15 180 18 
rect 177 18 180 21 
rect 177 21 180 24 
rect 177 24 180 27 
rect 177 27 180 30 
rect 177 30 180 33 
rect 177 33 180 36 
rect 177 36 180 39 
rect 177 39 180 42 
rect 177 42 180 45 
rect 177 45 180 48 
rect 177 48 180 51 
rect 177 51 180 54 
rect 177 54 180 57 
rect 177 57 180 60 
rect 177 60 180 63 
rect 177 63 180 66 
rect 177 66 180 69 
rect 177 69 180 72 
rect 177 72 180 75 
rect 177 75 180 78 
rect 177 78 180 81 
rect 177 81 180 84 
rect 177 84 180 87 
rect 177 87 180 90 
rect 177 90 180 93 
rect 177 93 180 96 
rect 177 96 180 99 
rect 177 99 180 102 
rect 177 102 180 105 
rect 177 105 180 108 
rect 177 108 180 111 
rect 177 111 180 114 
rect 177 114 180 117 
rect 177 117 180 120 
rect 177 120 180 123 
rect 177 123 180 126 
rect 177 126 180 129 
rect 177 129 180 132 
rect 177 132 180 135 
rect 177 135 180 138 
rect 177 138 180 141 
rect 177 141 180 144 
rect 177 144 180 147 
rect 177 147 180 150 
rect 177 150 180 153 
rect 177 153 180 156 
rect 177 156 180 159 
rect 177 159 180 162 
rect 177 162 180 165 
rect 177 165 180 168 
rect 177 168 180 171 
rect 177 171 180 174 
rect 177 174 180 177 
rect 177 177 180 180 
rect 177 180 180 183 
rect 177 183 180 186 
rect 177 186 180 189 
rect 177 189 180 192 
rect 177 192 180 195 
rect 177 195 180 198 
rect 177 198 180 201 
rect 177 201 180 204 
rect 177 204 180 207 
rect 177 207 180 210 
rect 177 210 180 213 
rect 177 213 180 216 
rect 177 216 180 219 
rect 177 219 180 222 
rect 177 222 180 225 
rect 177 225 180 228 
rect 177 228 180 231 
rect 177 231 180 234 
rect 177 234 180 237 
rect 177 237 180 240 
rect 177 240 180 243 
rect 177 243 180 246 
rect 177 246 180 249 
rect 177 249 180 252 
rect 177 252 180 255 
rect 177 255 180 258 
rect 177 258 180 261 
rect 177 261 180 264 
rect 177 264 180 267 
rect 177 267 180 270 
rect 177 270 180 273 
rect 177 273 180 276 
rect 177 276 180 279 
rect 177 279 180 282 
rect 177 282 180 285 
rect 177 285 180 288 
rect 177 288 180 291 
rect 177 291 180 294 
rect 177 294 180 297 
rect 177 297 180 300 
rect 177 300 180 303 
rect 177 303 180 306 
rect 177 306 180 309 
rect 177 309 180 312 
rect 177 312 180 315 
rect 177 315 180 318 
rect 177 318 180 321 
rect 177 321 180 324 
rect 177 324 180 327 
rect 177 327 180 330 
rect 177 330 180 333 
rect 177 333 180 336 
rect 177 336 180 339 
rect 177 339 180 342 
rect 177 342 180 345 
rect 177 345 180 348 
rect 177 348 180 351 
rect 177 351 180 354 
rect 177 354 180 357 
rect 177 357 180 360 
rect 177 360 180 363 
rect 177 363 180 366 
rect 177 366 180 369 
rect 177 369 180 372 
rect 177 372 180 375 
rect 177 375 180 378 
rect 177 378 180 381 
rect 177 381 180 384 
rect 177 384 180 387 
rect 177 387 180 390 
rect 177 390 180 393 
rect 177 393 180 396 
rect 177 396 180 399 
rect 177 399 180 402 
rect 177 402 180 405 
rect 177 405 180 408 
rect 177 408 180 411 
rect 177 411 180 414 
rect 177 414 180 417 
rect 177 417 180 420 
rect 177 420 180 423 
rect 177 423 180 426 
rect 177 426 180 429 
rect 177 429 180 432 
rect 177 432 180 435 
rect 177 435 180 438 
rect 177 438 180 441 
rect 177 441 180 444 
rect 177 444 180 447 
rect 177 447 180 450 
rect 177 450 180 453 
rect 177 453 180 456 
rect 177 456 180 459 
rect 177 459 180 462 
rect 177 462 180 465 
rect 177 465 180 468 
rect 177 468 180 471 
rect 177 471 180 474 
rect 177 474 180 477 
rect 177 477 180 480 
rect 177 480 180 483 
rect 177 483 180 486 
rect 177 486 180 489 
rect 177 489 180 492 
rect 177 492 180 495 
rect 177 495 180 498 
rect 177 498 180 501 
rect 177 501 180 504 
rect 177 504 180 507 
rect 177 507 180 510 
rect 180 0 183 3 
rect 180 3 183 6 
rect 180 6 183 9 
rect 180 9 183 12 
rect 180 12 183 15 
rect 180 15 183 18 
rect 180 18 183 21 
rect 180 21 183 24 
rect 180 24 183 27 
rect 180 27 183 30 
rect 180 30 183 33 
rect 180 33 183 36 
rect 180 36 183 39 
rect 180 39 183 42 
rect 180 42 183 45 
rect 180 45 183 48 
rect 180 48 183 51 
rect 180 51 183 54 
rect 180 54 183 57 
rect 180 57 183 60 
rect 180 60 183 63 
rect 180 63 183 66 
rect 180 66 183 69 
rect 180 69 183 72 
rect 180 72 183 75 
rect 180 75 183 78 
rect 180 78 183 81 
rect 180 81 183 84 
rect 180 84 183 87 
rect 180 87 183 90 
rect 180 90 183 93 
rect 180 93 183 96 
rect 180 96 183 99 
rect 180 99 183 102 
rect 180 102 183 105 
rect 180 105 183 108 
rect 180 108 183 111 
rect 180 111 183 114 
rect 180 114 183 117 
rect 180 117 183 120 
rect 180 120 183 123 
rect 180 123 183 126 
rect 180 126 183 129 
rect 180 129 183 132 
rect 180 132 183 135 
rect 180 135 183 138 
rect 180 138 183 141 
rect 180 141 183 144 
rect 180 144 183 147 
rect 180 147 183 150 
rect 180 150 183 153 
rect 180 153 183 156 
rect 180 156 183 159 
rect 180 159 183 162 
rect 180 162 183 165 
rect 180 165 183 168 
rect 180 168 183 171 
rect 180 171 183 174 
rect 180 174 183 177 
rect 180 177 183 180 
rect 180 180 183 183 
rect 180 183 183 186 
rect 180 186 183 189 
rect 180 189 183 192 
rect 180 192 183 195 
rect 180 195 183 198 
rect 180 198 183 201 
rect 180 201 183 204 
rect 180 204 183 207 
rect 180 207 183 210 
rect 180 210 183 213 
rect 180 213 183 216 
rect 180 216 183 219 
rect 180 219 183 222 
rect 180 222 183 225 
rect 180 225 183 228 
rect 180 228 183 231 
rect 180 231 183 234 
rect 180 234 183 237 
rect 180 237 183 240 
rect 180 240 183 243 
rect 180 243 183 246 
rect 180 246 183 249 
rect 180 249 183 252 
rect 180 252 183 255 
rect 180 255 183 258 
rect 180 258 183 261 
rect 180 261 183 264 
rect 180 264 183 267 
rect 180 267 183 270 
rect 180 270 183 273 
rect 180 273 183 276 
rect 180 276 183 279 
rect 180 279 183 282 
rect 180 282 183 285 
rect 180 285 183 288 
rect 180 288 183 291 
rect 180 291 183 294 
rect 180 294 183 297 
rect 180 297 183 300 
rect 180 300 183 303 
rect 180 303 183 306 
rect 180 306 183 309 
rect 180 309 183 312 
rect 180 312 183 315 
rect 180 315 183 318 
rect 180 318 183 321 
rect 180 321 183 324 
rect 180 324 183 327 
rect 180 327 183 330 
rect 180 330 183 333 
rect 180 333 183 336 
rect 180 336 183 339 
rect 180 339 183 342 
rect 180 342 183 345 
rect 180 345 183 348 
rect 180 348 183 351 
rect 180 351 183 354 
rect 180 354 183 357 
rect 180 357 183 360 
rect 180 360 183 363 
rect 180 363 183 366 
rect 180 366 183 369 
rect 180 369 183 372 
rect 180 372 183 375 
rect 180 375 183 378 
rect 180 378 183 381 
rect 180 381 183 384 
rect 180 384 183 387 
rect 180 387 183 390 
rect 180 390 183 393 
rect 180 393 183 396 
rect 180 396 183 399 
rect 180 399 183 402 
rect 180 402 183 405 
rect 180 405 183 408 
rect 180 408 183 411 
rect 180 411 183 414 
rect 180 414 183 417 
rect 180 417 183 420 
rect 180 420 183 423 
rect 180 423 183 426 
rect 180 426 183 429 
rect 180 429 183 432 
rect 180 432 183 435 
rect 180 435 183 438 
rect 180 438 183 441 
rect 180 441 183 444 
rect 180 444 183 447 
rect 180 447 183 450 
rect 180 450 183 453 
rect 180 453 183 456 
rect 180 456 183 459 
rect 180 459 183 462 
rect 180 462 183 465 
rect 180 465 183 468 
rect 180 468 183 471 
rect 180 471 183 474 
rect 180 474 183 477 
rect 180 477 183 480 
rect 180 480 183 483 
rect 180 483 183 486 
rect 180 486 183 489 
rect 180 489 183 492 
rect 180 492 183 495 
rect 180 495 183 498 
rect 180 498 183 501 
rect 180 501 183 504 
rect 180 504 183 507 
rect 180 507 183 510 
rect 183 0 186 3 
rect 183 3 186 6 
rect 183 6 186 9 
rect 183 9 186 12 
rect 183 12 186 15 
rect 183 15 186 18 
rect 183 18 186 21 
rect 183 21 186 24 
rect 183 24 186 27 
rect 183 27 186 30 
rect 183 30 186 33 
rect 183 33 186 36 
rect 183 36 186 39 
rect 183 39 186 42 
rect 183 42 186 45 
rect 183 45 186 48 
rect 183 48 186 51 
rect 183 51 186 54 
rect 183 54 186 57 
rect 183 57 186 60 
rect 183 60 186 63 
rect 183 63 186 66 
rect 183 66 186 69 
rect 183 69 186 72 
rect 183 72 186 75 
rect 183 75 186 78 
rect 183 78 186 81 
rect 183 81 186 84 
rect 183 84 186 87 
rect 183 87 186 90 
rect 183 90 186 93 
rect 183 93 186 96 
rect 183 96 186 99 
rect 183 99 186 102 
rect 183 102 186 105 
rect 183 105 186 108 
rect 183 108 186 111 
rect 183 111 186 114 
rect 183 114 186 117 
rect 183 117 186 120 
rect 183 120 186 123 
rect 183 123 186 126 
rect 183 126 186 129 
rect 183 129 186 132 
rect 183 132 186 135 
rect 183 135 186 138 
rect 183 138 186 141 
rect 183 141 186 144 
rect 183 144 186 147 
rect 183 147 186 150 
rect 183 150 186 153 
rect 183 153 186 156 
rect 183 156 186 159 
rect 183 159 186 162 
rect 183 162 186 165 
rect 183 165 186 168 
rect 183 168 186 171 
rect 183 171 186 174 
rect 183 174 186 177 
rect 183 177 186 180 
rect 183 180 186 183 
rect 183 183 186 186 
rect 183 186 186 189 
rect 183 189 186 192 
rect 183 192 186 195 
rect 183 195 186 198 
rect 183 198 186 201 
rect 183 201 186 204 
rect 183 204 186 207 
rect 183 207 186 210 
rect 183 210 186 213 
rect 183 213 186 216 
rect 183 216 186 219 
rect 183 219 186 222 
rect 183 222 186 225 
rect 183 225 186 228 
rect 183 228 186 231 
rect 183 231 186 234 
rect 183 234 186 237 
rect 183 237 186 240 
rect 183 240 186 243 
rect 183 243 186 246 
rect 183 246 186 249 
rect 183 249 186 252 
rect 183 252 186 255 
rect 183 255 186 258 
rect 183 258 186 261 
rect 183 261 186 264 
rect 183 264 186 267 
rect 183 267 186 270 
rect 183 270 186 273 
rect 183 273 186 276 
rect 183 276 186 279 
rect 183 279 186 282 
rect 183 282 186 285 
rect 183 285 186 288 
rect 183 288 186 291 
rect 183 291 186 294 
rect 183 294 186 297 
rect 183 297 186 300 
rect 183 300 186 303 
rect 183 303 186 306 
rect 183 306 186 309 
rect 183 309 186 312 
rect 183 312 186 315 
rect 183 315 186 318 
rect 183 318 186 321 
rect 183 321 186 324 
rect 183 324 186 327 
rect 183 327 186 330 
rect 183 330 186 333 
rect 183 333 186 336 
rect 183 336 186 339 
rect 183 339 186 342 
rect 183 342 186 345 
rect 183 345 186 348 
rect 183 348 186 351 
rect 183 351 186 354 
rect 183 354 186 357 
rect 183 357 186 360 
rect 183 360 186 363 
rect 183 363 186 366 
rect 183 366 186 369 
rect 183 369 186 372 
rect 183 372 186 375 
rect 183 375 186 378 
rect 183 378 186 381 
rect 183 381 186 384 
rect 183 384 186 387 
rect 183 387 186 390 
rect 183 390 186 393 
rect 183 393 186 396 
rect 183 396 186 399 
rect 183 399 186 402 
rect 183 402 186 405 
rect 183 405 186 408 
rect 183 408 186 411 
rect 183 411 186 414 
rect 183 414 186 417 
rect 183 417 186 420 
rect 183 420 186 423 
rect 183 423 186 426 
rect 183 426 186 429 
rect 183 429 186 432 
rect 183 432 186 435 
rect 183 435 186 438 
rect 183 438 186 441 
rect 183 441 186 444 
rect 183 444 186 447 
rect 183 447 186 450 
rect 183 450 186 453 
rect 183 453 186 456 
rect 183 456 186 459 
rect 183 459 186 462 
rect 183 462 186 465 
rect 183 465 186 468 
rect 183 468 186 471 
rect 183 471 186 474 
rect 183 474 186 477 
rect 183 477 186 480 
rect 183 480 186 483 
rect 183 483 186 486 
rect 183 486 186 489 
rect 183 489 186 492 
rect 183 492 186 495 
rect 183 495 186 498 
rect 183 498 186 501 
rect 183 501 186 504 
rect 183 504 186 507 
rect 183 507 186 510 
rect 186 0 189 3 
rect 186 3 189 6 
rect 186 6 189 9 
rect 186 9 189 12 
rect 186 12 189 15 
rect 186 15 189 18 
rect 186 18 189 21 
rect 186 21 189 24 
rect 186 24 189 27 
rect 186 27 189 30 
rect 186 30 189 33 
rect 186 33 189 36 
rect 186 36 189 39 
rect 186 39 189 42 
rect 186 42 189 45 
rect 186 45 189 48 
rect 186 48 189 51 
rect 186 51 189 54 
rect 186 54 189 57 
rect 186 57 189 60 
rect 186 60 189 63 
rect 186 63 189 66 
rect 186 66 189 69 
rect 186 69 189 72 
rect 186 72 189 75 
rect 186 75 189 78 
rect 186 78 189 81 
rect 186 81 189 84 
rect 186 84 189 87 
rect 186 87 189 90 
rect 186 90 189 93 
rect 186 93 189 96 
rect 186 96 189 99 
rect 186 99 189 102 
rect 186 102 189 105 
rect 186 105 189 108 
rect 186 108 189 111 
rect 186 111 189 114 
rect 186 114 189 117 
rect 186 117 189 120 
rect 186 120 189 123 
rect 186 123 189 126 
rect 186 126 189 129 
rect 186 129 189 132 
rect 186 132 189 135 
rect 186 135 189 138 
rect 186 138 189 141 
rect 186 141 189 144 
rect 186 144 189 147 
rect 186 147 189 150 
rect 186 150 189 153 
rect 186 153 189 156 
rect 186 156 189 159 
rect 186 159 189 162 
rect 186 162 189 165 
rect 186 165 189 168 
rect 186 168 189 171 
rect 186 171 189 174 
rect 186 174 189 177 
rect 186 177 189 180 
rect 186 180 189 183 
rect 186 183 189 186 
rect 186 186 189 189 
rect 186 189 189 192 
rect 186 192 189 195 
rect 186 195 189 198 
rect 186 198 189 201 
rect 186 201 189 204 
rect 186 204 189 207 
rect 186 207 189 210 
rect 186 210 189 213 
rect 186 213 189 216 
rect 186 216 189 219 
rect 186 219 189 222 
rect 186 222 189 225 
rect 186 225 189 228 
rect 186 228 189 231 
rect 186 231 189 234 
rect 186 234 189 237 
rect 186 237 189 240 
rect 186 240 189 243 
rect 186 243 189 246 
rect 186 246 189 249 
rect 186 249 189 252 
rect 186 252 189 255 
rect 186 255 189 258 
rect 186 258 189 261 
rect 186 261 189 264 
rect 186 264 189 267 
rect 186 267 189 270 
rect 186 270 189 273 
rect 186 273 189 276 
rect 186 276 189 279 
rect 186 279 189 282 
rect 186 282 189 285 
rect 186 285 189 288 
rect 186 288 189 291 
rect 186 291 189 294 
rect 186 294 189 297 
rect 186 297 189 300 
rect 186 300 189 303 
rect 186 303 189 306 
rect 186 306 189 309 
rect 186 309 189 312 
rect 186 312 189 315 
rect 186 315 189 318 
rect 186 318 189 321 
rect 186 321 189 324 
rect 186 324 189 327 
rect 186 327 189 330 
rect 186 330 189 333 
rect 186 333 189 336 
rect 186 336 189 339 
rect 186 339 189 342 
rect 186 342 189 345 
rect 186 345 189 348 
rect 186 348 189 351 
rect 186 351 189 354 
rect 186 354 189 357 
rect 186 357 189 360 
rect 186 360 189 363 
rect 186 363 189 366 
rect 186 366 189 369 
rect 186 369 189 372 
rect 186 372 189 375 
rect 186 375 189 378 
rect 186 378 189 381 
rect 186 381 189 384 
rect 186 384 189 387 
rect 186 387 189 390 
rect 186 390 189 393 
rect 186 393 189 396 
rect 186 396 189 399 
rect 186 399 189 402 
rect 186 402 189 405 
rect 186 405 189 408 
rect 186 408 189 411 
rect 186 411 189 414 
rect 186 414 189 417 
rect 186 417 189 420 
rect 186 420 189 423 
rect 186 423 189 426 
rect 186 426 189 429 
rect 186 429 189 432 
rect 186 432 189 435 
rect 186 435 189 438 
rect 186 438 189 441 
rect 186 441 189 444 
rect 186 444 189 447 
rect 186 447 189 450 
rect 186 450 189 453 
rect 186 453 189 456 
rect 186 456 189 459 
rect 186 459 189 462 
rect 186 462 189 465 
rect 186 465 189 468 
rect 186 468 189 471 
rect 186 471 189 474 
rect 186 474 189 477 
rect 186 477 189 480 
rect 186 480 189 483 
rect 186 483 189 486 
rect 186 486 189 489 
rect 186 489 189 492 
rect 186 492 189 495 
rect 186 495 189 498 
rect 186 498 189 501 
rect 186 501 189 504 
rect 186 504 189 507 
rect 186 507 189 510 
rect 189 0 192 3 
rect 189 3 192 6 
rect 189 6 192 9 
rect 189 9 192 12 
rect 189 12 192 15 
rect 189 15 192 18 
rect 189 18 192 21 
rect 189 21 192 24 
rect 189 24 192 27 
rect 189 27 192 30 
rect 189 30 192 33 
rect 189 36 192 39 
rect 189 39 192 42 
rect 189 42 192 45 
rect 189 45 192 48 
rect 189 48 192 51 
rect 189 51 192 54 
rect 189 54 192 57 
rect 189 57 192 60 
rect 189 60 192 63 
rect 189 63 192 66 
rect 189 66 192 69 
rect 189 69 192 72 
rect 189 72 192 75 
rect 189 75 192 78 
rect 189 78 192 81 
rect 189 84 192 87 
rect 189 87 192 90 
rect 189 93 192 96 
rect 189 96 192 99 
rect 189 99 192 102 
rect 189 102 192 105 
rect 189 105 192 108 
rect 189 108 192 111 
rect 189 111 192 114 
rect 189 114 192 117 
rect 189 117 192 120 
rect 189 120 192 123 
rect 189 123 192 126 
rect 189 126 192 129 
rect 189 132 192 135 
rect 189 135 192 138 
rect 189 138 192 141 
rect 189 141 192 144 
rect 189 144 192 147 
rect 189 147 192 150 
rect 189 150 192 153 
rect 189 153 192 156 
rect 189 156 192 159 
rect 189 159 192 162 
rect 189 162 192 165 
rect 189 165 192 168 
rect 189 168 192 171 
rect 189 171 192 174 
rect 189 174 192 177 
rect 189 177 192 180 
rect 189 180 192 183 
rect 189 183 192 186 
rect 189 186 192 189 
rect 189 189 192 192 
rect 189 192 192 195 
rect 189 195 192 198 
rect 189 198 192 201 
rect 189 201 192 204 
rect 189 204 192 207 
rect 189 207 192 210 
rect 189 210 192 213 
rect 189 213 192 216 
rect 189 216 192 219 
rect 189 219 192 222 
rect 189 222 192 225 
rect 189 225 192 228 
rect 189 228 192 231 
rect 189 231 192 234 
rect 189 234 192 237 
rect 189 237 192 240 
rect 189 240 192 243 
rect 189 243 192 246 
rect 189 246 192 249 
rect 189 249 192 252 
rect 189 252 192 255 
rect 189 255 192 258 
rect 189 258 192 261 
rect 189 261 192 264 
rect 189 264 192 267 
rect 189 267 192 270 
rect 189 270 192 273 
rect 189 273 192 276 
rect 189 276 192 279 
rect 189 279 192 282 
rect 189 282 192 285 
rect 189 285 192 288 
rect 189 288 192 291 
rect 189 291 192 294 
rect 189 294 192 297 
rect 189 297 192 300 
rect 189 300 192 303 
rect 189 303 192 306 
rect 189 306 192 309 
rect 189 309 192 312 
rect 189 312 192 315 
rect 189 315 192 318 
rect 189 318 192 321 
rect 189 321 192 324 
rect 189 324 192 327 
rect 189 327 192 330 
rect 189 330 192 333 
rect 189 333 192 336 
rect 189 336 192 339 
rect 189 339 192 342 
rect 189 342 192 345 
rect 189 345 192 348 
rect 189 348 192 351 
rect 189 351 192 354 
rect 189 354 192 357 
rect 189 357 192 360 
rect 189 360 192 363 
rect 189 363 192 366 
rect 189 366 192 369 
rect 189 369 192 372 
rect 189 372 192 375 
rect 189 375 192 378 
rect 189 378 192 381 
rect 189 381 192 384 
rect 189 384 192 387 
rect 189 387 192 390 
rect 189 390 192 393 
rect 189 393 192 396 
rect 189 396 192 399 
rect 189 399 192 402 
rect 189 402 192 405 
rect 189 405 192 408 
rect 189 408 192 411 
rect 189 411 192 414 
rect 189 414 192 417 
rect 189 417 192 420 
rect 189 420 192 423 
rect 189 423 192 426 
rect 189 429 192 432 
rect 189 432 192 435 
rect 189 435 192 438 
rect 189 438 192 441 
rect 189 441 192 444 
rect 189 444 192 447 
rect 189 447 192 450 
rect 189 450 192 453 
rect 189 453 192 456 
rect 189 456 192 459 
rect 189 459 192 462 
rect 189 462 192 465 
rect 189 465 192 468 
rect 189 468 192 471 
rect 189 471 192 474 
rect 189 477 192 480 
rect 189 480 192 483 
rect 189 483 192 486 
rect 189 486 192 489 
rect 189 489 192 492 
rect 189 492 192 495 
rect 189 495 192 498 
rect 189 498 192 501 
rect 189 501 192 504 
rect 189 504 192 507 
rect 189 507 192 510 
rect 192 0 195 3 
rect 192 3 195 6 
rect 192 6 195 9 
rect 192 9 195 12 
rect 192 12 195 15 
rect 192 15 195 18 
rect 192 18 195 21 
rect 192 21 195 24 
rect 192 24 195 27 
rect 192 27 195 30 
rect 192 30 195 33 
rect 192 33 195 36 
rect 192 36 195 39 
rect 192 39 195 42 
rect 192 42 195 45 
rect 192 45 195 48 
rect 192 48 195 51 
rect 192 51 195 54 
rect 192 54 195 57 
rect 192 57 195 60 
rect 192 60 195 63 
rect 192 63 195 66 
rect 192 66 195 69 
rect 192 69 195 72 
rect 192 72 195 75 
rect 192 75 195 78 
rect 192 78 195 81 
rect 192 81 195 84 
rect 192 84 195 87 
rect 192 87 195 90 
rect 192 90 195 93 
rect 192 93 195 96 
rect 192 96 195 99 
rect 192 99 195 102 
rect 192 102 195 105 
rect 192 105 195 108 
rect 192 108 195 111 
rect 192 111 195 114 
rect 192 114 195 117 
rect 192 117 195 120 
rect 192 120 195 123 
rect 192 123 195 126 
rect 192 126 195 129 
rect 192 129 195 132 
rect 192 132 195 135 
rect 192 135 195 138 
rect 192 138 195 141 
rect 192 141 195 144 
rect 192 144 195 147 
rect 192 147 195 150 
rect 192 150 195 153 
rect 192 153 195 156 
rect 192 156 195 159 
rect 192 159 195 162 
rect 192 162 195 165 
rect 192 165 195 168 
rect 192 168 195 171 
rect 192 171 195 174 
rect 192 174 195 177 
rect 192 177 195 180 
rect 192 180 195 183 
rect 192 183 195 186 
rect 192 186 195 189 
rect 192 189 195 192 
rect 192 192 195 195 
rect 192 195 195 198 
rect 192 198 195 201 
rect 192 201 195 204 
rect 192 204 195 207 
rect 192 207 195 210 
rect 192 210 195 213 
rect 192 213 195 216 
rect 192 216 195 219 
rect 192 219 195 222 
rect 192 222 195 225 
rect 192 225 195 228 
rect 192 228 195 231 
rect 192 231 195 234 
rect 192 234 195 237 
rect 192 237 195 240 
rect 192 240 195 243 
rect 192 243 195 246 
rect 192 246 195 249 
rect 192 249 195 252 
rect 192 252 195 255 
rect 192 255 195 258 
rect 192 258 195 261 
rect 192 261 195 264 
rect 192 264 195 267 
rect 192 267 195 270 
rect 192 270 195 273 
rect 192 273 195 276 
rect 192 276 195 279 
rect 192 279 195 282 
rect 192 282 195 285 
rect 192 285 195 288 
rect 192 288 195 291 
rect 192 291 195 294 
rect 192 294 195 297 
rect 192 297 195 300 
rect 192 300 195 303 
rect 192 303 195 306 
rect 192 306 195 309 
rect 192 309 195 312 
rect 192 312 195 315 
rect 192 315 195 318 
rect 192 318 195 321 
rect 192 321 195 324 
rect 192 324 195 327 
rect 192 327 195 330 
rect 192 330 195 333 
rect 192 333 195 336 
rect 192 336 195 339 
rect 192 339 195 342 
rect 192 342 195 345 
rect 192 345 195 348 
rect 192 348 195 351 
rect 192 351 195 354 
rect 192 354 195 357 
rect 192 357 195 360 
rect 192 360 195 363 
rect 192 363 195 366 
rect 192 366 195 369 
rect 192 369 195 372 
rect 192 372 195 375 
rect 192 375 195 378 
rect 192 378 195 381 
rect 192 381 195 384 
rect 192 384 195 387 
rect 192 387 195 390 
rect 192 390 195 393 
rect 192 393 195 396 
rect 192 396 195 399 
rect 192 399 195 402 
rect 192 402 195 405 
rect 192 405 195 408 
rect 192 408 195 411 
rect 192 411 195 414 
rect 192 414 195 417 
rect 192 417 195 420 
rect 192 420 195 423 
rect 192 423 195 426 
rect 192 426 195 429 
rect 192 429 195 432 
rect 192 432 195 435 
rect 192 435 195 438 
rect 192 438 195 441 
rect 192 441 195 444 
rect 192 444 195 447 
rect 192 447 195 450 
rect 192 450 195 453 
rect 192 453 195 456 
rect 192 456 195 459 
rect 192 459 195 462 
rect 192 462 195 465 
rect 192 465 195 468 
rect 192 468 195 471 
rect 192 471 195 474 
rect 192 474 195 477 
rect 192 477 195 480 
rect 192 480 195 483 
rect 192 483 195 486 
rect 192 486 195 489 
rect 192 489 195 492 
rect 192 492 195 495 
rect 192 495 195 498 
rect 192 498 195 501 
rect 192 501 195 504 
rect 192 504 195 507 
rect 192 507 195 510 
rect 195 0 198 3 
rect 195 3 198 6 
rect 195 6 198 9 
rect 195 9 198 12 
rect 195 12 198 15 
rect 195 15 198 18 
rect 195 18 198 21 
rect 195 21 198 24 
rect 195 24 198 27 
rect 195 27 198 30 
rect 195 30 198 33 
rect 195 33 198 36 
rect 195 36 198 39 
rect 195 39 198 42 
rect 195 42 198 45 
rect 195 45 198 48 
rect 195 48 198 51 
rect 195 51 198 54 
rect 195 54 198 57 
rect 195 57 198 60 
rect 195 60 198 63 
rect 195 63 198 66 
rect 195 66 198 69 
rect 195 69 198 72 
rect 195 72 198 75 
rect 195 75 198 78 
rect 195 78 198 81 
rect 195 81 198 84 
rect 195 84 198 87 
rect 195 87 198 90 
rect 195 90 198 93 
rect 195 93 198 96 
rect 195 96 198 99 
rect 195 99 198 102 
rect 195 102 198 105 
rect 195 105 198 108 
rect 195 108 198 111 
rect 195 111 198 114 
rect 195 114 198 117 
rect 195 117 198 120 
rect 195 120 198 123 
rect 195 123 198 126 
rect 195 126 198 129 
rect 195 129 198 132 
rect 195 132 198 135 
rect 195 135 198 138 
rect 195 138 198 141 
rect 195 141 198 144 
rect 195 144 198 147 
rect 195 147 198 150 
rect 195 150 198 153 
rect 195 153 198 156 
rect 195 156 198 159 
rect 195 159 198 162 
rect 195 162 198 165 
rect 195 165 198 168 
rect 195 168 198 171 
rect 195 171 198 174 
rect 195 174 198 177 
rect 195 177 198 180 
rect 195 180 198 183 
rect 195 183 198 186 
rect 195 186 198 189 
rect 195 189 198 192 
rect 195 192 198 195 
rect 195 195 198 198 
rect 195 198 198 201 
rect 195 201 198 204 
rect 195 204 198 207 
rect 195 207 198 210 
rect 195 210 198 213 
rect 195 213 198 216 
rect 195 216 198 219 
rect 195 219 198 222 
rect 195 222 198 225 
rect 195 225 198 228 
rect 195 228 198 231 
rect 195 231 198 234 
rect 195 234 198 237 
rect 195 237 198 240 
rect 195 240 198 243 
rect 195 243 198 246 
rect 195 246 198 249 
rect 195 249 198 252 
rect 195 252 198 255 
rect 195 255 198 258 
rect 195 258 198 261 
rect 195 261 198 264 
rect 195 264 198 267 
rect 195 267 198 270 
rect 195 270 198 273 
rect 195 273 198 276 
rect 195 276 198 279 
rect 195 279 198 282 
rect 195 282 198 285 
rect 195 285 198 288 
rect 195 288 198 291 
rect 195 291 198 294 
rect 195 294 198 297 
rect 195 297 198 300 
rect 195 300 198 303 
rect 195 303 198 306 
rect 195 306 198 309 
rect 195 309 198 312 
rect 195 312 198 315 
rect 195 315 198 318 
rect 195 318 198 321 
rect 195 321 198 324 
rect 195 324 198 327 
rect 195 327 198 330 
rect 195 330 198 333 
rect 195 333 198 336 
rect 195 336 198 339 
rect 195 339 198 342 
rect 195 342 198 345 
rect 195 345 198 348 
rect 195 348 198 351 
rect 195 351 198 354 
rect 195 354 198 357 
rect 195 357 198 360 
rect 195 360 198 363 
rect 195 363 198 366 
rect 195 366 198 369 
rect 195 369 198 372 
rect 195 372 198 375 
rect 195 375 198 378 
rect 195 378 198 381 
rect 195 381 198 384 
rect 195 384 198 387 
rect 195 387 198 390 
rect 195 390 198 393 
rect 195 393 198 396 
rect 195 396 198 399 
rect 195 399 198 402 
rect 195 402 198 405 
rect 195 405 198 408 
rect 195 408 198 411 
rect 195 411 198 414 
rect 195 414 198 417 
rect 195 417 198 420 
rect 195 420 198 423 
rect 195 423 198 426 
rect 195 426 198 429 
rect 195 429 198 432 
rect 195 432 198 435 
rect 195 435 198 438 
rect 195 438 198 441 
rect 195 441 198 444 
rect 195 444 198 447 
rect 195 447 198 450 
rect 195 450 198 453 
rect 195 453 198 456 
rect 195 456 198 459 
rect 195 459 198 462 
rect 195 462 198 465 
rect 195 465 198 468 
rect 195 468 198 471 
rect 195 471 198 474 
rect 195 474 198 477 
rect 195 477 198 480 
rect 195 480 198 483 
rect 195 483 198 486 
rect 195 486 198 489 
rect 195 489 198 492 
rect 195 492 198 495 
rect 195 495 198 498 
rect 195 498 198 501 
rect 195 501 198 504 
rect 195 504 198 507 
rect 195 507 198 510 
rect 198 0 201 3 
rect 198 3 201 6 
rect 198 6 201 9 
rect 198 9 201 12 
rect 198 12 201 15 
rect 198 15 201 18 
rect 198 18 201 21 
rect 198 21 201 24 
rect 198 24 201 27 
rect 198 27 201 30 
rect 198 30 201 33 
rect 198 33 201 36 
rect 198 36 201 39 
rect 198 39 201 42 
rect 198 42 201 45 
rect 198 45 201 48 
rect 198 48 201 51 
rect 198 51 201 54 
rect 198 54 201 57 
rect 198 57 201 60 
rect 198 60 201 63 
rect 198 63 201 66 
rect 198 66 201 69 
rect 198 69 201 72 
rect 198 72 201 75 
rect 198 75 201 78 
rect 198 78 201 81 
rect 198 81 201 84 
rect 198 84 201 87 
rect 198 87 201 90 
rect 198 90 201 93 
rect 198 93 201 96 
rect 198 96 201 99 
rect 198 99 201 102 
rect 198 102 201 105 
rect 198 105 201 108 
rect 198 108 201 111 
rect 198 111 201 114 
rect 198 114 201 117 
rect 198 117 201 120 
rect 198 120 201 123 
rect 198 123 201 126 
rect 198 126 201 129 
rect 198 129 201 132 
rect 198 132 201 135 
rect 198 135 201 138 
rect 198 138 201 141 
rect 198 141 201 144 
rect 198 144 201 147 
rect 198 147 201 150 
rect 198 150 201 153 
rect 198 153 201 156 
rect 198 156 201 159 
rect 198 159 201 162 
rect 198 162 201 165 
rect 198 165 201 168 
rect 198 168 201 171 
rect 198 171 201 174 
rect 198 174 201 177 
rect 198 177 201 180 
rect 198 180 201 183 
rect 198 183 201 186 
rect 198 186 201 189 
rect 198 189 201 192 
rect 198 192 201 195 
rect 198 195 201 198 
rect 198 198 201 201 
rect 198 201 201 204 
rect 198 204 201 207 
rect 198 207 201 210 
rect 198 210 201 213 
rect 198 213 201 216 
rect 198 216 201 219 
rect 198 219 201 222 
rect 198 222 201 225 
rect 198 225 201 228 
rect 198 228 201 231 
rect 198 231 201 234 
rect 198 234 201 237 
rect 198 237 201 240 
rect 198 240 201 243 
rect 198 243 201 246 
rect 198 246 201 249 
rect 198 249 201 252 
rect 198 252 201 255 
rect 198 255 201 258 
rect 198 258 201 261 
rect 198 261 201 264 
rect 198 264 201 267 
rect 198 267 201 270 
rect 198 270 201 273 
rect 198 273 201 276 
rect 198 276 201 279 
rect 198 279 201 282 
rect 198 282 201 285 
rect 198 285 201 288 
rect 198 288 201 291 
rect 198 291 201 294 
rect 198 294 201 297 
rect 198 297 201 300 
rect 198 300 201 303 
rect 198 303 201 306 
rect 198 306 201 309 
rect 198 309 201 312 
rect 198 312 201 315 
rect 198 315 201 318 
rect 198 318 201 321 
rect 198 321 201 324 
rect 198 324 201 327 
rect 198 327 201 330 
rect 198 330 201 333 
rect 198 333 201 336 
rect 198 336 201 339 
rect 198 339 201 342 
rect 198 342 201 345 
rect 198 345 201 348 
rect 198 348 201 351 
rect 198 351 201 354 
rect 198 354 201 357 
rect 198 357 201 360 
rect 198 360 201 363 
rect 198 363 201 366 
rect 198 366 201 369 
rect 198 369 201 372 
rect 198 372 201 375 
rect 198 375 201 378 
rect 198 378 201 381 
rect 198 381 201 384 
rect 198 384 201 387 
rect 198 387 201 390 
rect 198 390 201 393 
rect 198 393 201 396 
rect 198 396 201 399 
rect 198 399 201 402 
rect 198 402 201 405 
rect 198 405 201 408 
rect 198 408 201 411 
rect 198 411 201 414 
rect 198 414 201 417 
rect 198 417 201 420 
rect 198 420 201 423 
rect 198 423 201 426 
rect 198 426 201 429 
rect 198 429 201 432 
rect 198 432 201 435 
rect 198 435 201 438 
rect 198 438 201 441 
rect 198 441 201 444 
rect 198 444 201 447 
rect 198 447 201 450 
rect 198 450 201 453 
rect 198 453 201 456 
rect 198 456 201 459 
rect 198 459 201 462 
rect 198 462 201 465 
rect 198 465 201 468 
rect 198 468 201 471 
rect 198 471 201 474 
rect 198 474 201 477 
rect 198 477 201 480 
rect 198 480 201 483 
rect 198 483 201 486 
rect 198 486 201 489 
rect 198 489 201 492 
rect 198 492 201 495 
rect 198 495 201 498 
rect 198 498 201 501 
rect 198 501 201 504 
rect 198 504 201 507 
rect 198 507 201 510 
rect 201 0 204 3 
rect 201 3 204 6 
rect 201 6 204 9 
rect 201 9 204 12 
rect 201 12 204 15 
rect 201 15 204 18 
rect 201 18 204 21 
rect 201 21 204 24 
rect 201 24 204 27 
rect 201 27 204 30 
rect 201 30 204 33 
rect 201 33 204 36 
rect 201 36 204 39 
rect 201 39 204 42 
rect 201 42 204 45 
rect 201 45 204 48 
rect 201 48 204 51 
rect 201 51 204 54 
rect 201 54 204 57 
rect 201 57 204 60 
rect 201 60 204 63 
rect 201 63 204 66 
rect 201 66 204 69 
rect 201 69 204 72 
rect 201 72 204 75 
rect 201 75 204 78 
rect 201 78 204 81 
rect 201 81 204 84 
rect 201 84 204 87 
rect 201 87 204 90 
rect 201 90 204 93 
rect 201 93 204 96 
rect 201 96 204 99 
rect 201 99 204 102 
rect 201 102 204 105 
rect 201 105 204 108 
rect 201 108 204 111 
rect 201 111 204 114 
rect 201 114 204 117 
rect 201 117 204 120 
rect 201 120 204 123 
rect 201 123 204 126 
rect 201 126 204 129 
rect 201 129 204 132 
rect 201 132 204 135 
rect 201 135 204 138 
rect 201 138 204 141 
rect 201 141 204 144 
rect 201 144 204 147 
rect 201 147 204 150 
rect 201 150 204 153 
rect 201 153 204 156 
rect 201 156 204 159 
rect 201 159 204 162 
rect 201 162 204 165 
rect 201 165 204 168 
rect 201 168 204 171 
rect 201 171 204 174 
rect 201 174 204 177 
rect 201 177 204 180 
rect 201 180 204 183 
rect 201 183 204 186 
rect 201 186 204 189 
rect 201 189 204 192 
rect 201 192 204 195 
rect 201 195 204 198 
rect 201 198 204 201 
rect 201 201 204 204 
rect 201 204 204 207 
rect 201 207 204 210 
rect 201 210 204 213 
rect 201 213 204 216 
rect 201 216 204 219 
rect 201 219 204 222 
rect 201 222 204 225 
rect 201 225 204 228 
rect 201 228 204 231 
rect 201 231 204 234 
rect 201 234 204 237 
rect 201 237 204 240 
rect 201 240 204 243 
rect 201 243 204 246 
rect 201 246 204 249 
rect 201 249 204 252 
rect 201 252 204 255 
rect 201 255 204 258 
rect 201 258 204 261 
rect 201 261 204 264 
rect 201 264 204 267 
rect 201 267 204 270 
rect 201 270 204 273 
rect 201 273 204 276 
rect 201 276 204 279 
rect 201 279 204 282 
rect 201 282 204 285 
rect 201 285 204 288 
rect 201 288 204 291 
rect 201 291 204 294 
rect 201 294 204 297 
rect 201 297 204 300 
rect 201 300 204 303 
rect 201 303 204 306 
rect 201 306 204 309 
rect 201 309 204 312 
rect 201 312 204 315 
rect 201 315 204 318 
rect 201 318 204 321 
rect 201 321 204 324 
rect 201 324 204 327 
rect 201 327 204 330 
rect 201 330 204 333 
rect 201 333 204 336 
rect 201 336 204 339 
rect 201 339 204 342 
rect 201 342 204 345 
rect 201 345 204 348 
rect 201 348 204 351 
rect 201 351 204 354 
rect 201 354 204 357 
rect 201 357 204 360 
rect 201 360 204 363 
rect 201 363 204 366 
rect 201 366 204 369 
rect 201 369 204 372 
rect 201 372 204 375 
rect 201 375 204 378 
rect 201 378 204 381 
rect 201 381 204 384 
rect 201 384 204 387 
rect 201 387 204 390 
rect 201 390 204 393 
rect 201 393 204 396 
rect 201 396 204 399 
rect 201 399 204 402 
rect 201 402 204 405 
rect 201 405 204 408 
rect 201 408 204 411 
rect 201 411 204 414 
rect 201 414 204 417 
rect 201 417 204 420 
rect 201 420 204 423 
rect 201 423 204 426 
rect 201 426 204 429 
rect 201 429 204 432 
rect 201 432 204 435 
rect 201 435 204 438 
rect 201 438 204 441 
rect 201 441 204 444 
rect 201 444 204 447 
rect 201 447 204 450 
rect 201 450 204 453 
rect 201 453 204 456 
rect 201 456 204 459 
rect 201 459 204 462 
rect 201 462 204 465 
rect 201 465 204 468 
rect 201 468 204 471 
rect 201 471 204 474 
rect 201 474 204 477 
rect 201 477 204 480 
rect 201 480 204 483 
rect 201 483 204 486 
rect 201 486 204 489 
rect 201 489 204 492 
rect 201 492 204 495 
rect 201 495 204 498 
rect 201 498 204 501 
rect 201 501 204 504 
rect 201 504 204 507 
rect 201 507 204 510 
rect 204 0 207 3 
rect 204 3 207 6 
rect 204 6 207 9 
rect 204 9 207 12 
rect 204 12 207 15 
rect 204 15 207 18 
rect 204 18 207 21 
rect 204 21 207 24 
rect 204 24 207 27 
rect 204 27 207 30 
rect 204 30 207 33 
rect 204 33 207 36 
rect 204 36 207 39 
rect 204 39 207 42 
rect 204 42 207 45 
rect 204 45 207 48 
rect 204 48 207 51 
rect 204 51 207 54 
rect 204 54 207 57 
rect 204 57 207 60 
rect 204 60 207 63 
rect 204 63 207 66 
rect 204 66 207 69 
rect 204 69 207 72 
rect 204 72 207 75 
rect 204 75 207 78 
rect 204 78 207 81 
rect 204 81 207 84 
rect 204 84 207 87 
rect 204 87 207 90 
rect 204 90 207 93 
rect 204 93 207 96 
rect 204 96 207 99 
rect 204 99 207 102 
rect 204 102 207 105 
rect 204 105 207 108 
rect 204 108 207 111 
rect 204 111 207 114 
rect 204 114 207 117 
rect 204 117 207 120 
rect 204 120 207 123 
rect 204 123 207 126 
rect 204 126 207 129 
rect 204 129 207 132 
rect 204 132 207 135 
rect 204 135 207 138 
rect 204 138 207 141 
rect 204 141 207 144 
rect 204 144 207 147 
rect 204 147 207 150 
rect 204 150 207 153 
rect 204 153 207 156 
rect 204 156 207 159 
rect 204 159 207 162 
rect 204 162 207 165 
rect 204 165 207 168 
rect 204 168 207 171 
rect 204 171 207 174 
rect 204 174 207 177 
rect 204 177 207 180 
rect 204 180 207 183 
rect 204 183 207 186 
rect 204 186 207 189 
rect 204 189 207 192 
rect 204 192 207 195 
rect 204 195 207 198 
rect 204 198 207 201 
rect 204 201 207 204 
rect 204 204 207 207 
rect 204 207 207 210 
rect 204 210 207 213 
rect 204 213 207 216 
rect 204 216 207 219 
rect 204 219 207 222 
rect 204 222 207 225 
rect 204 225 207 228 
rect 204 228 207 231 
rect 204 231 207 234 
rect 204 234 207 237 
rect 204 237 207 240 
rect 204 240 207 243 
rect 204 243 207 246 
rect 204 246 207 249 
rect 204 249 207 252 
rect 204 252 207 255 
rect 204 255 207 258 
rect 204 258 207 261 
rect 204 261 207 264 
rect 204 264 207 267 
rect 204 267 207 270 
rect 204 270 207 273 
rect 204 273 207 276 
rect 204 276 207 279 
rect 204 279 207 282 
rect 204 282 207 285 
rect 204 285 207 288 
rect 204 288 207 291 
rect 204 291 207 294 
rect 204 294 207 297 
rect 204 297 207 300 
rect 204 300 207 303 
rect 204 303 207 306 
rect 204 306 207 309 
rect 204 309 207 312 
rect 204 312 207 315 
rect 204 315 207 318 
rect 204 318 207 321 
rect 204 321 207 324 
rect 204 324 207 327 
rect 204 327 207 330 
rect 204 330 207 333 
rect 204 333 207 336 
rect 204 336 207 339 
rect 204 339 207 342 
rect 204 342 207 345 
rect 204 345 207 348 
rect 204 348 207 351 
rect 204 351 207 354 
rect 204 354 207 357 
rect 204 357 207 360 
rect 204 360 207 363 
rect 204 363 207 366 
rect 204 366 207 369 
rect 204 369 207 372 
rect 204 372 207 375 
rect 204 375 207 378 
rect 204 378 207 381 
rect 204 381 207 384 
rect 204 384 207 387 
rect 204 387 207 390 
rect 204 390 207 393 
rect 204 393 207 396 
rect 204 396 207 399 
rect 204 399 207 402 
rect 204 402 207 405 
rect 204 405 207 408 
rect 204 408 207 411 
rect 204 411 207 414 
rect 204 414 207 417 
rect 204 417 207 420 
rect 204 420 207 423 
rect 204 423 207 426 
rect 204 426 207 429 
rect 204 429 207 432 
rect 204 432 207 435 
rect 204 435 207 438 
rect 204 438 207 441 
rect 204 441 207 444 
rect 204 444 207 447 
rect 204 447 207 450 
rect 204 450 207 453 
rect 204 453 207 456 
rect 204 456 207 459 
rect 204 459 207 462 
rect 204 462 207 465 
rect 204 465 207 468 
rect 204 468 207 471 
rect 204 471 207 474 
rect 204 474 207 477 
rect 204 477 207 480 
rect 204 480 207 483 
rect 204 483 207 486 
rect 204 486 207 489 
rect 204 489 207 492 
rect 204 492 207 495 
rect 204 495 207 498 
rect 204 498 207 501 
rect 204 501 207 504 
rect 204 504 207 507 
rect 204 507 207 510 
rect 207 0 210 3 
rect 207 3 210 6 
rect 207 6 210 9 
rect 207 9 210 12 
rect 207 12 210 15 
rect 207 15 210 18 
rect 207 18 210 21 
rect 207 21 210 24 
rect 207 24 210 27 
rect 207 27 210 30 
rect 207 30 210 33 
rect 207 33 210 36 
rect 207 36 210 39 
rect 207 39 210 42 
rect 207 42 210 45 
rect 207 45 210 48 
rect 207 48 210 51 
rect 207 51 210 54 
rect 207 54 210 57 
rect 207 57 210 60 
rect 207 60 210 63 
rect 207 63 210 66 
rect 207 66 210 69 
rect 207 69 210 72 
rect 207 72 210 75 
rect 207 75 210 78 
rect 207 78 210 81 
rect 207 81 210 84 
rect 207 84 210 87 
rect 207 87 210 90 
rect 207 90 210 93 
rect 207 93 210 96 
rect 207 96 210 99 
rect 207 99 210 102 
rect 207 102 210 105 
rect 207 105 210 108 
rect 207 108 210 111 
rect 207 111 210 114 
rect 207 114 210 117 
rect 207 117 210 120 
rect 207 120 210 123 
rect 207 123 210 126 
rect 207 126 210 129 
rect 207 129 210 132 
rect 207 132 210 135 
rect 207 135 210 138 
rect 207 138 210 141 
rect 207 141 210 144 
rect 207 144 210 147 
rect 207 147 210 150 
rect 207 150 210 153 
rect 207 153 210 156 
rect 207 156 210 159 
rect 207 159 210 162 
rect 207 162 210 165 
rect 207 165 210 168 
rect 207 168 210 171 
rect 207 171 210 174 
rect 207 174 210 177 
rect 207 177 210 180 
rect 207 180 210 183 
rect 207 183 210 186 
rect 207 186 210 189 
rect 207 189 210 192 
rect 207 192 210 195 
rect 207 195 210 198 
rect 207 198 210 201 
rect 207 201 210 204 
rect 207 204 210 207 
rect 207 207 210 210 
rect 207 210 210 213 
rect 207 213 210 216 
rect 207 216 210 219 
rect 207 219 210 222 
rect 207 222 210 225 
rect 207 225 210 228 
rect 207 228 210 231 
rect 207 231 210 234 
rect 207 234 210 237 
rect 207 237 210 240 
rect 207 240 210 243 
rect 207 243 210 246 
rect 207 246 210 249 
rect 207 249 210 252 
rect 207 252 210 255 
rect 207 255 210 258 
rect 207 258 210 261 
rect 207 261 210 264 
rect 207 264 210 267 
rect 207 267 210 270 
rect 207 270 210 273 
rect 207 273 210 276 
rect 207 276 210 279 
rect 207 279 210 282 
rect 207 282 210 285 
rect 207 285 210 288 
rect 207 288 210 291 
rect 207 291 210 294 
rect 207 294 210 297 
rect 207 297 210 300 
rect 207 300 210 303 
rect 207 303 210 306 
rect 207 306 210 309 
rect 207 309 210 312 
rect 207 312 210 315 
rect 207 315 210 318 
rect 207 318 210 321 
rect 207 321 210 324 
rect 207 324 210 327 
rect 207 327 210 330 
rect 207 330 210 333 
rect 207 333 210 336 
rect 207 336 210 339 
rect 207 339 210 342 
rect 207 342 210 345 
rect 207 345 210 348 
rect 207 348 210 351 
rect 207 351 210 354 
rect 207 354 210 357 
rect 207 357 210 360 
rect 207 360 210 363 
rect 207 363 210 366 
rect 207 366 210 369 
rect 207 369 210 372 
rect 207 372 210 375 
rect 207 375 210 378 
rect 207 378 210 381 
rect 207 381 210 384 
rect 207 384 210 387 
rect 207 387 210 390 
rect 207 390 210 393 
rect 207 393 210 396 
rect 207 396 210 399 
rect 207 399 210 402 
rect 207 402 210 405 
rect 207 405 210 408 
rect 207 408 210 411 
rect 207 411 210 414 
rect 207 414 210 417 
rect 207 417 210 420 
rect 207 420 210 423 
rect 207 423 210 426 
rect 207 426 210 429 
rect 207 429 210 432 
rect 207 432 210 435 
rect 207 435 210 438 
rect 207 438 210 441 
rect 207 441 210 444 
rect 207 444 210 447 
rect 207 447 210 450 
rect 207 450 210 453 
rect 207 453 210 456 
rect 207 456 210 459 
rect 207 459 210 462 
rect 207 462 210 465 
rect 207 465 210 468 
rect 207 468 210 471 
rect 207 471 210 474 
rect 207 474 210 477 
rect 207 477 210 480 
rect 207 480 210 483 
rect 207 483 210 486 
rect 207 486 210 489 
rect 207 489 210 492 
rect 207 492 210 495 
rect 207 495 210 498 
rect 207 498 210 501 
rect 207 501 210 504 
rect 207 504 210 507 
rect 207 507 210 510 
rect 210 0 213 3 
rect 210 3 213 6 
rect 210 6 213 9 
rect 210 9 213 12 
rect 210 12 213 15 
rect 210 15 213 18 
rect 210 18 213 21 
rect 210 21 213 24 
rect 210 24 213 27 
rect 210 27 213 30 
rect 210 30 213 33 
rect 210 33 213 36 
rect 210 36 213 39 
rect 210 39 213 42 
rect 210 42 213 45 
rect 210 45 213 48 
rect 210 48 213 51 
rect 210 51 213 54 
rect 210 54 213 57 
rect 210 57 213 60 
rect 210 60 213 63 
rect 210 63 213 66 
rect 210 66 213 69 
rect 210 69 213 72 
rect 210 72 213 75 
rect 210 75 213 78 
rect 210 78 213 81 
rect 210 81 213 84 
rect 210 84 213 87 
rect 210 87 213 90 
rect 210 90 213 93 
rect 210 93 213 96 
rect 210 96 213 99 
rect 210 99 213 102 
rect 210 102 213 105 
rect 210 105 213 108 
rect 210 108 213 111 
rect 210 111 213 114 
rect 210 114 213 117 
rect 210 117 213 120 
rect 210 120 213 123 
rect 210 123 213 126 
rect 210 126 213 129 
rect 210 129 213 132 
rect 210 132 213 135 
rect 210 135 213 138 
rect 210 138 213 141 
rect 210 141 213 144 
rect 210 144 213 147 
rect 210 147 213 150 
rect 210 150 213 153 
rect 210 153 213 156 
rect 210 156 213 159 
rect 210 159 213 162 
rect 210 162 213 165 
rect 210 165 213 168 
rect 210 168 213 171 
rect 210 171 213 174 
rect 210 174 213 177 
rect 210 177 213 180 
rect 210 180 213 183 
rect 210 183 213 186 
rect 210 186 213 189 
rect 210 189 213 192 
rect 210 192 213 195 
rect 210 195 213 198 
rect 210 198 213 201 
rect 210 201 213 204 
rect 210 204 213 207 
rect 210 207 213 210 
rect 210 210 213 213 
rect 210 213 213 216 
rect 210 216 213 219 
rect 210 219 213 222 
rect 210 222 213 225 
rect 210 225 213 228 
rect 210 228 213 231 
rect 210 231 213 234 
rect 210 234 213 237 
rect 210 237 213 240 
rect 210 240 213 243 
rect 210 243 213 246 
rect 210 246 213 249 
rect 210 249 213 252 
rect 210 252 213 255 
rect 210 255 213 258 
rect 210 258 213 261 
rect 210 261 213 264 
rect 210 264 213 267 
rect 210 267 213 270 
rect 210 270 213 273 
rect 210 273 213 276 
rect 210 276 213 279 
rect 210 279 213 282 
rect 210 282 213 285 
rect 210 285 213 288 
rect 210 288 213 291 
rect 210 291 213 294 
rect 210 294 213 297 
rect 210 297 213 300 
rect 210 300 213 303 
rect 210 303 213 306 
rect 210 306 213 309 
rect 210 309 213 312 
rect 210 312 213 315 
rect 210 315 213 318 
rect 210 318 213 321 
rect 210 321 213 324 
rect 210 324 213 327 
rect 210 327 213 330 
rect 210 330 213 333 
rect 210 333 213 336 
rect 210 336 213 339 
rect 210 339 213 342 
rect 210 342 213 345 
rect 210 345 213 348 
rect 210 348 213 351 
rect 210 351 213 354 
rect 210 354 213 357 
rect 210 357 213 360 
rect 210 360 213 363 
rect 210 363 213 366 
rect 210 366 213 369 
rect 210 369 213 372 
rect 210 372 213 375 
rect 210 375 213 378 
rect 210 378 213 381 
rect 210 381 213 384 
rect 210 384 213 387 
rect 210 387 213 390 
rect 210 390 213 393 
rect 210 393 213 396 
rect 210 396 213 399 
rect 210 399 213 402 
rect 210 402 213 405 
rect 210 405 213 408 
rect 210 408 213 411 
rect 210 411 213 414 
rect 210 414 213 417 
rect 210 417 213 420 
rect 210 420 213 423 
rect 210 423 213 426 
rect 210 426 213 429 
rect 210 429 213 432 
rect 210 432 213 435 
rect 210 435 213 438 
rect 210 438 213 441 
rect 210 441 213 444 
rect 210 444 213 447 
rect 210 447 213 450 
rect 210 450 213 453 
rect 210 453 213 456 
rect 210 456 213 459 
rect 210 459 213 462 
rect 210 462 213 465 
rect 210 465 213 468 
rect 210 468 213 471 
rect 210 471 213 474 
rect 210 474 213 477 
rect 210 477 213 480 
rect 210 480 213 483 
rect 210 483 213 486 
rect 210 486 213 489 
rect 210 489 213 492 
rect 210 492 213 495 
rect 210 495 213 498 
rect 210 498 213 501 
rect 210 501 213 504 
rect 210 504 213 507 
rect 210 507 213 510 
rect 213 0 216 3 
rect 213 3 216 6 
rect 213 6 216 9 
rect 213 9 216 12 
rect 213 12 216 15 
rect 213 15 216 18 
rect 213 18 216 21 
rect 213 21 216 24 
rect 213 24 216 27 
rect 213 27 216 30 
rect 213 30 216 33 
rect 213 33 216 36 
rect 213 36 216 39 
rect 213 39 216 42 
rect 213 42 216 45 
rect 213 45 216 48 
rect 213 48 216 51 
rect 213 51 216 54 
rect 213 54 216 57 
rect 213 57 216 60 
rect 213 60 216 63 
rect 213 63 216 66 
rect 213 66 216 69 
rect 213 69 216 72 
rect 213 72 216 75 
rect 213 75 216 78 
rect 213 78 216 81 
rect 213 81 216 84 
rect 213 84 216 87 
rect 213 87 216 90 
rect 213 90 216 93 
rect 213 93 216 96 
rect 213 96 216 99 
rect 213 99 216 102 
rect 213 102 216 105 
rect 213 105 216 108 
rect 213 108 216 111 
rect 213 111 216 114 
rect 213 114 216 117 
rect 213 117 216 120 
rect 213 120 216 123 
rect 213 123 216 126 
rect 213 126 216 129 
rect 213 129 216 132 
rect 213 132 216 135 
rect 213 135 216 138 
rect 213 138 216 141 
rect 213 141 216 144 
rect 213 144 216 147 
rect 213 147 216 150 
rect 213 150 216 153 
rect 213 153 216 156 
rect 213 156 216 159 
rect 213 159 216 162 
rect 213 162 216 165 
rect 213 165 216 168 
rect 213 168 216 171 
rect 213 171 216 174 
rect 213 174 216 177 
rect 213 177 216 180 
rect 213 180 216 183 
rect 213 183 216 186 
rect 213 186 216 189 
rect 213 189 216 192 
rect 213 192 216 195 
rect 213 195 216 198 
rect 213 198 216 201 
rect 213 201 216 204 
rect 213 204 216 207 
rect 213 207 216 210 
rect 213 210 216 213 
rect 213 213 216 216 
rect 213 216 216 219 
rect 213 219 216 222 
rect 213 222 216 225 
rect 213 225 216 228 
rect 213 228 216 231 
rect 213 231 216 234 
rect 213 234 216 237 
rect 213 237 216 240 
rect 213 240 216 243 
rect 213 243 216 246 
rect 213 246 216 249 
rect 213 249 216 252 
rect 213 252 216 255 
rect 213 255 216 258 
rect 213 258 216 261 
rect 213 261 216 264 
rect 213 264 216 267 
rect 213 267 216 270 
rect 213 270 216 273 
rect 213 273 216 276 
rect 213 276 216 279 
rect 213 279 216 282 
rect 213 282 216 285 
rect 213 285 216 288 
rect 213 288 216 291 
rect 213 291 216 294 
rect 213 294 216 297 
rect 213 297 216 300 
rect 213 300 216 303 
rect 213 303 216 306 
rect 213 306 216 309 
rect 213 309 216 312 
rect 213 312 216 315 
rect 213 315 216 318 
rect 213 318 216 321 
rect 213 321 216 324 
rect 213 324 216 327 
rect 213 327 216 330 
rect 213 330 216 333 
rect 213 333 216 336 
rect 213 336 216 339 
rect 213 339 216 342 
rect 213 342 216 345 
rect 213 345 216 348 
rect 213 348 216 351 
rect 213 351 216 354 
rect 213 354 216 357 
rect 213 357 216 360 
rect 213 360 216 363 
rect 213 363 216 366 
rect 213 366 216 369 
rect 213 369 216 372 
rect 213 372 216 375 
rect 213 375 216 378 
rect 213 378 216 381 
rect 213 381 216 384 
rect 213 384 216 387 
rect 213 387 216 390 
rect 213 390 216 393 
rect 213 393 216 396 
rect 213 396 216 399 
rect 213 399 216 402 
rect 213 402 216 405 
rect 213 405 216 408 
rect 213 408 216 411 
rect 213 411 216 414 
rect 213 414 216 417 
rect 213 417 216 420 
rect 213 420 216 423 
rect 213 423 216 426 
rect 213 426 216 429 
rect 213 429 216 432 
rect 213 432 216 435 
rect 213 435 216 438 
rect 213 438 216 441 
rect 213 441 216 444 
rect 213 444 216 447 
rect 213 447 216 450 
rect 213 450 216 453 
rect 213 453 216 456 
rect 213 456 216 459 
rect 213 459 216 462 
rect 213 462 216 465 
rect 213 465 216 468 
rect 213 468 216 471 
rect 213 471 216 474 
rect 213 474 216 477 
rect 213 477 216 480 
rect 213 480 216 483 
rect 213 483 216 486 
rect 213 486 216 489 
rect 213 489 216 492 
rect 213 492 216 495 
rect 213 495 216 498 
rect 213 498 216 501 
rect 213 501 216 504 
rect 213 504 216 507 
rect 213 507 216 510 
rect 216 0 219 3 
rect 216 3 219 6 
rect 216 6 219 9 
rect 216 9 219 12 
rect 216 12 219 15 
rect 216 15 219 18 
rect 216 18 219 21 
rect 216 21 219 24 
rect 216 24 219 27 
rect 216 27 219 30 
rect 216 30 219 33 
rect 216 33 219 36 
rect 216 36 219 39 
rect 216 39 219 42 
rect 216 42 219 45 
rect 216 45 219 48 
rect 216 48 219 51 
rect 216 51 219 54 
rect 216 54 219 57 
rect 216 57 219 60 
rect 216 60 219 63 
rect 216 63 219 66 
rect 216 66 219 69 
rect 216 69 219 72 
rect 216 72 219 75 
rect 216 75 219 78 
rect 216 78 219 81 
rect 216 81 219 84 
rect 216 84 219 87 
rect 216 87 219 90 
rect 216 90 219 93 
rect 216 93 219 96 
rect 216 96 219 99 
rect 216 99 219 102 
rect 216 102 219 105 
rect 216 105 219 108 
rect 216 108 219 111 
rect 216 111 219 114 
rect 216 114 219 117 
rect 216 117 219 120 
rect 216 120 219 123 
rect 216 123 219 126 
rect 216 126 219 129 
rect 216 129 219 132 
rect 216 132 219 135 
rect 216 135 219 138 
rect 216 138 219 141 
rect 216 141 219 144 
rect 216 144 219 147 
rect 216 147 219 150 
rect 216 150 219 153 
rect 216 153 219 156 
rect 216 156 219 159 
rect 216 159 219 162 
rect 216 162 219 165 
rect 216 165 219 168 
rect 216 168 219 171 
rect 216 171 219 174 
rect 216 174 219 177 
rect 216 177 219 180 
rect 216 180 219 183 
rect 216 183 219 186 
rect 216 186 219 189 
rect 216 189 219 192 
rect 216 192 219 195 
rect 216 195 219 198 
rect 216 198 219 201 
rect 216 201 219 204 
rect 216 204 219 207 
rect 216 207 219 210 
rect 216 210 219 213 
rect 216 213 219 216 
rect 216 216 219 219 
rect 216 219 219 222 
rect 216 222 219 225 
rect 216 225 219 228 
rect 216 228 219 231 
rect 216 231 219 234 
rect 216 234 219 237 
rect 216 237 219 240 
rect 216 240 219 243 
rect 216 243 219 246 
rect 216 246 219 249 
rect 216 249 219 252 
rect 216 252 219 255 
rect 216 255 219 258 
rect 216 258 219 261 
rect 216 261 219 264 
rect 216 264 219 267 
rect 216 267 219 270 
rect 216 270 219 273 
rect 216 273 219 276 
rect 216 276 219 279 
rect 216 279 219 282 
rect 216 282 219 285 
rect 216 285 219 288 
rect 216 288 219 291 
rect 216 291 219 294 
rect 216 294 219 297 
rect 216 297 219 300 
rect 216 300 219 303 
rect 216 303 219 306 
rect 216 306 219 309 
rect 216 309 219 312 
rect 216 312 219 315 
rect 216 315 219 318 
rect 216 318 219 321 
rect 216 321 219 324 
rect 216 324 219 327 
rect 216 327 219 330 
rect 216 330 219 333 
rect 216 333 219 336 
rect 216 336 219 339 
rect 216 339 219 342 
rect 216 342 219 345 
rect 216 345 219 348 
rect 216 348 219 351 
rect 216 351 219 354 
rect 216 354 219 357 
rect 216 357 219 360 
rect 216 360 219 363 
rect 216 363 219 366 
rect 216 366 219 369 
rect 216 369 219 372 
rect 216 372 219 375 
rect 216 375 219 378 
rect 216 378 219 381 
rect 216 381 219 384 
rect 216 384 219 387 
rect 216 387 219 390 
rect 216 390 219 393 
rect 216 393 219 396 
rect 216 396 219 399 
rect 216 399 219 402 
rect 216 402 219 405 
rect 216 405 219 408 
rect 216 408 219 411 
rect 216 411 219 414 
rect 216 414 219 417 
rect 216 417 219 420 
rect 216 420 219 423 
rect 216 423 219 426 
rect 216 426 219 429 
rect 216 429 219 432 
rect 216 432 219 435 
rect 216 435 219 438 
rect 216 438 219 441 
rect 216 441 219 444 
rect 216 444 219 447 
rect 216 447 219 450 
rect 216 450 219 453 
rect 216 453 219 456 
rect 216 456 219 459 
rect 216 459 219 462 
rect 216 462 219 465 
rect 216 465 219 468 
rect 216 468 219 471 
rect 216 471 219 474 
rect 216 474 219 477 
rect 216 477 219 480 
rect 216 480 219 483 
rect 216 483 219 486 
rect 216 486 219 489 
rect 216 489 219 492 
rect 216 492 219 495 
rect 216 495 219 498 
rect 216 498 219 501 
rect 216 501 219 504 
rect 216 504 219 507 
rect 216 507 219 510 
rect 219 0 222 3 
rect 219 3 222 6 
rect 219 6 222 9 
rect 219 9 222 12 
rect 219 12 222 15 
rect 219 15 222 18 
rect 219 18 222 21 
rect 219 21 222 24 
rect 219 24 222 27 
rect 219 27 222 30 
rect 219 30 222 33 
rect 219 33 222 36 
rect 219 36 222 39 
rect 219 39 222 42 
rect 219 42 222 45 
rect 219 45 222 48 
rect 219 48 222 51 
rect 219 51 222 54 
rect 219 54 222 57 
rect 219 57 222 60 
rect 219 60 222 63 
rect 219 63 222 66 
rect 219 66 222 69 
rect 219 69 222 72 
rect 219 72 222 75 
rect 219 75 222 78 
rect 219 78 222 81 
rect 219 81 222 84 
rect 219 84 222 87 
rect 219 87 222 90 
rect 219 90 222 93 
rect 219 93 222 96 
rect 219 96 222 99 
rect 219 99 222 102 
rect 219 102 222 105 
rect 219 105 222 108 
rect 219 108 222 111 
rect 219 111 222 114 
rect 219 114 222 117 
rect 219 117 222 120 
rect 219 120 222 123 
rect 219 123 222 126 
rect 219 126 222 129 
rect 219 129 222 132 
rect 219 132 222 135 
rect 219 135 222 138 
rect 219 138 222 141 
rect 219 141 222 144 
rect 219 144 222 147 
rect 219 147 222 150 
rect 219 150 222 153 
rect 219 153 222 156 
rect 219 156 222 159 
rect 219 159 222 162 
rect 219 162 222 165 
rect 219 165 222 168 
rect 219 168 222 171 
rect 219 171 222 174 
rect 219 174 222 177 
rect 219 177 222 180 
rect 219 180 222 183 
rect 219 183 222 186 
rect 219 186 222 189 
rect 219 189 222 192 
rect 219 192 222 195 
rect 219 195 222 198 
rect 219 198 222 201 
rect 219 201 222 204 
rect 219 204 222 207 
rect 219 207 222 210 
rect 219 210 222 213 
rect 219 213 222 216 
rect 219 216 222 219 
rect 219 219 222 222 
rect 219 222 222 225 
rect 219 225 222 228 
rect 219 228 222 231 
rect 219 231 222 234 
rect 219 234 222 237 
rect 219 237 222 240 
rect 219 240 222 243 
rect 219 243 222 246 
rect 219 246 222 249 
rect 219 249 222 252 
rect 219 252 222 255 
rect 219 255 222 258 
rect 219 258 222 261 
rect 219 261 222 264 
rect 219 264 222 267 
rect 219 267 222 270 
rect 219 270 222 273 
rect 219 273 222 276 
rect 219 276 222 279 
rect 219 279 222 282 
rect 219 282 222 285 
rect 219 285 222 288 
rect 219 288 222 291 
rect 219 291 222 294 
rect 219 294 222 297 
rect 219 297 222 300 
rect 219 300 222 303 
rect 219 303 222 306 
rect 219 306 222 309 
rect 219 309 222 312 
rect 219 312 222 315 
rect 219 315 222 318 
rect 219 318 222 321 
rect 219 321 222 324 
rect 219 324 222 327 
rect 219 327 222 330 
rect 219 330 222 333 
rect 219 333 222 336 
rect 219 336 222 339 
rect 219 339 222 342 
rect 219 342 222 345 
rect 219 345 222 348 
rect 219 348 222 351 
rect 219 351 222 354 
rect 219 354 222 357 
rect 219 357 222 360 
rect 219 360 222 363 
rect 219 363 222 366 
rect 219 366 222 369 
rect 219 369 222 372 
rect 219 372 222 375 
rect 219 375 222 378 
rect 219 378 222 381 
rect 219 381 222 384 
rect 219 384 222 387 
rect 219 387 222 390 
rect 219 390 222 393 
rect 219 393 222 396 
rect 219 396 222 399 
rect 219 399 222 402 
rect 219 402 222 405 
rect 219 405 222 408 
rect 219 408 222 411 
rect 219 411 222 414 
rect 219 414 222 417 
rect 219 417 222 420 
rect 219 420 222 423 
rect 219 423 222 426 
rect 219 426 222 429 
rect 219 429 222 432 
rect 219 432 222 435 
rect 219 435 222 438 
rect 219 438 222 441 
rect 219 441 222 444 
rect 219 444 222 447 
rect 219 447 222 450 
rect 219 450 222 453 
rect 219 453 222 456 
rect 219 456 222 459 
rect 219 459 222 462 
rect 219 462 222 465 
rect 219 465 222 468 
rect 219 468 222 471 
rect 219 471 222 474 
rect 219 474 222 477 
rect 219 477 222 480 
rect 219 480 222 483 
rect 219 483 222 486 
rect 219 486 222 489 
rect 219 489 222 492 
rect 219 492 222 495 
rect 219 495 222 498 
rect 219 498 222 501 
rect 219 501 222 504 
rect 219 504 222 507 
rect 219 507 222 510 
rect 222 0 225 3 
rect 222 3 225 6 
rect 222 6 225 9 
rect 222 9 225 12 
rect 222 12 225 15 
rect 222 15 225 18 
rect 222 18 225 21 
rect 222 21 225 24 
rect 222 24 225 27 
rect 222 27 225 30 
rect 222 30 225 33 
rect 222 33 225 36 
rect 222 36 225 39 
rect 222 39 225 42 
rect 222 42 225 45 
rect 222 45 225 48 
rect 222 48 225 51 
rect 222 51 225 54 
rect 222 54 225 57 
rect 222 57 225 60 
rect 222 60 225 63 
rect 222 63 225 66 
rect 222 66 225 69 
rect 222 69 225 72 
rect 222 72 225 75 
rect 222 75 225 78 
rect 222 78 225 81 
rect 222 81 225 84 
rect 222 84 225 87 
rect 222 87 225 90 
rect 222 90 225 93 
rect 222 93 225 96 
rect 222 96 225 99 
rect 222 99 225 102 
rect 222 102 225 105 
rect 222 105 225 108 
rect 222 108 225 111 
rect 222 111 225 114 
rect 222 114 225 117 
rect 222 117 225 120 
rect 222 120 225 123 
rect 222 123 225 126 
rect 222 126 225 129 
rect 222 129 225 132 
rect 222 132 225 135 
rect 222 135 225 138 
rect 222 138 225 141 
rect 222 141 225 144 
rect 222 144 225 147 
rect 222 147 225 150 
rect 222 150 225 153 
rect 222 153 225 156 
rect 222 156 225 159 
rect 222 159 225 162 
rect 222 162 225 165 
rect 222 165 225 168 
rect 222 168 225 171 
rect 222 171 225 174 
rect 222 174 225 177 
rect 222 177 225 180 
rect 222 180 225 183 
rect 222 183 225 186 
rect 222 186 225 189 
rect 222 189 225 192 
rect 222 192 225 195 
rect 222 195 225 198 
rect 222 198 225 201 
rect 222 201 225 204 
rect 222 204 225 207 
rect 222 207 225 210 
rect 222 210 225 213 
rect 222 213 225 216 
rect 222 216 225 219 
rect 222 219 225 222 
rect 222 222 225 225 
rect 222 225 225 228 
rect 222 228 225 231 
rect 222 231 225 234 
rect 222 237 225 240 
rect 222 240 225 243 
rect 222 243 225 246 
rect 222 246 225 249 
rect 222 249 225 252 
rect 222 252 225 255 
rect 222 255 225 258 
rect 222 258 225 261 
rect 222 261 225 264 
rect 222 264 225 267 
rect 222 267 225 270 
rect 222 270 225 273 
rect 222 273 225 276 
rect 222 276 225 279 
rect 222 279 225 282 
rect 222 285 225 288 
rect 222 288 225 291 
rect 222 291 225 294 
rect 222 294 225 297 
rect 222 297 225 300 
rect 222 300 225 303 
rect 222 303 225 306 
rect 222 306 225 309 
rect 222 309 225 312 
rect 222 312 225 315 
rect 222 315 225 318 
rect 222 318 225 321 
rect 222 321 225 324 
rect 222 324 225 327 
rect 222 327 225 330 
rect 222 330 225 333 
rect 222 333 225 336 
rect 222 336 225 339 
rect 222 339 225 342 
rect 222 342 225 345 
rect 222 345 225 348 
rect 222 348 225 351 
rect 222 351 225 354 
rect 222 354 225 357 
rect 222 357 225 360 
rect 222 360 225 363 
rect 222 363 225 366 
rect 222 366 225 369 
rect 222 369 225 372 
rect 222 372 225 375 
rect 222 375 225 378 
rect 222 378 225 381 
rect 222 381 225 384 
rect 222 384 225 387 
rect 222 387 225 390 
rect 222 390 225 393 
rect 222 393 225 396 
rect 222 396 225 399 
rect 222 399 225 402 
rect 222 402 225 405 
rect 222 405 225 408 
rect 222 408 225 411 
rect 222 411 225 414 
rect 222 414 225 417 
rect 222 417 225 420 
rect 222 420 225 423 
rect 222 423 225 426 
rect 222 426 225 429 
rect 222 429 225 432 
rect 222 432 225 435 
rect 222 435 225 438 
rect 222 438 225 441 
rect 222 441 225 444 
rect 222 444 225 447 
rect 222 447 225 450 
rect 222 450 225 453 
rect 222 453 225 456 
rect 222 456 225 459 
rect 222 459 225 462 
rect 222 462 225 465 
rect 222 465 225 468 
rect 222 468 225 471 
rect 222 471 225 474 
rect 222 474 225 477 
rect 222 477 225 480 
rect 222 480 225 483 
rect 222 483 225 486 
rect 222 486 225 489 
rect 222 489 225 492 
rect 222 492 225 495 
rect 222 495 225 498 
rect 222 498 225 501 
rect 222 501 225 504 
rect 222 504 225 507 
rect 222 507 225 510 
rect 225 0 228 3 
rect 225 3 228 6 
rect 225 6 228 9 
rect 225 9 228 12 
rect 225 12 228 15 
rect 225 15 228 18 
rect 225 18 228 21 
rect 225 21 228 24 
rect 225 24 228 27 
rect 225 27 228 30 
rect 225 30 228 33 
rect 225 33 228 36 
rect 225 36 228 39 
rect 225 39 228 42 
rect 225 42 228 45 
rect 225 45 228 48 
rect 225 48 228 51 
rect 225 51 228 54 
rect 225 54 228 57 
rect 225 57 228 60 
rect 225 60 228 63 
rect 225 63 228 66 
rect 225 66 228 69 
rect 225 69 228 72 
rect 225 72 228 75 
rect 225 75 228 78 
rect 225 78 228 81 
rect 225 81 228 84 
rect 225 84 228 87 
rect 225 87 228 90 
rect 225 90 228 93 
rect 225 93 228 96 
rect 225 96 228 99 
rect 225 99 228 102 
rect 225 102 228 105 
rect 225 105 228 108 
rect 225 108 228 111 
rect 225 111 228 114 
rect 225 114 228 117 
rect 225 117 228 120 
rect 225 120 228 123 
rect 225 123 228 126 
rect 225 126 228 129 
rect 225 129 228 132 
rect 225 132 228 135 
rect 225 135 228 138 
rect 225 138 228 141 
rect 225 141 228 144 
rect 225 144 228 147 
rect 225 147 228 150 
rect 225 150 228 153 
rect 225 153 228 156 
rect 225 156 228 159 
rect 225 159 228 162 
rect 225 162 228 165 
rect 225 165 228 168 
rect 225 168 228 171 
rect 225 171 228 174 
rect 225 174 228 177 
rect 225 177 228 180 
rect 225 180 228 183 
rect 225 183 228 186 
rect 225 186 228 189 
rect 225 189 228 192 
rect 225 192 228 195 
rect 225 195 228 198 
rect 225 198 228 201 
rect 225 201 228 204 
rect 225 204 228 207 
rect 225 207 228 210 
rect 225 210 228 213 
rect 225 213 228 216 
rect 225 216 228 219 
rect 225 219 228 222 
rect 225 222 228 225 
rect 225 225 228 228 
rect 225 228 228 231 
rect 225 231 228 234 
rect 225 234 228 237 
rect 225 237 228 240 
rect 225 240 228 243 
rect 225 243 228 246 
rect 225 246 228 249 
rect 225 249 228 252 
rect 225 252 228 255 
rect 225 255 228 258 
rect 225 258 228 261 
rect 225 261 228 264 
rect 225 264 228 267 
rect 225 267 228 270 
rect 225 270 228 273 
rect 225 273 228 276 
rect 225 276 228 279 
rect 225 279 228 282 
rect 225 282 228 285 
rect 225 285 228 288 
rect 225 288 228 291 
rect 225 291 228 294 
rect 225 294 228 297 
rect 225 297 228 300 
rect 225 300 228 303 
rect 225 303 228 306 
rect 225 306 228 309 
rect 225 309 228 312 
rect 225 312 228 315 
rect 225 315 228 318 
rect 225 318 228 321 
rect 225 321 228 324 
rect 225 324 228 327 
rect 225 327 228 330 
rect 225 330 228 333 
rect 225 333 228 336 
rect 225 336 228 339 
rect 225 339 228 342 
rect 225 342 228 345 
rect 225 345 228 348 
rect 225 348 228 351 
rect 225 351 228 354 
rect 225 354 228 357 
rect 225 357 228 360 
rect 225 360 228 363 
rect 225 363 228 366 
rect 225 366 228 369 
rect 225 369 228 372 
rect 225 372 228 375 
rect 225 375 228 378 
rect 225 378 228 381 
rect 225 381 228 384 
rect 225 384 228 387 
rect 225 387 228 390 
rect 225 390 228 393 
rect 225 393 228 396 
rect 225 396 228 399 
rect 225 399 228 402 
rect 225 402 228 405 
rect 225 405 228 408 
rect 225 408 228 411 
rect 225 411 228 414 
rect 225 414 228 417 
rect 225 417 228 420 
rect 225 420 228 423 
rect 225 423 228 426 
rect 225 426 228 429 
rect 225 429 228 432 
rect 225 432 228 435 
rect 225 435 228 438 
rect 225 438 228 441 
rect 225 441 228 444 
rect 225 444 228 447 
rect 225 447 228 450 
rect 225 450 228 453 
rect 225 453 228 456 
rect 225 456 228 459 
rect 225 459 228 462 
rect 225 462 228 465 
rect 225 465 228 468 
rect 225 468 228 471 
rect 225 471 228 474 
rect 225 474 228 477 
rect 225 477 228 480 
rect 225 480 228 483 
rect 225 483 228 486 
rect 225 486 228 489 
rect 225 489 228 492 
rect 225 492 228 495 
rect 225 495 228 498 
rect 225 498 228 501 
rect 225 501 228 504 
rect 225 504 228 507 
rect 225 507 228 510 
rect 228 0 231 3 
rect 228 3 231 6 
rect 228 6 231 9 
rect 228 9 231 12 
rect 228 12 231 15 
rect 228 15 231 18 
rect 228 18 231 21 
rect 228 21 231 24 
rect 228 24 231 27 
rect 228 27 231 30 
rect 228 30 231 33 
rect 228 33 231 36 
rect 228 36 231 39 
rect 228 39 231 42 
rect 228 42 231 45 
rect 228 45 231 48 
rect 228 48 231 51 
rect 228 51 231 54 
rect 228 54 231 57 
rect 228 57 231 60 
rect 228 60 231 63 
rect 228 63 231 66 
rect 228 66 231 69 
rect 228 69 231 72 
rect 228 72 231 75 
rect 228 75 231 78 
rect 228 78 231 81 
rect 228 81 231 84 
rect 228 84 231 87 
rect 228 87 231 90 
rect 228 90 231 93 
rect 228 93 231 96 
rect 228 96 231 99 
rect 228 99 231 102 
rect 228 102 231 105 
rect 228 105 231 108 
rect 228 108 231 111 
rect 228 111 231 114 
rect 228 114 231 117 
rect 228 117 231 120 
rect 228 120 231 123 
rect 228 123 231 126 
rect 228 126 231 129 
rect 228 129 231 132 
rect 228 132 231 135 
rect 228 135 231 138 
rect 228 138 231 141 
rect 228 141 231 144 
rect 228 144 231 147 
rect 228 147 231 150 
rect 228 150 231 153 
rect 228 153 231 156 
rect 228 156 231 159 
rect 228 159 231 162 
rect 228 162 231 165 
rect 228 165 231 168 
rect 228 168 231 171 
rect 228 171 231 174 
rect 228 174 231 177 
rect 228 177 231 180 
rect 228 180 231 183 
rect 228 183 231 186 
rect 228 186 231 189 
rect 228 189 231 192 
rect 228 192 231 195 
rect 228 195 231 198 
rect 228 198 231 201 
rect 228 201 231 204 
rect 228 204 231 207 
rect 228 207 231 210 
rect 228 210 231 213 
rect 228 213 231 216 
rect 228 216 231 219 
rect 228 219 231 222 
rect 228 222 231 225 
rect 228 225 231 228 
rect 228 228 231 231 
rect 228 231 231 234 
rect 228 234 231 237 
rect 228 237 231 240 
rect 228 240 231 243 
rect 228 243 231 246 
rect 228 246 231 249 
rect 228 249 231 252 
rect 228 252 231 255 
rect 228 255 231 258 
rect 228 258 231 261 
rect 228 261 231 264 
rect 228 264 231 267 
rect 228 267 231 270 
rect 228 270 231 273 
rect 228 273 231 276 
rect 228 276 231 279 
rect 228 279 231 282 
rect 228 282 231 285 
rect 228 285 231 288 
rect 228 288 231 291 
rect 228 291 231 294 
rect 228 294 231 297 
rect 228 297 231 300 
rect 228 300 231 303 
rect 228 303 231 306 
rect 228 306 231 309 
rect 228 309 231 312 
rect 228 312 231 315 
rect 228 315 231 318 
rect 228 318 231 321 
rect 228 321 231 324 
rect 228 324 231 327 
rect 228 327 231 330 
rect 228 330 231 333 
rect 228 333 231 336 
rect 228 336 231 339 
rect 228 339 231 342 
rect 228 342 231 345 
rect 228 345 231 348 
rect 228 348 231 351 
rect 228 351 231 354 
rect 228 354 231 357 
rect 228 357 231 360 
rect 228 360 231 363 
rect 228 363 231 366 
rect 228 366 231 369 
rect 228 369 231 372 
rect 228 372 231 375 
rect 228 375 231 378 
rect 228 378 231 381 
rect 228 381 231 384 
rect 228 384 231 387 
rect 228 387 231 390 
rect 228 390 231 393 
rect 228 393 231 396 
rect 228 396 231 399 
rect 228 399 231 402 
rect 228 402 231 405 
rect 228 405 231 408 
rect 228 408 231 411 
rect 228 411 231 414 
rect 228 414 231 417 
rect 228 417 231 420 
rect 228 420 231 423 
rect 228 423 231 426 
rect 228 426 231 429 
rect 228 429 231 432 
rect 228 432 231 435 
rect 228 435 231 438 
rect 228 438 231 441 
rect 228 441 231 444 
rect 228 444 231 447 
rect 228 447 231 450 
rect 228 450 231 453 
rect 228 453 231 456 
rect 228 456 231 459 
rect 228 459 231 462 
rect 228 462 231 465 
rect 228 465 231 468 
rect 228 468 231 471 
rect 228 471 231 474 
rect 228 474 231 477 
rect 228 477 231 480 
rect 228 480 231 483 
rect 228 483 231 486 
rect 228 486 231 489 
rect 228 489 231 492 
rect 228 492 231 495 
rect 228 495 231 498 
rect 228 498 231 501 
rect 228 501 231 504 
rect 228 504 231 507 
rect 228 507 231 510 
rect 231 0 234 3 
rect 231 3 234 6 
rect 231 6 234 9 
rect 231 9 234 12 
rect 231 12 234 15 
rect 231 15 234 18 
rect 231 18 234 21 
rect 231 21 234 24 
rect 231 24 234 27 
rect 231 27 234 30 
rect 231 30 234 33 
rect 231 33 234 36 
rect 231 36 234 39 
rect 231 39 234 42 
rect 231 42 234 45 
rect 231 45 234 48 
rect 231 48 234 51 
rect 231 51 234 54 
rect 231 54 234 57 
rect 231 57 234 60 
rect 231 60 234 63 
rect 231 63 234 66 
rect 231 66 234 69 
rect 231 69 234 72 
rect 231 72 234 75 
rect 231 75 234 78 
rect 231 78 234 81 
rect 231 81 234 84 
rect 231 84 234 87 
rect 231 87 234 90 
rect 231 90 234 93 
rect 231 93 234 96 
rect 231 96 234 99 
rect 231 99 234 102 
rect 231 102 234 105 
rect 231 105 234 108 
rect 231 108 234 111 
rect 231 111 234 114 
rect 231 114 234 117 
rect 231 117 234 120 
rect 231 120 234 123 
rect 231 123 234 126 
rect 231 126 234 129 
rect 231 129 234 132 
rect 231 132 234 135 
rect 231 135 234 138 
rect 231 138 234 141 
rect 231 141 234 144 
rect 231 144 234 147 
rect 231 147 234 150 
rect 231 150 234 153 
rect 231 153 234 156 
rect 231 156 234 159 
rect 231 159 234 162 
rect 231 162 234 165 
rect 231 165 234 168 
rect 231 168 234 171 
rect 231 171 234 174 
rect 231 174 234 177 
rect 231 177 234 180 
rect 231 180 234 183 
rect 231 183 234 186 
rect 231 186 234 189 
rect 231 189 234 192 
rect 231 192 234 195 
rect 231 195 234 198 
rect 231 198 234 201 
rect 231 201 234 204 
rect 231 204 234 207 
rect 231 207 234 210 
rect 231 210 234 213 
rect 231 213 234 216 
rect 231 216 234 219 
rect 231 219 234 222 
rect 231 222 234 225 
rect 231 225 234 228 
rect 231 228 234 231 
rect 231 231 234 234 
rect 231 234 234 237 
rect 231 237 234 240 
rect 231 240 234 243 
rect 231 243 234 246 
rect 231 246 234 249 
rect 231 249 234 252 
rect 231 252 234 255 
rect 231 255 234 258 
rect 231 258 234 261 
rect 231 261 234 264 
rect 231 264 234 267 
rect 231 267 234 270 
rect 231 270 234 273 
rect 231 273 234 276 
rect 231 276 234 279 
rect 231 279 234 282 
rect 231 282 234 285 
rect 231 285 234 288 
rect 231 288 234 291 
rect 231 291 234 294 
rect 231 294 234 297 
rect 231 297 234 300 
rect 231 300 234 303 
rect 231 303 234 306 
rect 231 306 234 309 
rect 231 309 234 312 
rect 231 312 234 315 
rect 231 315 234 318 
rect 231 318 234 321 
rect 231 321 234 324 
rect 231 324 234 327 
rect 231 327 234 330 
rect 231 330 234 333 
rect 231 333 234 336 
rect 231 336 234 339 
rect 231 339 234 342 
rect 231 342 234 345 
rect 231 345 234 348 
rect 231 348 234 351 
rect 231 351 234 354 
rect 231 354 234 357 
rect 231 357 234 360 
rect 231 360 234 363 
rect 231 363 234 366 
rect 231 366 234 369 
rect 231 369 234 372 
rect 231 372 234 375 
rect 231 375 234 378 
rect 231 378 234 381 
rect 231 381 234 384 
rect 231 384 234 387 
rect 231 387 234 390 
rect 231 390 234 393 
rect 231 393 234 396 
rect 231 396 234 399 
rect 231 399 234 402 
rect 231 402 234 405 
rect 231 405 234 408 
rect 231 408 234 411 
rect 231 411 234 414 
rect 231 414 234 417 
rect 231 417 234 420 
rect 231 420 234 423 
rect 231 423 234 426 
rect 231 426 234 429 
rect 231 429 234 432 
rect 231 432 234 435 
rect 231 435 234 438 
rect 231 438 234 441 
rect 231 441 234 444 
rect 231 444 234 447 
rect 231 447 234 450 
rect 231 450 234 453 
rect 231 453 234 456 
rect 231 456 234 459 
rect 231 459 234 462 
rect 231 462 234 465 
rect 231 465 234 468 
rect 231 468 234 471 
rect 231 471 234 474 
rect 231 474 234 477 
rect 231 477 234 480 
rect 231 480 234 483 
rect 231 483 234 486 
rect 231 486 234 489 
rect 231 489 234 492 
rect 231 492 234 495 
rect 231 495 234 498 
rect 231 498 234 501 
rect 231 501 234 504 
rect 231 504 234 507 
rect 231 507 234 510 
rect 234 0 237 3 
rect 234 3 237 6 
rect 234 6 237 9 
rect 234 9 237 12 
rect 234 12 237 15 
rect 234 15 237 18 
rect 234 18 237 21 
rect 234 21 237 24 
rect 234 24 237 27 
rect 234 27 237 30 
rect 234 30 237 33 
rect 234 33 237 36 
rect 234 36 237 39 
rect 234 39 237 42 
rect 234 42 237 45 
rect 234 45 237 48 
rect 234 48 237 51 
rect 234 51 237 54 
rect 234 54 237 57 
rect 234 57 237 60 
rect 234 60 237 63 
rect 234 63 237 66 
rect 234 66 237 69 
rect 234 69 237 72 
rect 234 72 237 75 
rect 234 75 237 78 
rect 234 78 237 81 
rect 234 81 237 84 
rect 234 84 237 87 
rect 234 87 237 90 
rect 234 90 237 93 
rect 234 93 237 96 
rect 234 96 237 99 
rect 234 99 237 102 
rect 234 102 237 105 
rect 234 105 237 108 
rect 234 108 237 111 
rect 234 111 237 114 
rect 234 114 237 117 
rect 234 117 237 120 
rect 234 120 237 123 
rect 234 123 237 126 
rect 234 126 237 129 
rect 234 129 237 132 
rect 234 132 237 135 
rect 234 135 237 138 
rect 234 138 237 141 
rect 234 141 237 144 
rect 234 144 237 147 
rect 234 147 237 150 
rect 234 150 237 153 
rect 234 153 237 156 
rect 234 156 237 159 
rect 234 159 237 162 
rect 234 162 237 165 
rect 234 165 237 168 
rect 234 168 237 171 
rect 234 171 237 174 
rect 234 174 237 177 
rect 234 177 237 180 
rect 234 180 237 183 
rect 234 183 237 186 
rect 234 186 237 189 
rect 234 189 237 192 
rect 234 192 237 195 
rect 234 195 237 198 
rect 234 198 237 201 
rect 234 201 237 204 
rect 234 204 237 207 
rect 234 207 237 210 
rect 234 210 237 213 
rect 234 213 237 216 
rect 234 216 237 219 
rect 234 219 237 222 
rect 234 222 237 225 
rect 234 225 237 228 
rect 234 228 237 231 
rect 234 231 237 234 
rect 234 234 237 237 
rect 234 237 237 240 
rect 234 240 237 243 
rect 234 243 237 246 
rect 234 246 237 249 
rect 234 249 237 252 
rect 234 252 237 255 
rect 234 255 237 258 
rect 234 258 237 261 
rect 234 261 237 264 
rect 234 264 237 267 
rect 234 267 237 270 
rect 234 270 237 273 
rect 234 273 237 276 
rect 234 276 237 279 
rect 234 279 237 282 
rect 234 282 237 285 
rect 234 285 237 288 
rect 234 288 237 291 
rect 234 291 237 294 
rect 234 294 237 297 
rect 234 297 237 300 
rect 234 300 237 303 
rect 234 303 237 306 
rect 234 306 237 309 
rect 234 309 237 312 
rect 234 312 237 315 
rect 234 315 237 318 
rect 234 318 237 321 
rect 234 321 237 324 
rect 234 324 237 327 
rect 234 327 237 330 
rect 234 330 237 333 
rect 234 333 237 336 
rect 234 336 237 339 
rect 234 339 237 342 
rect 234 342 237 345 
rect 234 345 237 348 
rect 234 348 237 351 
rect 234 351 237 354 
rect 234 354 237 357 
rect 234 357 237 360 
rect 234 360 237 363 
rect 234 363 237 366 
rect 234 366 237 369 
rect 234 369 237 372 
rect 234 372 237 375 
rect 234 375 237 378 
rect 234 378 237 381 
rect 234 381 237 384 
rect 234 384 237 387 
rect 234 387 237 390 
rect 234 390 237 393 
rect 234 393 237 396 
rect 234 396 237 399 
rect 234 399 237 402 
rect 234 402 237 405 
rect 234 405 237 408 
rect 234 408 237 411 
rect 234 411 237 414 
rect 234 414 237 417 
rect 234 417 237 420 
rect 234 420 237 423 
rect 234 423 237 426 
rect 234 426 237 429 
rect 234 429 237 432 
rect 234 432 237 435 
rect 234 435 237 438 
rect 234 438 237 441 
rect 234 441 237 444 
rect 234 444 237 447 
rect 234 447 237 450 
rect 234 450 237 453 
rect 234 453 237 456 
rect 234 456 237 459 
rect 234 459 237 462 
rect 234 462 237 465 
rect 234 465 237 468 
rect 234 468 237 471 
rect 234 471 237 474 
rect 234 474 237 477 
rect 234 477 237 480 
rect 234 480 237 483 
rect 234 483 237 486 
rect 234 486 237 489 
rect 234 489 237 492 
rect 234 492 237 495 
rect 234 495 237 498 
rect 234 498 237 501 
rect 234 501 237 504 
rect 234 504 237 507 
rect 234 507 237 510 
rect 237 0 240 3 
rect 237 3 240 6 
rect 237 6 240 9 
rect 237 9 240 12 
rect 237 12 240 15 
rect 237 15 240 18 
rect 237 18 240 21 
rect 237 21 240 24 
rect 237 24 240 27 
rect 237 27 240 30 
rect 237 30 240 33 
rect 237 33 240 36 
rect 237 36 240 39 
rect 237 39 240 42 
rect 237 42 240 45 
rect 237 45 240 48 
rect 237 48 240 51 
rect 237 51 240 54 
rect 237 54 240 57 
rect 237 57 240 60 
rect 237 60 240 63 
rect 237 63 240 66 
rect 237 66 240 69 
rect 237 69 240 72 
rect 237 72 240 75 
rect 237 75 240 78 
rect 237 78 240 81 
rect 237 81 240 84 
rect 237 84 240 87 
rect 237 87 240 90 
rect 237 90 240 93 
rect 237 93 240 96 
rect 237 96 240 99 
rect 237 99 240 102 
rect 237 102 240 105 
rect 237 105 240 108 
rect 237 108 240 111 
rect 237 111 240 114 
rect 237 114 240 117 
rect 237 117 240 120 
rect 237 120 240 123 
rect 237 123 240 126 
rect 237 126 240 129 
rect 237 129 240 132 
rect 237 132 240 135 
rect 237 135 240 138 
rect 237 138 240 141 
rect 237 141 240 144 
rect 237 144 240 147 
rect 237 147 240 150 
rect 237 150 240 153 
rect 237 153 240 156 
rect 237 156 240 159 
rect 237 159 240 162 
rect 237 162 240 165 
rect 237 165 240 168 
rect 237 168 240 171 
rect 237 171 240 174 
rect 237 174 240 177 
rect 237 177 240 180 
rect 237 180 240 183 
rect 237 183 240 186 
rect 237 186 240 189 
rect 237 189 240 192 
rect 237 192 240 195 
rect 237 195 240 198 
rect 237 198 240 201 
rect 237 201 240 204 
rect 237 204 240 207 
rect 237 207 240 210 
rect 237 210 240 213 
rect 237 213 240 216 
rect 237 216 240 219 
rect 237 219 240 222 
rect 237 222 240 225 
rect 237 228 240 231 
rect 237 231 240 234 
rect 237 234 240 237 
rect 237 237 240 240 
rect 237 240 240 243 
rect 237 243 240 246 
rect 237 246 240 249 
rect 237 249 240 252 
rect 237 252 240 255 
rect 237 255 240 258 
rect 237 258 240 261 
rect 237 261 240 264 
rect 237 264 240 267 
rect 237 267 240 270 
rect 237 270 240 273 
rect 237 273 240 276 
rect 237 276 240 279 
rect 237 279 240 282 
rect 237 282 240 285 
rect 237 285 240 288 
rect 237 288 240 291 
rect 237 291 240 294 
rect 237 294 240 297 
rect 237 297 240 300 
rect 237 300 240 303 
rect 237 303 240 306 
rect 237 306 240 309 
rect 237 309 240 312 
rect 237 312 240 315 
rect 237 315 240 318 
rect 237 318 240 321 
rect 237 321 240 324 
rect 237 324 240 327 
rect 237 327 240 330 
rect 237 333 240 336 
rect 237 336 240 339 
rect 237 339 240 342 
rect 237 342 240 345 
rect 237 345 240 348 
rect 237 348 240 351 
rect 237 351 240 354 
rect 237 354 240 357 
rect 237 357 240 360 
rect 237 360 240 363 
rect 237 363 240 366 
rect 237 366 240 369 
rect 237 369 240 372 
rect 237 372 240 375 
rect 237 375 240 378 
rect 237 378 240 381 
rect 237 381 240 384 
rect 237 384 240 387 
rect 237 387 240 390 
rect 237 390 240 393 
rect 237 393 240 396 
rect 237 396 240 399 
rect 237 399 240 402 
rect 237 402 240 405 
rect 237 405 240 408 
rect 237 408 240 411 
rect 237 411 240 414 
rect 237 414 240 417 
rect 237 417 240 420 
rect 237 420 240 423 
rect 237 423 240 426 
rect 237 426 240 429 
rect 237 429 240 432 
rect 237 432 240 435 
rect 237 435 240 438 
rect 237 438 240 441 
rect 237 441 240 444 
rect 237 444 240 447 
rect 237 447 240 450 
rect 237 450 240 453 
rect 237 453 240 456 
rect 237 456 240 459 
rect 237 459 240 462 
rect 237 462 240 465 
rect 237 465 240 468 
rect 237 468 240 471 
rect 237 471 240 474 
rect 237 474 240 477 
rect 237 477 240 480 
rect 237 480 240 483 
rect 237 483 240 486 
rect 237 486 240 489 
rect 237 489 240 492 
rect 237 492 240 495 
rect 237 495 240 498 
rect 237 498 240 501 
rect 237 501 240 504 
rect 237 504 240 507 
rect 237 507 240 510 
rect 240 0 243 3 
rect 240 3 243 6 
rect 240 6 243 9 
rect 240 9 243 12 
rect 240 12 243 15 
rect 240 15 243 18 
rect 240 18 243 21 
rect 240 21 243 24 
rect 240 24 243 27 
rect 240 27 243 30 
rect 240 30 243 33 
rect 240 33 243 36 
rect 240 36 243 39 
rect 240 39 243 42 
rect 240 42 243 45 
rect 240 45 243 48 
rect 240 48 243 51 
rect 240 51 243 54 
rect 240 54 243 57 
rect 240 57 243 60 
rect 240 60 243 63 
rect 240 63 243 66 
rect 240 66 243 69 
rect 240 69 243 72 
rect 240 72 243 75 
rect 240 75 243 78 
rect 240 78 243 81 
rect 240 81 243 84 
rect 240 84 243 87 
rect 240 87 243 90 
rect 240 90 243 93 
rect 240 93 243 96 
rect 240 96 243 99 
rect 240 99 243 102 
rect 240 102 243 105 
rect 240 105 243 108 
rect 240 108 243 111 
rect 240 111 243 114 
rect 240 114 243 117 
rect 240 117 243 120 
rect 240 120 243 123 
rect 240 123 243 126 
rect 240 126 243 129 
rect 240 129 243 132 
rect 240 132 243 135 
rect 240 135 243 138 
rect 240 138 243 141 
rect 240 141 243 144 
rect 240 144 243 147 
rect 240 147 243 150 
rect 240 150 243 153 
rect 240 153 243 156 
rect 240 156 243 159 
rect 240 159 243 162 
rect 240 162 243 165 
rect 240 165 243 168 
rect 240 168 243 171 
rect 240 171 243 174 
rect 240 174 243 177 
rect 240 177 243 180 
rect 240 180 243 183 
rect 240 183 243 186 
rect 240 186 243 189 
rect 240 189 243 192 
rect 240 192 243 195 
rect 240 195 243 198 
rect 240 198 243 201 
rect 240 201 243 204 
rect 240 204 243 207 
rect 240 207 243 210 
rect 240 210 243 213 
rect 240 213 243 216 
rect 240 216 243 219 
rect 240 219 243 222 
rect 240 222 243 225 
rect 240 225 243 228 
rect 240 228 243 231 
rect 240 231 243 234 
rect 240 234 243 237 
rect 240 237 243 240 
rect 240 240 243 243 
rect 240 243 243 246 
rect 240 246 243 249 
rect 240 249 243 252 
rect 240 252 243 255 
rect 240 255 243 258 
rect 240 258 243 261 
rect 240 261 243 264 
rect 240 264 243 267 
rect 240 267 243 270 
rect 240 270 243 273 
rect 240 273 243 276 
rect 240 276 243 279 
rect 240 279 243 282 
rect 240 282 243 285 
rect 240 285 243 288 
rect 240 288 243 291 
rect 240 291 243 294 
rect 240 294 243 297 
rect 240 297 243 300 
rect 240 300 243 303 
rect 240 303 243 306 
rect 240 306 243 309 
rect 240 309 243 312 
rect 240 312 243 315 
rect 240 315 243 318 
rect 240 318 243 321 
rect 240 321 243 324 
rect 240 324 243 327 
rect 240 327 243 330 
rect 240 330 243 333 
rect 240 333 243 336 
rect 240 336 243 339 
rect 240 339 243 342 
rect 240 342 243 345 
rect 240 345 243 348 
rect 240 348 243 351 
rect 240 351 243 354 
rect 240 354 243 357 
rect 240 357 243 360 
rect 240 360 243 363 
rect 240 363 243 366 
rect 240 366 243 369 
rect 240 369 243 372 
rect 240 372 243 375 
rect 240 375 243 378 
rect 240 378 243 381 
rect 240 381 243 384 
rect 240 384 243 387 
rect 240 387 243 390 
rect 240 390 243 393 
rect 240 393 243 396 
rect 240 396 243 399 
rect 240 399 243 402 
rect 240 402 243 405 
rect 240 405 243 408 
rect 240 408 243 411 
rect 240 411 243 414 
rect 240 414 243 417 
rect 240 417 243 420 
rect 240 420 243 423 
rect 240 423 243 426 
rect 240 426 243 429 
rect 240 429 243 432 
rect 240 432 243 435 
rect 240 435 243 438 
rect 240 438 243 441 
rect 240 441 243 444 
rect 240 444 243 447 
rect 240 447 243 450 
rect 240 450 243 453 
rect 240 453 243 456 
rect 240 456 243 459 
rect 240 459 243 462 
rect 240 462 243 465 
rect 240 465 243 468 
rect 240 468 243 471 
rect 240 471 243 474 
rect 240 474 243 477 
rect 240 477 243 480 
rect 240 480 243 483 
rect 240 483 243 486 
rect 240 486 243 489 
rect 240 489 243 492 
rect 240 492 243 495 
rect 240 495 243 498 
rect 240 498 243 501 
rect 240 501 243 504 
rect 240 504 243 507 
rect 240 507 243 510 
rect 243 0 246 3 
rect 243 3 246 6 
rect 243 6 246 9 
rect 243 9 246 12 
rect 243 12 246 15 
rect 243 15 246 18 
rect 243 18 246 21 
rect 243 21 246 24 
rect 243 24 246 27 
rect 243 27 246 30 
rect 243 30 246 33 
rect 243 33 246 36 
rect 243 36 246 39 
rect 243 39 246 42 
rect 243 42 246 45 
rect 243 45 246 48 
rect 243 48 246 51 
rect 243 51 246 54 
rect 243 54 246 57 
rect 243 57 246 60 
rect 243 60 246 63 
rect 243 63 246 66 
rect 243 66 246 69 
rect 243 69 246 72 
rect 243 72 246 75 
rect 243 75 246 78 
rect 243 78 246 81 
rect 243 81 246 84 
rect 243 84 246 87 
rect 243 87 246 90 
rect 243 90 246 93 
rect 243 93 246 96 
rect 243 96 246 99 
rect 243 99 246 102 
rect 243 102 246 105 
rect 243 105 246 108 
rect 243 108 246 111 
rect 243 111 246 114 
rect 243 114 246 117 
rect 243 117 246 120 
rect 243 120 246 123 
rect 243 123 246 126 
rect 243 126 246 129 
rect 243 129 246 132 
rect 243 132 246 135 
rect 243 135 246 138 
rect 243 138 246 141 
rect 243 141 246 144 
rect 243 144 246 147 
rect 243 147 246 150 
rect 243 150 246 153 
rect 243 153 246 156 
rect 243 156 246 159 
rect 243 159 246 162 
rect 243 162 246 165 
rect 243 165 246 168 
rect 243 168 246 171 
rect 243 171 246 174 
rect 243 174 246 177 
rect 243 177 246 180 
rect 243 180 246 183 
rect 243 183 246 186 
rect 243 186 246 189 
rect 243 189 246 192 
rect 243 192 246 195 
rect 243 195 246 198 
rect 243 198 246 201 
rect 243 201 246 204 
rect 243 204 246 207 
rect 243 207 246 210 
rect 243 210 246 213 
rect 243 213 246 216 
rect 243 216 246 219 
rect 243 219 246 222 
rect 243 222 246 225 
rect 243 225 246 228 
rect 243 228 246 231 
rect 243 231 246 234 
rect 243 234 246 237 
rect 243 237 246 240 
rect 243 240 246 243 
rect 243 243 246 246 
rect 243 246 246 249 
rect 243 249 246 252 
rect 243 252 246 255 
rect 243 255 246 258 
rect 243 258 246 261 
rect 243 261 246 264 
rect 243 264 246 267 
rect 243 267 246 270 
rect 243 270 246 273 
rect 243 273 246 276 
rect 243 276 246 279 
rect 243 279 246 282 
rect 243 282 246 285 
rect 243 285 246 288 
rect 243 288 246 291 
rect 243 291 246 294 
rect 243 294 246 297 
rect 243 297 246 300 
rect 243 300 246 303 
rect 243 303 246 306 
rect 243 306 246 309 
rect 243 309 246 312 
rect 243 312 246 315 
rect 243 315 246 318 
rect 243 318 246 321 
rect 243 321 246 324 
rect 243 324 246 327 
rect 243 327 246 330 
rect 243 330 246 333 
rect 243 333 246 336 
rect 243 336 246 339 
rect 243 339 246 342 
rect 243 342 246 345 
rect 243 345 246 348 
rect 243 348 246 351 
rect 243 351 246 354 
rect 243 354 246 357 
rect 243 357 246 360 
rect 243 360 246 363 
rect 243 363 246 366 
rect 243 366 246 369 
rect 243 369 246 372 
rect 243 372 246 375 
rect 243 375 246 378 
rect 243 378 246 381 
rect 243 381 246 384 
rect 243 384 246 387 
rect 243 387 246 390 
rect 243 390 246 393 
rect 243 393 246 396 
rect 243 396 246 399 
rect 243 399 246 402 
rect 243 402 246 405 
rect 243 405 246 408 
rect 243 408 246 411 
rect 243 411 246 414 
rect 243 414 246 417 
rect 243 417 246 420 
rect 243 420 246 423 
rect 243 423 246 426 
rect 243 426 246 429 
rect 243 429 246 432 
rect 243 432 246 435 
rect 243 435 246 438 
rect 243 438 246 441 
rect 243 441 246 444 
rect 243 444 246 447 
rect 243 447 246 450 
rect 243 450 246 453 
rect 243 453 246 456 
rect 243 456 246 459 
rect 243 459 246 462 
rect 243 462 246 465 
rect 243 465 246 468 
rect 243 468 246 471 
rect 243 471 246 474 
rect 243 474 246 477 
rect 243 477 246 480 
rect 243 480 246 483 
rect 243 483 246 486 
rect 243 486 246 489 
rect 243 489 246 492 
rect 243 492 246 495 
rect 243 495 246 498 
rect 243 498 246 501 
rect 243 501 246 504 
rect 243 504 246 507 
rect 243 507 246 510 
rect 246 0 249 3 
rect 246 3 249 6 
rect 246 6 249 9 
rect 246 9 249 12 
rect 246 12 249 15 
rect 246 15 249 18 
rect 246 18 249 21 
rect 246 21 249 24 
rect 246 24 249 27 
rect 246 27 249 30 
rect 246 30 249 33 
rect 246 33 249 36 
rect 246 36 249 39 
rect 246 39 249 42 
rect 246 42 249 45 
rect 246 45 249 48 
rect 246 48 249 51 
rect 246 51 249 54 
rect 246 54 249 57 
rect 246 57 249 60 
rect 246 60 249 63 
rect 246 63 249 66 
rect 246 66 249 69 
rect 246 69 249 72 
rect 246 72 249 75 
rect 246 75 249 78 
rect 246 78 249 81 
rect 246 81 249 84 
rect 246 84 249 87 
rect 246 87 249 90 
rect 246 90 249 93 
rect 246 93 249 96 
rect 246 96 249 99 
rect 246 99 249 102 
rect 246 102 249 105 
rect 246 105 249 108 
rect 246 108 249 111 
rect 246 111 249 114 
rect 246 114 249 117 
rect 246 117 249 120 
rect 246 120 249 123 
rect 246 123 249 126 
rect 246 126 249 129 
rect 246 129 249 132 
rect 246 132 249 135 
rect 246 135 249 138 
rect 246 138 249 141 
rect 246 141 249 144 
rect 246 144 249 147 
rect 246 147 249 150 
rect 246 150 249 153 
rect 246 153 249 156 
rect 246 156 249 159 
rect 246 159 249 162 
rect 246 162 249 165 
rect 246 165 249 168 
rect 246 168 249 171 
rect 246 171 249 174 
rect 246 174 249 177 
rect 246 177 249 180 
rect 246 180 249 183 
rect 246 183 249 186 
rect 246 186 249 189 
rect 246 189 249 192 
rect 246 192 249 195 
rect 246 195 249 198 
rect 246 198 249 201 
rect 246 201 249 204 
rect 246 204 249 207 
rect 246 207 249 210 
rect 246 210 249 213 
rect 246 213 249 216 
rect 246 216 249 219 
rect 246 219 249 222 
rect 246 222 249 225 
rect 246 225 249 228 
rect 246 228 249 231 
rect 246 231 249 234 
rect 246 234 249 237 
rect 246 237 249 240 
rect 246 240 249 243 
rect 246 243 249 246 
rect 246 246 249 249 
rect 246 249 249 252 
rect 246 252 249 255 
rect 246 255 249 258 
rect 246 258 249 261 
rect 246 261 249 264 
rect 246 264 249 267 
rect 246 267 249 270 
rect 246 270 249 273 
rect 246 273 249 276 
rect 246 276 249 279 
rect 246 279 249 282 
rect 246 282 249 285 
rect 246 285 249 288 
rect 246 288 249 291 
rect 246 291 249 294 
rect 246 294 249 297 
rect 246 297 249 300 
rect 246 300 249 303 
rect 246 303 249 306 
rect 246 306 249 309 
rect 246 309 249 312 
rect 246 312 249 315 
rect 246 315 249 318 
rect 246 318 249 321 
rect 246 321 249 324 
rect 246 324 249 327 
rect 246 327 249 330 
rect 246 330 249 333 
rect 246 333 249 336 
rect 246 336 249 339 
rect 246 339 249 342 
rect 246 342 249 345 
rect 246 345 249 348 
rect 246 348 249 351 
rect 246 351 249 354 
rect 246 354 249 357 
rect 246 357 249 360 
rect 246 360 249 363 
rect 246 363 249 366 
rect 246 366 249 369 
rect 246 369 249 372 
rect 246 372 249 375 
rect 246 375 249 378 
rect 246 378 249 381 
rect 246 381 249 384 
rect 246 384 249 387 
rect 246 387 249 390 
rect 246 390 249 393 
rect 246 393 249 396 
rect 246 396 249 399 
rect 246 399 249 402 
rect 246 402 249 405 
rect 246 405 249 408 
rect 246 408 249 411 
rect 246 411 249 414 
rect 246 414 249 417 
rect 246 417 249 420 
rect 246 420 249 423 
rect 246 423 249 426 
rect 246 426 249 429 
rect 246 429 249 432 
rect 246 432 249 435 
rect 246 435 249 438 
rect 246 438 249 441 
rect 246 441 249 444 
rect 246 444 249 447 
rect 246 447 249 450 
rect 246 450 249 453 
rect 246 453 249 456 
rect 246 456 249 459 
rect 246 459 249 462 
rect 246 462 249 465 
rect 246 465 249 468 
rect 246 468 249 471 
rect 246 471 249 474 
rect 246 474 249 477 
rect 246 477 249 480 
rect 246 480 249 483 
rect 246 483 249 486 
rect 246 486 249 489 
rect 246 489 249 492 
rect 246 492 249 495 
rect 246 495 249 498 
rect 246 498 249 501 
rect 246 501 249 504 
rect 246 504 249 507 
rect 246 507 249 510 
rect 249 0 252 3 
rect 249 3 252 6 
rect 249 6 252 9 
rect 249 9 252 12 
rect 249 12 252 15 
rect 249 15 252 18 
rect 249 18 252 21 
rect 249 21 252 24 
rect 249 24 252 27 
rect 249 27 252 30 
rect 249 30 252 33 
rect 249 33 252 36 
rect 249 36 252 39 
rect 249 39 252 42 
rect 249 42 252 45 
rect 249 45 252 48 
rect 249 48 252 51 
rect 249 51 252 54 
rect 249 54 252 57 
rect 249 57 252 60 
rect 249 60 252 63 
rect 249 63 252 66 
rect 249 66 252 69 
rect 249 69 252 72 
rect 249 72 252 75 
rect 249 75 252 78 
rect 249 78 252 81 
rect 249 81 252 84 
rect 249 84 252 87 
rect 249 87 252 90 
rect 249 90 252 93 
rect 249 93 252 96 
rect 249 96 252 99 
rect 249 99 252 102 
rect 249 102 252 105 
rect 249 105 252 108 
rect 249 108 252 111 
rect 249 111 252 114 
rect 249 114 252 117 
rect 249 117 252 120 
rect 249 120 252 123 
rect 249 123 252 126 
rect 249 126 252 129 
rect 249 129 252 132 
rect 249 132 252 135 
rect 249 135 252 138 
rect 249 138 252 141 
rect 249 141 252 144 
rect 249 144 252 147 
rect 249 147 252 150 
rect 249 150 252 153 
rect 249 153 252 156 
rect 249 156 252 159 
rect 249 159 252 162 
rect 249 162 252 165 
rect 249 165 252 168 
rect 249 168 252 171 
rect 249 171 252 174 
rect 249 174 252 177 
rect 249 177 252 180 
rect 249 180 252 183 
rect 249 183 252 186 
rect 249 186 252 189 
rect 249 189 252 192 
rect 249 192 252 195 
rect 249 195 252 198 
rect 249 198 252 201 
rect 249 201 252 204 
rect 249 204 252 207 
rect 249 207 252 210 
rect 249 210 252 213 
rect 249 213 252 216 
rect 249 216 252 219 
rect 249 219 252 222 
rect 249 222 252 225 
rect 249 225 252 228 
rect 249 228 252 231 
rect 249 231 252 234 
rect 249 234 252 237 
rect 249 237 252 240 
rect 249 240 252 243 
rect 249 243 252 246 
rect 249 246 252 249 
rect 249 249 252 252 
rect 249 252 252 255 
rect 249 255 252 258 
rect 249 258 252 261 
rect 249 261 252 264 
rect 249 264 252 267 
rect 249 267 252 270 
rect 249 270 252 273 
rect 249 273 252 276 
rect 249 276 252 279 
rect 249 279 252 282 
rect 249 282 252 285 
rect 249 285 252 288 
rect 249 288 252 291 
rect 249 291 252 294 
rect 249 294 252 297 
rect 249 297 252 300 
rect 249 300 252 303 
rect 249 303 252 306 
rect 249 306 252 309 
rect 249 309 252 312 
rect 249 312 252 315 
rect 249 315 252 318 
rect 249 318 252 321 
rect 249 321 252 324 
rect 249 324 252 327 
rect 249 327 252 330 
rect 249 330 252 333 
rect 249 333 252 336 
rect 249 336 252 339 
rect 249 339 252 342 
rect 249 342 252 345 
rect 249 345 252 348 
rect 249 348 252 351 
rect 249 351 252 354 
rect 249 354 252 357 
rect 249 357 252 360 
rect 249 360 252 363 
rect 249 363 252 366 
rect 249 366 252 369 
rect 249 369 252 372 
rect 249 372 252 375 
rect 249 375 252 378 
rect 249 378 252 381 
rect 249 381 252 384 
rect 249 384 252 387 
rect 249 387 252 390 
rect 249 390 252 393 
rect 249 393 252 396 
rect 249 396 252 399 
rect 249 399 252 402 
rect 249 402 252 405 
rect 249 405 252 408 
rect 249 408 252 411 
rect 249 411 252 414 
rect 249 414 252 417 
rect 249 417 252 420 
rect 249 420 252 423 
rect 249 423 252 426 
rect 249 426 252 429 
rect 249 429 252 432 
rect 249 432 252 435 
rect 249 435 252 438 
rect 249 438 252 441 
rect 249 441 252 444 
rect 249 444 252 447 
rect 249 447 252 450 
rect 249 450 252 453 
rect 249 453 252 456 
rect 249 456 252 459 
rect 249 459 252 462 
rect 249 462 252 465 
rect 249 465 252 468 
rect 249 468 252 471 
rect 249 471 252 474 
rect 249 474 252 477 
rect 249 477 252 480 
rect 249 480 252 483 
rect 249 483 252 486 
rect 249 486 252 489 
rect 249 489 252 492 
rect 249 492 252 495 
rect 249 495 252 498 
rect 249 498 252 501 
rect 249 501 252 504 
rect 249 504 252 507 
rect 249 507 252 510 
rect 252 0 255 3 
rect 252 3 255 6 
rect 252 6 255 9 
rect 252 9 255 12 
rect 252 12 255 15 
rect 252 15 255 18 
rect 252 18 255 21 
rect 252 21 255 24 
rect 252 24 255 27 
rect 252 27 255 30 
rect 252 30 255 33 
rect 252 33 255 36 
rect 252 36 255 39 
rect 252 39 255 42 
rect 252 42 255 45 
rect 252 45 255 48 
rect 252 48 255 51 
rect 252 51 255 54 
rect 252 54 255 57 
rect 252 57 255 60 
rect 252 60 255 63 
rect 252 63 255 66 
rect 252 66 255 69 
rect 252 69 255 72 
rect 252 72 255 75 
rect 252 75 255 78 
rect 252 78 255 81 
rect 252 81 255 84 
rect 252 84 255 87 
rect 252 87 255 90 
rect 252 90 255 93 
rect 252 93 255 96 
rect 252 96 255 99 
rect 252 99 255 102 
rect 252 102 255 105 
rect 252 105 255 108 
rect 252 108 255 111 
rect 252 111 255 114 
rect 252 114 255 117 
rect 252 117 255 120 
rect 252 120 255 123 
rect 252 123 255 126 
rect 252 126 255 129 
rect 252 129 255 132 
rect 252 132 255 135 
rect 252 135 255 138 
rect 252 138 255 141 
rect 252 141 255 144 
rect 252 144 255 147 
rect 252 147 255 150 
rect 252 150 255 153 
rect 252 153 255 156 
rect 252 156 255 159 
rect 252 159 255 162 
rect 252 162 255 165 
rect 252 165 255 168 
rect 252 168 255 171 
rect 252 171 255 174 
rect 252 174 255 177 
rect 252 177 255 180 
rect 252 180 255 183 
rect 252 183 255 186 
rect 252 186 255 189 
rect 252 189 255 192 
rect 252 192 255 195 
rect 252 195 255 198 
rect 252 198 255 201 
rect 252 201 255 204 
rect 252 204 255 207 
rect 252 207 255 210 
rect 252 210 255 213 
rect 252 213 255 216 
rect 252 216 255 219 
rect 252 219 255 222 
rect 252 222 255 225 
rect 252 225 255 228 
rect 252 228 255 231 
rect 252 231 255 234 
rect 252 234 255 237 
rect 252 237 255 240 
rect 252 240 255 243 
rect 252 243 255 246 
rect 252 246 255 249 
rect 252 249 255 252 
rect 252 252 255 255 
rect 252 255 255 258 
rect 252 258 255 261 
rect 252 261 255 264 
rect 252 264 255 267 
rect 252 267 255 270 
rect 252 270 255 273 
rect 252 273 255 276 
rect 252 276 255 279 
rect 252 279 255 282 
rect 252 282 255 285 
rect 252 285 255 288 
rect 252 288 255 291 
rect 252 291 255 294 
rect 252 294 255 297 
rect 252 297 255 300 
rect 252 300 255 303 
rect 252 303 255 306 
rect 252 306 255 309 
rect 252 309 255 312 
rect 252 312 255 315 
rect 252 315 255 318 
rect 252 318 255 321 
rect 252 321 255 324 
rect 252 324 255 327 
rect 252 327 255 330 
rect 252 330 255 333 
rect 252 333 255 336 
rect 252 336 255 339 
rect 252 339 255 342 
rect 252 342 255 345 
rect 252 345 255 348 
rect 252 348 255 351 
rect 252 351 255 354 
rect 252 354 255 357 
rect 252 357 255 360 
rect 252 360 255 363 
rect 252 363 255 366 
rect 252 366 255 369 
rect 252 369 255 372 
rect 252 372 255 375 
rect 252 375 255 378 
rect 252 378 255 381 
rect 252 381 255 384 
rect 252 384 255 387 
rect 252 387 255 390 
rect 252 390 255 393 
rect 252 393 255 396 
rect 252 396 255 399 
rect 252 399 255 402 
rect 252 402 255 405 
rect 252 405 255 408 
rect 252 408 255 411 
rect 252 411 255 414 
rect 252 414 255 417 
rect 252 417 255 420 
rect 252 420 255 423 
rect 252 423 255 426 
rect 252 426 255 429 
rect 252 429 255 432 
rect 252 432 255 435 
rect 252 435 255 438 
rect 252 438 255 441 
rect 252 441 255 444 
rect 252 444 255 447 
rect 252 447 255 450 
rect 252 450 255 453 
rect 252 453 255 456 
rect 252 456 255 459 
rect 252 459 255 462 
rect 252 462 255 465 
rect 252 465 255 468 
rect 252 468 255 471 
rect 252 471 255 474 
rect 252 474 255 477 
rect 252 477 255 480 
rect 252 480 255 483 
rect 252 483 255 486 
rect 252 486 255 489 
rect 252 489 255 492 
rect 252 492 255 495 
rect 252 495 255 498 
rect 252 498 255 501 
rect 252 501 255 504 
rect 252 504 255 507 
rect 252 507 255 510 
rect 255 0 258 3 
rect 255 3 258 6 
rect 255 6 258 9 
rect 255 9 258 12 
rect 255 12 258 15 
rect 255 15 258 18 
rect 255 18 258 21 
rect 255 21 258 24 
rect 255 24 258 27 
rect 255 27 258 30 
rect 255 30 258 33 
rect 255 33 258 36 
rect 255 36 258 39 
rect 255 39 258 42 
rect 255 42 258 45 
rect 255 45 258 48 
rect 255 48 258 51 
rect 255 51 258 54 
rect 255 54 258 57 
rect 255 57 258 60 
rect 255 60 258 63 
rect 255 63 258 66 
rect 255 66 258 69 
rect 255 69 258 72 
rect 255 72 258 75 
rect 255 75 258 78 
rect 255 78 258 81 
rect 255 81 258 84 
rect 255 84 258 87 
rect 255 87 258 90 
rect 255 90 258 93 
rect 255 93 258 96 
rect 255 96 258 99 
rect 255 99 258 102 
rect 255 102 258 105 
rect 255 105 258 108 
rect 255 108 258 111 
rect 255 111 258 114 
rect 255 114 258 117 
rect 255 117 258 120 
rect 255 120 258 123 
rect 255 123 258 126 
rect 255 126 258 129 
rect 255 129 258 132 
rect 255 132 258 135 
rect 255 135 258 138 
rect 255 138 258 141 
rect 255 141 258 144 
rect 255 144 258 147 
rect 255 147 258 150 
rect 255 150 258 153 
rect 255 153 258 156 
rect 255 156 258 159 
rect 255 159 258 162 
rect 255 162 258 165 
rect 255 165 258 168 
rect 255 168 258 171 
rect 255 171 258 174 
rect 255 174 258 177 
rect 255 177 258 180 
rect 255 180 258 183 
rect 255 183 258 186 
rect 255 186 258 189 
rect 255 189 258 192 
rect 255 192 258 195 
rect 255 195 258 198 
rect 255 198 258 201 
rect 255 201 258 204 
rect 255 204 258 207 
rect 255 207 258 210 
rect 255 210 258 213 
rect 255 213 258 216 
rect 255 216 258 219 
rect 255 219 258 222 
rect 255 222 258 225 
rect 255 225 258 228 
rect 255 228 258 231 
rect 255 231 258 234 
rect 255 234 258 237 
rect 255 237 258 240 
rect 255 240 258 243 
rect 255 243 258 246 
rect 255 246 258 249 
rect 255 249 258 252 
rect 255 252 258 255 
rect 255 255 258 258 
rect 255 258 258 261 
rect 255 261 258 264 
rect 255 264 258 267 
rect 255 267 258 270 
rect 255 270 258 273 
rect 255 273 258 276 
rect 255 276 258 279 
rect 255 279 258 282 
rect 255 282 258 285 
rect 255 285 258 288 
rect 255 288 258 291 
rect 255 291 258 294 
rect 255 294 258 297 
rect 255 297 258 300 
rect 255 300 258 303 
rect 255 303 258 306 
rect 255 306 258 309 
rect 255 309 258 312 
rect 255 312 258 315 
rect 255 315 258 318 
rect 255 318 258 321 
rect 255 321 258 324 
rect 255 324 258 327 
rect 255 327 258 330 
rect 255 330 258 333 
rect 255 333 258 336 
rect 255 336 258 339 
rect 255 339 258 342 
rect 255 342 258 345 
rect 255 345 258 348 
rect 255 348 258 351 
rect 255 351 258 354 
rect 255 354 258 357 
rect 255 357 258 360 
rect 255 360 258 363 
rect 255 363 258 366 
rect 255 366 258 369 
rect 255 369 258 372 
rect 255 372 258 375 
rect 255 375 258 378 
rect 255 378 258 381 
rect 255 381 258 384 
rect 255 384 258 387 
rect 255 387 258 390 
rect 255 390 258 393 
rect 255 393 258 396 
rect 255 396 258 399 
rect 255 399 258 402 
rect 255 402 258 405 
rect 255 405 258 408 
rect 255 408 258 411 
rect 255 411 258 414 
rect 255 414 258 417 
rect 255 417 258 420 
rect 255 420 258 423 
rect 255 423 258 426 
rect 255 426 258 429 
rect 255 429 258 432 
rect 255 432 258 435 
rect 255 435 258 438 
rect 255 438 258 441 
rect 255 441 258 444 
rect 255 444 258 447 
rect 255 447 258 450 
rect 255 450 258 453 
rect 255 453 258 456 
rect 255 456 258 459 
rect 255 459 258 462 
rect 255 462 258 465 
rect 255 465 258 468 
rect 255 468 258 471 
rect 255 471 258 474 
rect 255 474 258 477 
rect 255 477 258 480 
rect 255 480 258 483 
rect 255 483 258 486 
rect 255 486 258 489 
rect 255 489 258 492 
rect 255 492 258 495 
rect 255 495 258 498 
rect 255 498 258 501 
rect 255 501 258 504 
rect 255 504 258 507 
rect 255 507 258 510 
rect 258 0 261 3 
rect 258 3 261 6 
rect 258 6 261 9 
rect 258 9 261 12 
rect 258 12 261 15 
rect 258 15 261 18 
rect 258 18 261 21 
rect 258 21 261 24 
rect 258 24 261 27 
rect 258 27 261 30 
rect 258 30 261 33 
rect 258 33 261 36 
rect 258 36 261 39 
rect 258 39 261 42 
rect 258 42 261 45 
rect 258 45 261 48 
rect 258 48 261 51 
rect 258 51 261 54 
rect 258 54 261 57 
rect 258 57 261 60 
rect 258 60 261 63 
rect 258 63 261 66 
rect 258 66 261 69 
rect 258 69 261 72 
rect 258 72 261 75 
rect 258 75 261 78 
rect 258 78 261 81 
rect 258 81 261 84 
rect 258 84 261 87 
rect 258 87 261 90 
rect 258 90 261 93 
rect 258 93 261 96 
rect 258 96 261 99 
rect 258 99 261 102 
rect 258 102 261 105 
rect 258 105 261 108 
rect 258 108 261 111 
rect 258 111 261 114 
rect 258 114 261 117 
rect 258 117 261 120 
rect 258 120 261 123 
rect 258 123 261 126 
rect 258 126 261 129 
rect 258 129 261 132 
rect 258 132 261 135 
rect 258 135 261 138 
rect 258 138 261 141 
rect 258 141 261 144 
rect 258 144 261 147 
rect 258 147 261 150 
rect 258 150 261 153 
rect 258 153 261 156 
rect 258 156 261 159 
rect 258 159 261 162 
rect 258 162 261 165 
rect 258 165 261 168 
rect 258 168 261 171 
rect 258 171 261 174 
rect 258 174 261 177 
rect 258 177 261 180 
rect 258 180 261 183 
rect 258 183 261 186 
rect 258 186 261 189 
rect 258 189 261 192 
rect 258 192 261 195 
rect 258 195 261 198 
rect 258 198 261 201 
rect 258 201 261 204 
rect 258 204 261 207 
rect 258 207 261 210 
rect 258 210 261 213 
rect 258 213 261 216 
rect 258 216 261 219 
rect 258 219 261 222 
rect 258 222 261 225 
rect 258 225 261 228 
rect 258 228 261 231 
rect 258 231 261 234 
rect 258 234 261 237 
rect 258 237 261 240 
rect 258 240 261 243 
rect 258 243 261 246 
rect 258 246 261 249 
rect 258 249 261 252 
rect 258 252 261 255 
rect 258 255 261 258 
rect 258 258 261 261 
rect 258 261 261 264 
rect 258 264 261 267 
rect 258 267 261 270 
rect 258 270 261 273 
rect 258 273 261 276 
rect 258 276 261 279 
rect 258 279 261 282 
rect 258 282 261 285 
rect 258 285 261 288 
rect 258 288 261 291 
rect 258 291 261 294 
rect 258 294 261 297 
rect 258 297 261 300 
rect 258 300 261 303 
rect 258 303 261 306 
rect 258 306 261 309 
rect 258 309 261 312 
rect 258 312 261 315 
rect 258 315 261 318 
rect 258 318 261 321 
rect 258 321 261 324 
rect 258 324 261 327 
rect 258 327 261 330 
rect 258 330 261 333 
rect 258 333 261 336 
rect 258 336 261 339 
rect 258 339 261 342 
rect 258 342 261 345 
rect 258 345 261 348 
rect 258 348 261 351 
rect 258 351 261 354 
rect 258 354 261 357 
rect 258 357 261 360 
rect 258 360 261 363 
rect 258 363 261 366 
rect 258 366 261 369 
rect 258 369 261 372 
rect 258 372 261 375 
rect 258 375 261 378 
rect 258 378 261 381 
rect 258 381 261 384 
rect 258 384 261 387 
rect 258 387 261 390 
rect 258 390 261 393 
rect 258 393 261 396 
rect 258 396 261 399 
rect 258 399 261 402 
rect 258 402 261 405 
rect 258 405 261 408 
rect 258 408 261 411 
rect 258 411 261 414 
rect 258 414 261 417 
rect 258 417 261 420 
rect 258 420 261 423 
rect 258 423 261 426 
rect 258 426 261 429 
rect 258 429 261 432 
rect 258 432 261 435 
rect 258 435 261 438 
rect 258 438 261 441 
rect 258 441 261 444 
rect 258 444 261 447 
rect 258 447 261 450 
rect 258 450 261 453 
rect 258 453 261 456 
rect 258 456 261 459 
rect 258 459 261 462 
rect 258 462 261 465 
rect 258 465 261 468 
rect 258 468 261 471 
rect 258 471 261 474 
rect 258 474 261 477 
rect 258 477 261 480 
rect 258 480 261 483 
rect 258 483 261 486 
rect 258 486 261 489 
rect 258 489 261 492 
rect 258 492 261 495 
rect 258 495 261 498 
rect 258 498 261 501 
rect 258 501 261 504 
rect 258 504 261 507 
rect 258 507 261 510 
rect 261 0 264 3 
rect 261 3 264 6 
rect 261 6 264 9 
rect 261 9 264 12 
rect 261 12 264 15 
rect 261 15 264 18 
rect 261 18 264 21 
rect 261 21 264 24 
rect 261 24 264 27 
rect 261 27 264 30 
rect 261 30 264 33 
rect 261 33 264 36 
rect 261 36 264 39 
rect 261 39 264 42 
rect 261 42 264 45 
rect 261 45 264 48 
rect 261 48 264 51 
rect 261 51 264 54 
rect 261 54 264 57 
rect 261 57 264 60 
rect 261 60 264 63 
rect 261 63 264 66 
rect 261 66 264 69 
rect 261 69 264 72 
rect 261 72 264 75 
rect 261 75 264 78 
rect 261 78 264 81 
rect 261 81 264 84 
rect 261 84 264 87 
rect 261 87 264 90 
rect 261 90 264 93 
rect 261 93 264 96 
rect 261 96 264 99 
rect 261 99 264 102 
rect 261 102 264 105 
rect 261 105 264 108 
rect 261 108 264 111 
rect 261 111 264 114 
rect 261 114 264 117 
rect 261 117 264 120 
rect 261 120 264 123 
rect 261 123 264 126 
rect 261 126 264 129 
rect 261 129 264 132 
rect 261 132 264 135 
rect 261 135 264 138 
rect 261 138 264 141 
rect 261 141 264 144 
rect 261 144 264 147 
rect 261 147 264 150 
rect 261 150 264 153 
rect 261 153 264 156 
rect 261 156 264 159 
rect 261 159 264 162 
rect 261 162 264 165 
rect 261 165 264 168 
rect 261 168 264 171 
rect 261 171 264 174 
rect 261 174 264 177 
rect 261 177 264 180 
rect 261 180 264 183 
rect 261 183 264 186 
rect 261 186 264 189 
rect 261 189 264 192 
rect 261 192 264 195 
rect 261 195 264 198 
rect 261 198 264 201 
rect 261 201 264 204 
rect 261 204 264 207 
rect 261 207 264 210 
rect 261 210 264 213 
rect 261 213 264 216 
rect 261 216 264 219 
rect 261 219 264 222 
rect 261 222 264 225 
rect 261 225 264 228 
rect 261 228 264 231 
rect 261 231 264 234 
rect 261 234 264 237 
rect 261 237 264 240 
rect 261 240 264 243 
rect 261 243 264 246 
rect 261 246 264 249 
rect 261 249 264 252 
rect 261 252 264 255 
rect 261 255 264 258 
rect 261 258 264 261 
rect 261 261 264 264 
rect 261 264 264 267 
rect 261 267 264 270 
rect 261 270 264 273 
rect 261 273 264 276 
rect 261 276 264 279 
rect 261 279 264 282 
rect 261 282 264 285 
rect 261 285 264 288 
rect 261 288 264 291 
rect 261 291 264 294 
rect 261 294 264 297 
rect 261 297 264 300 
rect 261 300 264 303 
rect 261 303 264 306 
rect 261 306 264 309 
rect 261 309 264 312 
rect 261 312 264 315 
rect 261 315 264 318 
rect 261 318 264 321 
rect 261 321 264 324 
rect 261 324 264 327 
rect 261 327 264 330 
rect 261 330 264 333 
rect 261 333 264 336 
rect 261 336 264 339 
rect 261 339 264 342 
rect 261 342 264 345 
rect 261 345 264 348 
rect 261 348 264 351 
rect 261 351 264 354 
rect 261 354 264 357 
rect 261 357 264 360 
rect 261 360 264 363 
rect 261 363 264 366 
rect 261 366 264 369 
rect 261 369 264 372 
rect 261 372 264 375 
rect 261 375 264 378 
rect 261 378 264 381 
rect 261 381 264 384 
rect 261 384 264 387 
rect 261 387 264 390 
rect 261 390 264 393 
rect 261 393 264 396 
rect 261 396 264 399 
rect 261 399 264 402 
rect 261 402 264 405 
rect 261 405 264 408 
rect 261 408 264 411 
rect 261 411 264 414 
rect 261 414 264 417 
rect 261 417 264 420 
rect 261 420 264 423 
rect 261 423 264 426 
rect 261 426 264 429 
rect 261 429 264 432 
rect 261 432 264 435 
rect 261 435 264 438 
rect 261 438 264 441 
rect 261 441 264 444 
rect 261 444 264 447 
rect 261 447 264 450 
rect 261 450 264 453 
rect 261 453 264 456 
rect 261 456 264 459 
rect 261 459 264 462 
rect 261 462 264 465 
rect 261 465 264 468 
rect 261 468 264 471 
rect 261 471 264 474 
rect 261 474 264 477 
rect 261 477 264 480 
rect 261 480 264 483 
rect 261 483 264 486 
rect 261 486 264 489 
rect 261 489 264 492 
rect 261 492 264 495 
rect 261 495 264 498 
rect 261 498 264 501 
rect 261 501 264 504 
rect 261 504 264 507 
rect 261 507 264 510 
rect 264 0 267 3 
rect 264 3 267 6 
rect 264 6 267 9 
rect 264 9 267 12 
rect 264 12 267 15 
rect 264 15 267 18 
rect 264 18 267 21 
rect 264 21 267 24 
rect 264 24 267 27 
rect 264 27 267 30 
rect 264 30 267 33 
rect 264 33 267 36 
rect 264 36 267 39 
rect 264 39 267 42 
rect 264 42 267 45 
rect 264 45 267 48 
rect 264 48 267 51 
rect 264 51 267 54 
rect 264 54 267 57 
rect 264 57 267 60 
rect 264 60 267 63 
rect 264 63 267 66 
rect 264 66 267 69 
rect 264 69 267 72 
rect 264 72 267 75 
rect 264 75 267 78 
rect 264 78 267 81 
rect 264 81 267 84 
rect 264 84 267 87 
rect 264 87 267 90 
rect 264 90 267 93 
rect 264 93 267 96 
rect 264 96 267 99 
rect 264 99 267 102 
rect 264 102 267 105 
rect 264 105 267 108 
rect 264 108 267 111 
rect 264 111 267 114 
rect 264 114 267 117 
rect 264 117 267 120 
rect 264 120 267 123 
rect 264 123 267 126 
rect 264 126 267 129 
rect 264 129 267 132 
rect 264 132 267 135 
rect 264 135 267 138 
rect 264 138 267 141 
rect 264 141 267 144 
rect 264 144 267 147 
rect 264 147 267 150 
rect 264 150 267 153 
rect 264 153 267 156 
rect 264 156 267 159 
rect 264 159 267 162 
rect 264 162 267 165 
rect 264 165 267 168 
rect 264 168 267 171 
rect 264 171 267 174 
rect 264 174 267 177 
rect 264 177 267 180 
rect 264 180 267 183 
rect 264 183 267 186 
rect 264 186 267 189 
rect 264 189 267 192 
rect 264 192 267 195 
rect 264 195 267 198 
rect 264 198 267 201 
rect 264 201 267 204 
rect 264 204 267 207 
rect 264 207 267 210 
rect 264 210 267 213 
rect 264 213 267 216 
rect 264 216 267 219 
rect 264 219 267 222 
rect 264 222 267 225 
rect 264 225 267 228 
rect 264 228 267 231 
rect 264 231 267 234 
rect 264 234 267 237 
rect 264 237 267 240 
rect 264 240 267 243 
rect 264 243 267 246 
rect 264 246 267 249 
rect 264 249 267 252 
rect 264 252 267 255 
rect 264 255 267 258 
rect 264 258 267 261 
rect 264 261 267 264 
rect 264 264 267 267 
rect 264 267 267 270 
rect 264 270 267 273 
rect 264 273 267 276 
rect 264 276 267 279 
rect 264 279 267 282 
rect 264 282 267 285 
rect 264 285 267 288 
rect 264 288 267 291 
rect 264 291 267 294 
rect 264 294 267 297 
rect 264 297 267 300 
rect 264 300 267 303 
rect 264 303 267 306 
rect 264 306 267 309 
rect 264 309 267 312 
rect 264 312 267 315 
rect 264 315 267 318 
rect 264 318 267 321 
rect 264 321 267 324 
rect 264 324 267 327 
rect 264 327 267 330 
rect 264 330 267 333 
rect 264 333 267 336 
rect 264 336 267 339 
rect 264 339 267 342 
rect 264 342 267 345 
rect 264 345 267 348 
rect 264 348 267 351 
rect 264 351 267 354 
rect 264 354 267 357 
rect 264 357 267 360 
rect 264 360 267 363 
rect 264 363 267 366 
rect 264 366 267 369 
rect 264 369 267 372 
rect 264 372 267 375 
rect 264 375 267 378 
rect 264 378 267 381 
rect 264 381 267 384 
rect 264 384 267 387 
rect 264 387 267 390 
rect 264 390 267 393 
rect 264 393 267 396 
rect 264 396 267 399 
rect 264 399 267 402 
rect 264 402 267 405 
rect 264 405 267 408 
rect 264 408 267 411 
rect 264 411 267 414 
rect 264 414 267 417 
rect 264 417 267 420 
rect 264 420 267 423 
rect 264 423 267 426 
rect 264 426 267 429 
rect 264 429 267 432 
rect 264 432 267 435 
rect 264 435 267 438 
rect 264 438 267 441 
rect 264 441 267 444 
rect 264 444 267 447 
rect 264 447 267 450 
rect 264 450 267 453 
rect 264 453 267 456 
rect 264 456 267 459 
rect 264 459 267 462 
rect 264 462 267 465 
rect 264 465 267 468 
rect 264 468 267 471 
rect 264 471 267 474 
rect 264 474 267 477 
rect 264 477 267 480 
rect 264 480 267 483 
rect 264 483 267 486 
rect 264 486 267 489 
rect 264 489 267 492 
rect 264 492 267 495 
rect 264 495 267 498 
rect 264 498 267 501 
rect 264 501 267 504 
rect 264 504 267 507 
rect 264 507 267 510 
rect 267 0 270 3 
rect 267 3 270 6 
rect 267 6 270 9 
rect 267 9 270 12 
rect 267 12 270 15 
rect 267 15 270 18 
rect 267 18 270 21 
rect 267 21 270 24 
rect 267 24 270 27 
rect 267 27 270 30 
rect 267 30 270 33 
rect 267 33 270 36 
rect 267 36 270 39 
rect 267 39 270 42 
rect 267 42 270 45 
rect 267 45 270 48 
rect 267 48 270 51 
rect 267 51 270 54 
rect 267 54 270 57 
rect 267 57 270 60 
rect 267 60 270 63 
rect 267 63 270 66 
rect 267 66 270 69 
rect 267 69 270 72 
rect 267 72 270 75 
rect 267 75 270 78 
rect 267 78 270 81 
rect 267 81 270 84 
rect 267 84 270 87 
rect 267 87 270 90 
rect 267 90 270 93 
rect 267 93 270 96 
rect 267 96 270 99 
rect 267 99 270 102 
rect 267 102 270 105 
rect 267 105 270 108 
rect 267 108 270 111 
rect 267 111 270 114 
rect 267 114 270 117 
rect 267 117 270 120 
rect 267 120 270 123 
rect 267 123 270 126 
rect 267 126 270 129 
rect 267 129 270 132 
rect 267 132 270 135 
rect 267 135 270 138 
rect 267 138 270 141 
rect 267 141 270 144 
rect 267 144 270 147 
rect 267 147 270 150 
rect 267 150 270 153 
rect 267 153 270 156 
rect 267 156 270 159 
rect 267 159 270 162 
rect 267 162 270 165 
rect 267 165 270 168 
rect 267 168 270 171 
rect 267 171 270 174 
rect 267 174 270 177 
rect 267 177 270 180 
rect 267 180 270 183 
rect 267 183 270 186 
rect 267 186 270 189 
rect 267 189 270 192 
rect 267 192 270 195 
rect 267 195 270 198 
rect 267 198 270 201 
rect 267 201 270 204 
rect 267 204 270 207 
rect 267 207 270 210 
rect 267 210 270 213 
rect 267 213 270 216 
rect 267 216 270 219 
rect 267 219 270 222 
rect 267 222 270 225 
rect 267 225 270 228 
rect 267 228 270 231 
rect 267 231 270 234 
rect 267 234 270 237 
rect 267 237 270 240 
rect 267 240 270 243 
rect 267 243 270 246 
rect 267 246 270 249 
rect 267 249 270 252 
rect 267 252 270 255 
rect 267 255 270 258 
rect 267 258 270 261 
rect 267 261 270 264 
rect 267 264 270 267 
rect 267 267 270 270 
rect 267 270 270 273 
rect 267 273 270 276 
rect 267 276 270 279 
rect 267 279 270 282 
rect 267 282 270 285 
rect 267 285 270 288 
rect 267 288 270 291 
rect 267 291 270 294 
rect 267 294 270 297 
rect 267 297 270 300 
rect 267 300 270 303 
rect 267 303 270 306 
rect 267 306 270 309 
rect 267 309 270 312 
rect 267 312 270 315 
rect 267 315 270 318 
rect 267 318 270 321 
rect 267 321 270 324 
rect 267 324 270 327 
rect 267 327 270 330 
rect 267 330 270 333 
rect 267 333 270 336 
rect 267 336 270 339 
rect 267 339 270 342 
rect 267 342 270 345 
rect 267 345 270 348 
rect 267 348 270 351 
rect 267 351 270 354 
rect 267 354 270 357 
rect 267 357 270 360 
rect 267 360 270 363 
rect 267 363 270 366 
rect 267 366 270 369 
rect 267 369 270 372 
rect 267 372 270 375 
rect 267 375 270 378 
rect 267 378 270 381 
rect 267 381 270 384 
rect 267 384 270 387 
rect 267 387 270 390 
rect 267 390 270 393 
rect 267 393 270 396 
rect 267 396 270 399 
rect 267 399 270 402 
rect 267 402 270 405 
rect 267 405 270 408 
rect 267 408 270 411 
rect 267 411 270 414 
rect 267 414 270 417 
rect 267 417 270 420 
rect 267 420 270 423 
rect 267 423 270 426 
rect 267 426 270 429 
rect 267 429 270 432 
rect 267 432 270 435 
rect 267 435 270 438 
rect 267 438 270 441 
rect 267 441 270 444 
rect 267 444 270 447 
rect 267 447 270 450 
rect 267 450 270 453 
rect 267 453 270 456 
rect 267 456 270 459 
rect 267 459 270 462 
rect 267 462 270 465 
rect 267 465 270 468 
rect 267 468 270 471 
rect 267 471 270 474 
rect 267 474 270 477 
rect 267 477 270 480 
rect 267 480 270 483 
rect 267 483 270 486 
rect 267 486 270 489 
rect 267 489 270 492 
rect 267 492 270 495 
rect 267 495 270 498 
rect 267 498 270 501 
rect 267 501 270 504 
rect 267 504 270 507 
rect 267 507 270 510 
rect 270 0 273 3 
rect 270 3 273 6 
rect 270 6 273 9 
rect 270 9 273 12 
rect 270 12 273 15 
rect 270 15 273 18 
rect 270 18 273 21 
rect 270 21 273 24 
rect 270 24 273 27 
rect 270 27 273 30 
rect 270 30 273 33 
rect 270 33 273 36 
rect 270 36 273 39 
rect 270 39 273 42 
rect 270 42 273 45 
rect 270 45 273 48 
rect 270 48 273 51 
rect 270 51 273 54 
rect 270 54 273 57 
rect 270 57 273 60 
rect 270 60 273 63 
rect 270 63 273 66 
rect 270 66 273 69 
rect 270 69 273 72 
rect 270 72 273 75 
rect 270 75 273 78 
rect 270 78 273 81 
rect 270 84 273 87 
rect 270 87 273 90 
rect 270 90 273 93 
rect 270 93 273 96 
rect 270 96 273 99 
rect 270 99 273 102 
rect 270 102 273 105 
rect 270 105 273 108 
rect 270 108 273 111 
rect 270 111 273 114 
rect 270 114 273 117 
rect 270 117 273 120 
rect 270 120 273 123 
rect 270 123 273 126 
rect 270 126 273 129 
rect 270 129 273 132 
rect 270 132 273 135 
rect 270 135 273 138 
rect 270 138 273 141 
rect 270 141 273 144 
rect 270 144 273 147 
rect 270 147 273 150 
rect 270 150 273 153 
rect 270 153 273 156 
rect 270 156 273 159 
rect 270 159 273 162 
rect 270 162 273 165 
rect 270 165 273 168 
rect 270 168 273 171 
rect 270 171 273 174 
rect 270 174 273 177 
rect 270 180 273 183 
rect 270 183 273 186 
rect 270 186 273 189 
rect 270 189 273 192 
rect 270 192 273 195 
rect 270 195 273 198 
rect 270 198 273 201 
rect 270 201 273 204 
rect 270 204 273 207 
rect 270 207 273 210 
rect 270 210 273 213 
rect 270 213 273 216 
rect 270 216 273 219 
rect 270 219 273 222 
rect 270 222 273 225 
rect 270 225 273 228 
rect 270 228 273 231 
rect 270 231 273 234 
rect 270 234 273 237 
rect 270 237 273 240 
rect 270 240 273 243 
rect 270 243 273 246 
rect 270 246 273 249 
rect 270 249 273 252 
rect 270 252 273 255 
rect 270 255 273 258 
rect 270 258 273 261 
rect 270 261 273 264 
rect 270 264 273 267 
rect 270 267 273 270 
rect 270 270 273 273 
rect 270 273 273 276 
rect 270 276 273 279 
rect 270 279 273 282 
rect 270 282 273 285 
rect 270 285 273 288 
rect 270 288 273 291 
rect 270 291 273 294 
rect 270 294 273 297 
rect 270 297 273 300 
rect 270 300 273 303 
rect 270 303 273 306 
rect 270 306 273 309 
rect 270 309 273 312 
rect 270 312 273 315 
rect 270 315 273 318 
rect 270 318 273 321 
rect 270 321 273 324 
rect 270 324 273 327 
rect 270 327 273 330 
rect 270 330 273 333 
rect 270 333 273 336 
rect 270 336 273 339 
rect 270 339 273 342 
rect 270 342 273 345 
rect 270 345 273 348 
rect 270 348 273 351 
rect 270 351 273 354 
rect 270 354 273 357 
rect 270 357 273 360 
rect 270 360 273 363 
rect 270 363 273 366 
rect 270 366 273 369 
rect 270 369 273 372 
rect 270 372 273 375 
rect 270 375 273 378 
rect 270 381 273 384 
rect 270 384 273 387 
rect 270 387 273 390 
rect 270 390 273 393 
rect 270 393 273 396 
rect 270 396 273 399 
rect 270 399 273 402 
rect 270 402 273 405 
rect 270 405 273 408 
rect 270 408 273 411 
rect 270 411 273 414 
rect 270 414 273 417 
rect 270 420 273 423 
rect 270 423 273 426 
rect 270 429 273 432 
rect 270 432 273 435 
rect 270 435 273 438 
rect 270 438 273 441 
rect 270 441 273 444 
rect 270 444 273 447 
rect 270 447 273 450 
rect 270 450 273 453 
rect 270 453 273 456 
rect 270 456 273 459 
rect 270 459 273 462 
rect 270 462 273 465 
rect 270 468 273 471 
rect 270 471 273 474 
rect 270 477 273 480 
rect 270 480 273 483 
rect 270 483 273 486 
rect 270 486 273 489 
rect 270 489 273 492 
rect 270 492 273 495 
rect 270 495 273 498 
rect 270 498 273 501 
rect 270 501 273 504 
rect 270 504 273 507 
rect 270 507 273 510 
rect 273 0 276 3 
rect 273 3 276 6 
rect 273 6 276 9 
rect 273 9 276 12 
rect 273 12 276 15 
rect 273 15 276 18 
rect 273 18 276 21 
rect 273 21 276 24 
rect 273 24 276 27 
rect 273 27 276 30 
rect 273 30 276 33 
rect 273 33 276 36 
rect 273 36 276 39 
rect 273 39 276 42 
rect 273 42 276 45 
rect 273 45 276 48 
rect 273 48 276 51 
rect 273 51 276 54 
rect 273 54 276 57 
rect 273 57 276 60 
rect 273 60 276 63 
rect 273 63 276 66 
rect 273 66 276 69 
rect 273 69 276 72 
rect 273 72 276 75 
rect 273 75 276 78 
rect 273 78 276 81 
rect 273 81 276 84 
rect 273 84 276 87 
rect 273 87 276 90 
rect 273 90 276 93 
rect 273 93 276 96 
rect 273 96 276 99 
rect 273 99 276 102 
rect 273 102 276 105 
rect 273 105 276 108 
rect 273 108 276 111 
rect 273 111 276 114 
rect 273 114 276 117 
rect 273 117 276 120 
rect 273 120 276 123 
rect 273 123 276 126 
rect 273 126 276 129 
rect 273 129 276 132 
rect 273 132 276 135 
rect 273 135 276 138 
rect 273 138 276 141 
rect 273 141 276 144 
rect 273 144 276 147 
rect 273 147 276 150 
rect 273 150 276 153 
rect 273 153 276 156 
rect 273 156 276 159 
rect 273 159 276 162 
rect 273 162 276 165 
rect 273 165 276 168 
rect 273 168 276 171 
rect 273 171 276 174 
rect 273 174 276 177 
rect 273 177 276 180 
rect 273 180 276 183 
rect 273 183 276 186 
rect 273 186 276 189 
rect 273 189 276 192 
rect 273 192 276 195 
rect 273 195 276 198 
rect 273 198 276 201 
rect 273 201 276 204 
rect 273 204 276 207 
rect 273 207 276 210 
rect 273 210 276 213 
rect 273 213 276 216 
rect 273 216 276 219 
rect 273 219 276 222 
rect 273 222 276 225 
rect 273 225 276 228 
rect 273 228 276 231 
rect 273 231 276 234 
rect 273 234 276 237 
rect 273 237 276 240 
rect 273 240 276 243 
rect 273 243 276 246 
rect 273 246 276 249 
rect 273 249 276 252 
rect 273 252 276 255 
rect 273 255 276 258 
rect 273 258 276 261 
rect 273 261 276 264 
rect 273 264 276 267 
rect 273 267 276 270 
rect 273 270 276 273 
rect 273 273 276 276 
rect 273 276 276 279 
rect 273 279 276 282 
rect 273 282 276 285 
rect 273 285 276 288 
rect 273 288 276 291 
rect 273 291 276 294 
rect 273 294 276 297 
rect 273 297 276 300 
rect 273 300 276 303 
rect 273 303 276 306 
rect 273 306 276 309 
rect 273 309 276 312 
rect 273 312 276 315 
rect 273 315 276 318 
rect 273 318 276 321 
rect 273 321 276 324 
rect 273 324 276 327 
rect 273 327 276 330 
rect 273 330 276 333 
rect 273 333 276 336 
rect 273 336 276 339 
rect 273 339 276 342 
rect 273 342 276 345 
rect 273 345 276 348 
rect 273 348 276 351 
rect 273 351 276 354 
rect 273 354 276 357 
rect 273 357 276 360 
rect 273 360 276 363 
rect 273 363 276 366 
rect 273 366 276 369 
rect 273 369 276 372 
rect 273 372 276 375 
rect 273 375 276 378 
rect 273 378 276 381 
rect 273 381 276 384 
rect 273 384 276 387 
rect 273 387 276 390 
rect 273 390 276 393 
rect 273 393 276 396 
rect 273 396 276 399 
rect 273 399 276 402 
rect 273 402 276 405 
rect 273 405 276 408 
rect 273 408 276 411 
rect 273 411 276 414 
rect 273 414 276 417 
rect 273 417 276 420 
rect 273 420 276 423 
rect 273 423 276 426 
rect 273 426 276 429 
rect 273 429 276 432 
rect 273 432 276 435 
rect 273 435 276 438 
rect 273 438 276 441 
rect 273 441 276 444 
rect 273 444 276 447 
rect 273 447 276 450 
rect 273 450 276 453 
rect 273 453 276 456 
rect 273 456 276 459 
rect 273 459 276 462 
rect 273 462 276 465 
rect 273 465 276 468 
rect 273 468 276 471 
rect 273 471 276 474 
rect 273 474 276 477 
rect 273 477 276 480 
rect 273 480 276 483 
rect 273 483 276 486 
rect 273 486 276 489 
rect 273 489 276 492 
rect 273 492 276 495 
rect 273 495 276 498 
rect 273 498 276 501 
rect 273 501 276 504 
rect 273 504 276 507 
rect 273 507 276 510 
rect 276 0 279 3 
rect 276 3 279 6 
rect 276 6 279 9 
rect 276 9 279 12 
rect 276 12 279 15 
rect 276 15 279 18 
rect 276 18 279 21 
rect 276 21 279 24 
rect 276 24 279 27 
rect 276 27 279 30 
rect 276 30 279 33 
rect 276 33 279 36 
rect 276 36 279 39 
rect 276 39 279 42 
rect 276 42 279 45 
rect 276 45 279 48 
rect 276 48 279 51 
rect 276 51 279 54 
rect 276 54 279 57 
rect 276 57 279 60 
rect 276 60 279 63 
rect 276 63 279 66 
rect 276 66 279 69 
rect 276 69 279 72 
rect 276 72 279 75 
rect 276 75 279 78 
rect 276 78 279 81 
rect 276 81 279 84 
rect 276 84 279 87 
rect 276 87 279 90 
rect 276 90 279 93 
rect 276 93 279 96 
rect 276 96 279 99 
rect 276 99 279 102 
rect 276 102 279 105 
rect 276 105 279 108 
rect 276 108 279 111 
rect 276 111 279 114 
rect 276 114 279 117 
rect 276 117 279 120 
rect 276 120 279 123 
rect 276 123 279 126 
rect 276 126 279 129 
rect 276 129 279 132 
rect 276 132 279 135 
rect 276 135 279 138 
rect 276 138 279 141 
rect 276 141 279 144 
rect 276 144 279 147 
rect 276 147 279 150 
rect 276 150 279 153 
rect 276 153 279 156 
rect 276 156 279 159 
rect 276 159 279 162 
rect 276 162 279 165 
rect 276 165 279 168 
rect 276 168 279 171 
rect 276 171 279 174 
rect 276 174 279 177 
rect 276 177 279 180 
rect 276 180 279 183 
rect 276 183 279 186 
rect 276 186 279 189 
rect 276 189 279 192 
rect 276 192 279 195 
rect 276 195 279 198 
rect 276 198 279 201 
rect 276 201 279 204 
rect 276 204 279 207 
rect 276 207 279 210 
rect 276 210 279 213 
rect 276 213 279 216 
rect 276 216 279 219 
rect 276 219 279 222 
rect 276 222 279 225 
rect 276 225 279 228 
rect 276 228 279 231 
rect 276 231 279 234 
rect 276 234 279 237 
rect 276 237 279 240 
rect 276 240 279 243 
rect 276 243 279 246 
rect 276 246 279 249 
rect 276 249 279 252 
rect 276 252 279 255 
rect 276 255 279 258 
rect 276 258 279 261 
rect 276 261 279 264 
rect 276 264 279 267 
rect 276 267 279 270 
rect 276 270 279 273 
rect 276 273 279 276 
rect 276 276 279 279 
rect 276 279 279 282 
rect 276 282 279 285 
rect 276 285 279 288 
rect 276 288 279 291 
rect 276 291 279 294 
rect 276 294 279 297 
rect 276 297 279 300 
rect 276 300 279 303 
rect 276 303 279 306 
rect 276 306 279 309 
rect 276 309 279 312 
rect 276 312 279 315 
rect 276 315 279 318 
rect 276 318 279 321 
rect 276 321 279 324 
rect 276 324 279 327 
rect 276 327 279 330 
rect 276 330 279 333 
rect 276 333 279 336 
rect 276 336 279 339 
rect 276 339 279 342 
rect 276 342 279 345 
rect 276 345 279 348 
rect 276 348 279 351 
rect 276 351 279 354 
rect 276 354 279 357 
rect 276 357 279 360 
rect 276 360 279 363 
rect 276 363 279 366 
rect 276 366 279 369 
rect 276 369 279 372 
rect 276 372 279 375 
rect 276 375 279 378 
rect 276 378 279 381 
rect 276 381 279 384 
rect 276 384 279 387 
rect 276 387 279 390 
rect 276 390 279 393 
rect 276 393 279 396 
rect 276 396 279 399 
rect 276 399 279 402 
rect 276 402 279 405 
rect 276 405 279 408 
rect 276 408 279 411 
rect 276 411 279 414 
rect 276 414 279 417 
rect 276 417 279 420 
rect 276 420 279 423 
rect 276 423 279 426 
rect 276 426 279 429 
rect 276 429 279 432 
rect 276 432 279 435 
rect 276 435 279 438 
rect 276 438 279 441 
rect 276 441 279 444 
rect 276 444 279 447 
rect 276 447 279 450 
rect 276 450 279 453 
rect 276 453 279 456 
rect 276 456 279 459 
rect 276 459 279 462 
rect 276 462 279 465 
rect 276 465 279 468 
rect 276 468 279 471 
rect 276 471 279 474 
rect 276 474 279 477 
rect 276 477 279 480 
rect 276 480 279 483 
rect 276 483 279 486 
rect 276 486 279 489 
rect 276 489 279 492 
rect 276 492 279 495 
rect 276 495 279 498 
rect 276 498 279 501 
rect 276 501 279 504 
rect 276 504 279 507 
rect 276 507 279 510 
rect 279 0 282 3 
rect 279 3 282 6 
rect 279 6 282 9 
rect 279 9 282 12 
rect 279 12 282 15 
rect 279 15 282 18 
rect 279 18 282 21 
rect 279 21 282 24 
rect 279 24 282 27 
rect 279 27 282 30 
rect 279 30 282 33 
rect 279 33 282 36 
rect 279 36 282 39 
rect 279 39 282 42 
rect 279 42 282 45 
rect 279 45 282 48 
rect 279 48 282 51 
rect 279 51 282 54 
rect 279 54 282 57 
rect 279 57 282 60 
rect 279 60 282 63 
rect 279 63 282 66 
rect 279 66 282 69 
rect 279 69 282 72 
rect 279 72 282 75 
rect 279 75 282 78 
rect 279 78 282 81 
rect 279 81 282 84 
rect 279 84 282 87 
rect 279 87 282 90 
rect 279 90 282 93 
rect 279 93 282 96 
rect 279 96 282 99 
rect 279 99 282 102 
rect 279 102 282 105 
rect 279 105 282 108 
rect 279 108 282 111 
rect 279 111 282 114 
rect 279 114 282 117 
rect 279 117 282 120 
rect 279 120 282 123 
rect 279 123 282 126 
rect 279 126 282 129 
rect 279 129 282 132 
rect 279 132 282 135 
rect 279 135 282 138 
rect 279 138 282 141 
rect 279 141 282 144 
rect 279 144 282 147 
rect 279 147 282 150 
rect 279 150 282 153 
rect 279 153 282 156 
rect 279 156 282 159 
rect 279 159 282 162 
rect 279 162 282 165 
rect 279 165 282 168 
rect 279 168 282 171 
rect 279 171 282 174 
rect 279 174 282 177 
rect 279 177 282 180 
rect 279 180 282 183 
rect 279 183 282 186 
rect 279 186 282 189 
rect 279 189 282 192 
rect 279 192 282 195 
rect 279 195 282 198 
rect 279 198 282 201 
rect 279 201 282 204 
rect 279 204 282 207 
rect 279 207 282 210 
rect 279 210 282 213 
rect 279 213 282 216 
rect 279 216 282 219 
rect 279 219 282 222 
rect 279 222 282 225 
rect 279 225 282 228 
rect 279 228 282 231 
rect 279 231 282 234 
rect 279 234 282 237 
rect 279 237 282 240 
rect 279 240 282 243 
rect 279 243 282 246 
rect 279 246 282 249 
rect 279 249 282 252 
rect 279 252 282 255 
rect 279 255 282 258 
rect 279 258 282 261 
rect 279 261 282 264 
rect 279 264 282 267 
rect 279 267 282 270 
rect 279 270 282 273 
rect 279 273 282 276 
rect 279 276 282 279 
rect 279 279 282 282 
rect 279 282 282 285 
rect 279 285 282 288 
rect 279 288 282 291 
rect 279 291 282 294 
rect 279 294 282 297 
rect 279 297 282 300 
rect 279 300 282 303 
rect 279 303 282 306 
rect 279 306 282 309 
rect 279 309 282 312 
rect 279 312 282 315 
rect 279 315 282 318 
rect 279 318 282 321 
rect 279 321 282 324 
rect 279 324 282 327 
rect 279 327 282 330 
rect 279 330 282 333 
rect 279 333 282 336 
rect 279 336 282 339 
rect 279 339 282 342 
rect 279 342 282 345 
rect 279 345 282 348 
rect 279 348 282 351 
rect 279 351 282 354 
rect 279 354 282 357 
rect 279 357 282 360 
rect 279 360 282 363 
rect 279 363 282 366 
rect 279 366 282 369 
rect 279 369 282 372 
rect 279 372 282 375 
rect 279 375 282 378 
rect 279 378 282 381 
rect 279 381 282 384 
rect 279 384 282 387 
rect 279 387 282 390 
rect 279 390 282 393 
rect 279 393 282 396 
rect 279 396 282 399 
rect 279 399 282 402 
rect 279 402 282 405 
rect 279 405 282 408 
rect 279 408 282 411 
rect 279 411 282 414 
rect 279 414 282 417 
rect 279 417 282 420 
rect 279 420 282 423 
rect 279 423 282 426 
rect 279 426 282 429 
rect 279 429 282 432 
rect 279 432 282 435 
rect 279 435 282 438 
rect 279 438 282 441 
rect 279 441 282 444 
rect 279 444 282 447 
rect 279 447 282 450 
rect 279 450 282 453 
rect 279 453 282 456 
rect 279 456 282 459 
rect 279 459 282 462 
rect 279 462 282 465 
rect 279 465 282 468 
rect 279 468 282 471 
rect 279 471 282 474 
rect 279 474 282 477 
rect 279 477 282 480 
rect 279 480 282 483 
rect 279 483 282 486 
rect 279 486 282 489 
rect 279 489 282 492 
rect 279 492 282 495 
rect 279 495 282 498 
rect 279 498 282 501 
rect 279 501 282 504 
rect 279 504 282 507 
rect 279 507 282 510 
rect 282 0 285 3 
rect 282 3 285 6 
rect 282 6 285 9 
rect 282 9 285 12 
rect 282 12 285 15 
rect 282 15 285 18 
rect 282 18 285 21 
rect 282 21 285 24 
rect 282 24 285 27 
rect 282 27 285 30 
rect 282 30 285 33 
rect 282 33 285 36 
rect 282 36 285 39 
rect 282 39 285 42 
rect 282 42 285 45 
rect 282 45 285 48 
rect 282 48 285 51 
rect 282 51 285 54 
rect 282 54 285 57 
rect 282 57 285 60 
rect 282 60 285 63 
rect 282 63 285 66 
rect 282 66 285 69 
rect 282 69 285 72 
rect 282 72 285 75 
rect 282 75 285 78 
rect 282 78 285 81 
rect 282 81 285 84 
rect 282 84 285 87 
rect 282 87 285 90 
rect 282 90 285 93 
rect 282 93 285 96 
rect 282 96 285 99 
rect 282 99 285 102 
rect 282 102 285 105 
rect 282 105 285 108 
rect 282 108 285 111 
rect 282 111 285 114 
rect 282 114 285 117 
rect 282 117 285 120 
rect 282 120 285 123 
rect 282 123 285 126 
rect 282 126 285 129 
rect 282 129 285 132 
rect 282 132 285 135 
rect 282 135 285 138 
rect 282 138 285 141 
rect 282 141 285 144 
rect 282 144 285 147 
rect 282 147 285 150 
rect 282 150 285 153 
rect 282 153 285 156 
rect 282 156 285 159 
rect 282 159 285 162 
rect 282 162 285 165 
rect 282 165 285 168 
rect 282 168 285 171 
rect 282 171 285 174 
rect 282 174 285 177 
rect 282 177 285 180 
rect 282 180 285 183 
rect 282 183 285 186 
rect 282 186 285 189 
rect 282 189 285 192 
rect 282 192 285 195 
rect 282 195 285 198 
rect 282 198 285 201 
rect 282 201 285 204 
rect 282 204 285 207 
rect 282 207 285 210 
rect 282 210 285 213 
rect 282 213 285 216 
rect 282 216 285 219 
rect 282 219 285 222 
rect 282 222 285 225 
rect 282 225 285 228 
rect 282 228 285 231 
rect 282 231 285 234 
rect 282 234 285 237 
rect 282 237 285 240 
rect 282 240 285 243 
rect 282 243 285 246 
rect 282 246 285 249 
rect 282 249 285 252 
rect 282 252 285 255 
rect 282 255 285 258 
rect 282 258 285 261 
rect 282 261 285 264 
rect 282 264 285 267 
rect 282 267 285 270 
rect 282 270 285 273 
rect 282 273 285 276 
rect 282 276 285 279 
rect 282 279 285 282 
rect 282 282 285 285 
rect 282 285 285 288 
rect 282 288 285 291 
rect 282 291 285 294 
rect 282 294 285 297 
rect 282 297 285 300 
rect 282 300 285 303 
rect 282 303 285 306 
rect 282 306 285 309 
rect 282 309 285 312 
rect 282 312 285 315 
rect 282 315 285 318 
rect 282 318 285 321 
rect 282 321 285 324 
rect 282 324 285 327 
rect 282 327 285 330 
rect 282 330 285 333 
rect 282 333 285 336 
rect 282 336 285 339 
rect 282 339 285 342 
rect 282 342 285 345 
rect 282 345 285 348 
rect 282 348 285 351 
rect 282 351 285 354 
rect 282 354 285 357 
rect 282 357 285 360 
rect 282 360 285 363 
rect 282 363 285 366 
rect 282 366 285 369 
rect 282 369 285 372 
rect 282 372 285 375 
rect 282 375 285 378 
rect 282 378 285 381 
rect 282 381 285 384 
rect 282 384 285 387 
rect 282 387 285 390 
rect 282 390 285 393 
rect 282 393 285 396 
rect 282 396 285 399 
rect 282 399 285 402 
rect 282 402 285 405 
rect 282 405 285 408 
rect 282 408 285 411 
rect 282 411 285 414 
rect 282 414 285 417 
rect 282 417 285 420 
rect 282 420 285 423 
rect 282 423 285 426 
rect 282 426 285 429 
rect 282 429 285 432 
rect 282 432 285 435 
rect 282 435 285 438 
rect 282 438 285 441 
rect 282 441 285 444 
rect 282 444 285 447 
rect 282 447 285 450 
rect 282 450 285 453 
rect 282 453 285 456 
rect 282 456 285 459 
rect 282 459 285 462 
rect 282 462 285 465 
rect 282 465 285 468 
rect 282 468 285 471 
rect 282 471 285 474 
rect 282 474 285 477 
rect 282 477 285 480 
rect 282 480 285 483 
rect 282 483 285 486 
rect 282 486 285 489 
rect 282 489 285 492 
rect 282 492 285 495 
rect 282 495 285 498 
rect 282 498 285 501 
rect 282 501 285 504 
rect 282 504 285 507 
rect 282 507 285 510 
rect 285 0 288 3 
rect 285 3 288 6 
rect 285 6 288 9 
rect 285 9 288 12 
rect 285 12 288 15 
rect 285 15 288 18 
rect 285 18 288 21 
rect 285 21 288 24 
rect 285 24 288 27 
rect 285 27 288 30 
rect 285 30 288 33 
rect 285 33 288 36 
rect 285 36 288 39 
rect 285 39 288 42 
rect 285 42 288 45 
rect 285 45 288 48 
rect 285 48 288 51 
rect 285 51 288 54 
rect 285 54 288 57 
rect 285 57 288 60 
rect 285 60 288 63 
rect 285 63 288 66 
rect 285 66 288 69 
rect 285 69 288 72 
rect 285 72 288 75 
rect 285 75 288 78 
rect 285 78 288 81 
rect 285 84 288 87 
rect 285 87 288 90 
rect 285 93 288 96 
rect 285 96 288 99 
rect 285 99 288 102 
rect 285 102 288 105 
rect 285 105 288 108 
rect 285 108 288 111 
rect 285 111 288 114 
rect 285 114 288 117 
rect 285 117 288 120 
rect 285 120 288 123 
rect 285 123 288 126 
rect 285 126 288 129 
rect 285 129 288 132 
rect 285 132 288 135 
rect 285 135 288 138 
rect 285 138 288 141 
rect 285 141 288 144 
rect 285 144 288 147 
rect 285 147 288 150 
rect 285 150 288 153 
rect 285 153 288 156 
rect 285 156 288 159 
rect 285 159 288 162 
rect 285 162 288 165 
rect 285 165 288 168 
rect 285 168 288 171 
rect 285 171 288 174 
rect 285 174 288 177 
rect 285 177 288 180 
rect 285 180 288 183 
rect 285 183 288 186 
rect 285 189 288 192 
rect 285 192 288 195 
rect 285 195 288 198 
rect 285 198 288 201 
rect 285 201 288 204 
rect 285 204 288 207 
rect 285 207 288 210 
rect 285 210 288 213 
rect 285 213 288 216 
rect 285 216 288 219 
rect 285 219 288 222 
rect 285 222 288 225 
rect 285 225 288 228 
rect 285 228 288 231 
rect 285 231 288 234 
rect 285 234 288 237 
rect 285 237 288 240 
rect 285 240 288 243 
rect 285 243 288 246 
rect 285 246 288 249 
rect 285 249 288 252 
rect 285 252 288 255 
rect 285 255 288 258 
rect 285 258 288 261 
rect 285 261 288 264 
rect 285 264 288 267 
rect 285 267 288 270 
rect 285 270 288 273 
rect 285 273 288 276 
rect 285 276 288 279 
rect 285 279 288 282 
rect 285 282 288 285 
rect 285 285 288 288 
rect 285 288 288 291 
rect 285 291 288 294 
rect 285 294 288 297 
rect 285 297 288 300 
rect 285 300 288 303 
rect 285 303 288 306 
rect 285 306 288 309 
rect 285 309 288 312 
rect 285 312 288 315 
rect 285 315 288 318 
rect 285 318 288 321 
rect 285 321 288 324 
rect 285 324 288 327 
rect 285 327 288 330 
rect 285 330 288 333 
rect 285 333 288 336 
rect 285 336 288 339 
rect 285 339 288 342 
rect 285 342 288 345 
rect 285 345 288 348 
rect 285 348 288 351 
rect 285 351 288 354 
rect 285 354 288 357 
rect 285 357 288 360 
rect 285 360 288 363 
rect 285 363 288 366 
rect 285 366 288 369 
rect 285 369 288 372 
rect 285 372 288 375 
rect 285 375 288 378 
rect 285 378 288 381 
rect 285 381 288 384 
rect 285 384 288 387 
rect 285 387 288 390 
rect 285 390 288 393 
rect 285 393 288 396 
rect 285 396 288 399 
rect 285 399 288 402 
rect 285 402 288 405 
rect 285 405 288 408 
rect 285 408 288 411 
rect 285 411 288 414 
rect 285 414 288 417 
rect 285 417 288 420 
rect 285 420 288 423 
rect 285 423 288 426 
rect 285 429 288 432 
rect 285 432 288 435 
rect 285 435 288 438 
rect 285 438 288 441 
rect 285 441 288 444 
rect 285 444 288 447 
rect 285 447 288 450 
rect 285 450 288 453 
rect 285 453 288 456 
rect 285 456 288 459 
rect 285 459 288 462 
rect 285 462 288 465 
rect 285 468 288 471 
rect 285 471 288 474 
rect 285 474 288 477 
rect 285 477 288 480 
rect 285 480 288 483 
rect 285 483 288 486 
rect 285 486 288 489 
rect 285 489 288 492 
rect 285 492 288 495 
rect 285 495 288 498 
rect 285 498 288 501 
rect 285 501 288 504 
rect 285 504 288 507 
rect 285 507 288 510 
rect 288 0 291 3 
rect 288 3 291 6 
rect 288 6 291 9 
rect 288 9 291 12 
rect 288 12 291 15 
rect 288 15 291 18 
rect 288 18 291 21 
rect 288 21 291 24 
rect 288 24 291 27 
rect 288 27 291 30 
rect 288 30 291 33 
rect 288 33 291 36 
rect 288 36 291 39 
rect 288 39 291 42 
rect 288 42 291 45 
rect 288 45 291 48 
rect 288 48 291 51 
rect 288 51 291 54 
rect 288 54 291 57 
rect 288 57 291 60 
rect 288 60 291 63 
rect 288 63 291 66 
rect 288 66 291 69 
rect 288 69 291 72 
rect 288 72 291 75 
rect 288 75 291 78 
rect 288 78 291 81 
rect 288 81 291 84 
rect 288 84 291 87 
rect 288 87 291 90 
rect 288 90 291 93 
rect 288 93 291 96 
rect 288 96 291 99 
rect 288 99 291 102 
rect 288 102 291 105 
rect 288 105 291 108 
rect 288 108 291 111 
rect 288 111 291 114 
rect 288 114 291 117 
rect 288 117 291 120 
rect 288 120 291 123 
rect 288 123 291 126 
rect 288 126 291 129 
rect 288 129 291 132 
rect 288 132 291 135 
rect 288 135 291 138 
rect 288 138 291 141 
rect 288 141 291 144 
rect 288 144 291 147 
rect 288 147 291 150 
rect 288 150 291 153 
rect 288 153 291 156 
rect 288 156 291 159 
rect 288 159 291 162 
rect 288 162 291 165 
rect 288 165 291 168 
rect 288 168 291 171 
rect 288 171 291 174 
rect 288 174 291 177 
rect 288 177 291 180 
rect 288 180 291 183 
rect 288 183 291 186 
rect 288 186 291 189 
rect 288 189 291 192 
rect 288 192 291 195 
rect 288 195 291 198 
rect 288 198 291 201 
rect 288 201 291 204 
rect 288 204 291 207 
rect 288 207 291 210 
rect 288 210 291 213 
rect 288 213 291 216 
rect 288 216 291 219 
rect 288 219 291 222 
rect 288 222 291 225 
rect 288 225 291 228 
rect 288 228 291 231 
rect 288 231 291 234 
rect 288 234 291 237 
rect 288 237 291 240 
rect 288 240 291 243 
rect 288 243 291 246 
rect 288 246 291 249 
rect 288 249 291 252 
rect 288 252 291 255 
rect 288 255 291 258 
rect 288 258 291 261 
rect 288 261 291 264 
rect 288 264 291 267 
rect 288 267 291 270 
rect 288 270 291 273 
rect 288 273 291 276 
rect 288 276 291 279 
rect 288 279 291 282 
rect 288 282 291 285 
rect 288 285 291 288 
rect 288 288 291 291 
rect 288 291 291 294 
rect 288 294 291 297 
rect 288 297 291 300 
rect 288 300 291 303 
rect 288 303 291 306 
rect 288 306 291 309 
rect 288 309 291 312 
rect 288 312 291 315 
rect 288 315 291 318 
rect 288 318 291 321 
rect 288 321 291 324 
rect 288 324 291 327 
rect 288 327 291 330 
rect 288 330 291 333 
rect 288 333 291 336 
rect 288 336 291 339 
rect 288 339 291 342 
rect 288 342 291 345 
rect 288 345 291 348 
rect 288 348 291 351 
rect 288 351 291 354 
rect 288 354 291 357 
rect 288 357 291 360 
rect 288 360 291 363 
rect 288 363 291 366 
rect 288 366 291 369 
rect 288 369 291 372 
rect 288 372 291 375 
rect 288 375 291 378 
rect 288 378 291 381 
rect 288 381 291 384 
rect 288 384 291 387 
rect 288 387 291 390 
rect 288 390 291 393 
rect 288 393 291 396 
rect 288 396 291 399 
rect 288 399 291 402 
rect 288 402 291 405 
rect 288 405 291 408 
rect 288 408 291 411 
rect 288 411 291 414 
rect 288 414 291 417 
rect 288 417 291 420 
rect 288 420 291 423 
rect 288 423 291 426 
rect 288 426 291 429 
rect 288 429 291 432 
rect 288 432 291 435 
rect 288 435 291 438 
rect 288 438 291 441 
rect 288 441 291 444 
rect 288 444 291 447 
rect 288 447 291 450 
rect 288 450 291 453 
rect 288 453 291 456 
rect 288 456 291 459 
rect 288 459 291 462 
rect 288 462 291 465 
rect 288 465 291 468 
rect 288 468 291 471 
rect 288 471 291 474 
rect 288 474 291 477 
rect 288 477 291 480 
rect 288 480 291 483 
rect 288 483 291 486 
rect 288 486 291 489 
rect 288 489 291 492 
rect 288 492 291 495 
rect 288 495 291 498 
rect 288 498 291 501 
rect 288 501 291 504 
rect 288 504 291 507 
rect 288 507 291 510 
rect 291 0 294 3 
rect 291 3 294 6 
rect 291 6 294 9 
rect 291 9 294 12 
rect 291 12 294 15 
rect 291 15 294 18 
rect 291 18 294 21 
rect 291 21 294 24 
rect 291 24 294 27 
rect 291 27 294 30 
rect 291 30 294 33 
rect 291 33 294 36 
rect 291 36 294 39 
rect 291 39 294 42 
rect 291 42 294 45 
rect 291 45 294 48 
rect 291 48 294 51 
rect 291 51 294 54 
rect 291 54 294 57 
rect 291 57 294 60 
rect 291 60 294 63 
rect 291 63 294 66 
rect 291 66 294 69 
rect 291 69 294 72 
rect 291 72 294 75 
rect 291 75 294 78 
rect 291 78 294 81 
rect 291 81 294 84 
rect 291 84 294 87 
rect 291 87 294 90 
rect 291 90 294 93 
rect 291 93 294 96 
rect 291 96 294 99 
rect 291 99 294 102 
rect 291 102 294 105 
rect 291 105 294 108 
rect 291 108 294 111 
rect 291 111 294 114 
rect 291 114 294 117 
rect 291 117 294 120 
rect 291 120 294 123 
rect 291 123 294 126 
rect 291 126 294 129 
rect 291 129 294 132 
rect 291 132 294 135 
rect 291 135 294 138 
rect 291 138 294 141 
rect 291 141 294 144 
rect 291 144 294 147 
rect 291 147 294 150 
rect 291 150 294 153 
rect 291 153 294 156 
rect 291 156 294 159 
rect 291 159 294 162 
rect 291 162 294 165 
rect 291 165 294 168 
rect 291 168 294 171 
rect 291 171 294 174 
rect 291 174 294 177 
rect 291 177 294 180 
rect 291 180 294 183 
rect 291 183 294 186 
rect 291 186 294 189 
rect 291 189 294 192 
rect 291 192 294 195 
rect 291 195 294 198 
rect 291 198 294 201 
rect 291 201 294 204 
rect 291 204 294 207 
rect 291 207 294 210 
rect 291 210 294 213 
rect 291 213 294 216 
rect 291 216 294 219 
rect 291 219 294 222 
rect 291 222 294 225 
rect 291 225 294 228 
rect 291 228 294 231 
rect 291 231 294 234 
rect 291 234 294 237 
rect 291 237 294 240 
rect 291 240 294 243 
rect 291 243 294 246 
rect 291 246 294 249 
rect 291 249 294 252 
rect 291 252 294 255 
rect 291 255 294 258 
rect 291 258 294 261 
rect 291 261 294 264 
rect 291 264 294 267 
rect 291 267 294 270 
rect 291 270 294 273 
rect 291 273 294 276 
rect 291 276 294 279 
rect 291 279 294 282 
rect 291 282 294 285 
rect 291 285 294 288 
rect 291 288 294 291 
rect 291 291 294 294 
rect 291 294 294 297 
rect 291 297 294 300 
rect 291 300 294 303 
rect 291 303 294 306 
rect 291 306 294 309 
rect 291 309 294 312 
rect 291 312 294 315 
rect 291 315 294 318 
rect 291 318 294 321 
rect 291 321 294 324 
rect 291 324 294 327 
rect 291 327 294 330 
rect 291 330 294 333 
rect 291 333 294 336 
rect 291 336 294 339 
rect 291 339 294 342 
rect 291 342 294 345 
rect 291 345 294 348 
rect 291 348 294 351 
rect 291 351 294 354 
rect 291 354 294 357 
rect 291 357 294 360 
rect 291 360 294 363 
rect 291 363 294 366 
rect 291 366 294 369 
rect 291 369 294 372 
rect 291 372 294 375 
rect 291 375 294 378 
rect 291 378 294 381 
rect 291 381 294 384 
rect 291 384 294 387 
rect 291 387 294 390 
rect 291 390 294 393 
rect 291 393 294 396 
rect 291 396 294 399 
rect 291 399 294 402 
rect 291 402 294 405 
rect 291 405 294 408 
rect 291 408 294 411 
rect 291 411 294 414 
rect 291 414 294 417 
rect 291 417 294 420 
rect 291 420 294 423 
rect 291 423 294 426 
rect 291 426 294 429 
rect 291 429 294 432 
rect 291 432 294 435 
rect 291 435 294 438 
rect 291 438 294 441 
rect 291 441 294 444 
rect 291 444 294 447 
rect 291 447 294 450 
rect 291 450 294 453 
rect 291 453 294 456 
rect 291 456 294 459 
rect 291 459 294 462 
rect 291 462 294 465 
rect 291 465 294 468 
rect 291 468 294 471 
rect 291 471 294 474 
rect 291 474 294 477 
rect 291 477 294 480 
rect 291 480 294 483 
rect 291 483 294 486 
rect 291 486 294 489 
rect 291 489 294 492 
rect 291 492 294 495 
rect 291 495 294 498 
rect 291 498 294 501 
rect 291 501 294 504 
rect 291 504 294 507 
rect 291 507 294 510 
rect 294 0 297 3 
rect 294 3 297 6 
rect 294 6 297 9 
rect 294 9 297 12 
rect 294 12 297 15 
rect 294 15 297 18 
rect 294 18 297 21 
rect 294 21 297 24 
rect 294 24 297 27 
rect 294 27 297 30 
rect 294 30 297 33 
rect 294 33 297 36 
rect 294 36 297 39 
rect 294 39 297 42 
rect 294 42 297 45 
rect 294 45 297 48 
rect 294 48 297 51 
rect 294 51 297 54 
rect 294 54 297 57 
rect 294 57 297 60 
rect 294 60 297 63 
rect 294 63 297 66 
rect 294 66 297 69 
rect 294 69 297 72 
rect 294 72 297 75 
rect 294 75 297 78 
rect 294 78 297 81 
rect 294 81 297 84 
rect 294 84 297 87 
rect 294 87 297 90 
rect 294 90 297 93 
rect 294 93 297 96 
rect 294 96 297 99 
rect 294 99 297 102 
rect 294 102 297 105 
rect 294 105 297 108 
rect 294 108 297 111 
rect 294 111 297 114 
rect 294 114 297 117 
rect 294 117 297 120 
rect 294 120 297 123 
rect 294 123 297 126 
rect 294 126 297 129 
rect 294 129 297 132 
rect 294 132 297 135 
rect 294 135 297 138 
rect 294 138 297 141 
rect 294 141 297 144 
rect 294 144 297 147 
rect 294 147 297 150 
rect 294 150 297 153 
rect 294 153 297 156 
rect 294 156 297 159 
rect 294 159 297 162 
rect 294 162 297 165 
rect 294 165 297 168 
rect 294 168 297 171 
rect 294 171 297 174 
rect 294 174 297 177 
rect 294 177 297 180 
rect 294 180 297 183 
rect 294 183 297 186 
rect 294 186 297 189 
rect 294 189 297 192 
rect 294 192 297 195 
rect 294 195 297 198 
rect 294 198 297 201 
rect 294 201 297 204 
rect 294 204 297 207 
rect 294 207 297 210 
rect 294 210 297 213 
rect 294 213 297 216 
rect 294 216 297 219 
rect 294 219 297 222 
rect 294 222 297 225 
rect 294 225 297 228 
rect 294 228 297 231 
rect 294 231 297 234 
rect 294 234 297 237 
rect 294 237 297 240 
rect 294 240 297 243 
rect 294 243 297 246 
rect 294 246 297 249 
rect 294 249 297 252 
rect 294 252 297 255 
rect 294 255 297 258 
rect 294 258 297 261 
rect 294 261 297 264 
rect 294 264 297 267 
rect 294 267 297 270 
rect 294 270 297 273 
rect 294 273 297 276 
rect 294 276 297 279 
rect 294 279 297 282 
rect 294 282 297 285 
rect 294 285 297 288 
rect 294 288 297 291 
rect 294 291 297 294 
rect 294 294 297 297 
rect 294 297 297 300 
rect 294 300 297 303 
rect 294 303 297 306 
rect 294 306 297 309 
rect 294 309 297 312 
rect 294 312 297 315 
rect 294 315 297 318 
rect 294 318 297 321 
rect 294 321 297 324 
rect 294 324 297 327 
rect 294 327 297 330 
rect 294 330 297 333 
rect 294 333 297 336 
rect 294 336 297 339 
rect 294 339 297 342 
rect 294 342 297 345 
rect 294 345 297 348 
rect 294 348 297 351 
rect 294 351 297 354 
rect 294 354 297 357 
rect 294 357 297 360 
rect 294 360 297 363 
rect 294 363 297 366 
rect 294 366 297 369 
rect 294 369 297 372 
rect 294 372 297 375 
rect 294 375 297 378 
rect 294 378 297 381 
rect 294 381 297 384 
rect 294 384 297 387 
rect 294 387 297 390 
rect 294 390 297 393 
rect 294 393 297 396 
rect 294 396 297 399 
rect 294 399 297 402 
rect 294 402 297 405 
rect 294 405 297 408 
rect 294 408 297 411 
rect 294 411 297 414 
rect 294 414 297 417 
rect 294 417 297 420 
rect 294 420 297 423 
rect 294 423 297 426 
rect 294 426 297 429 
rect 294 429 297 432 
rect 294 432 297 435 
rect 294 435 297 438 
rect 294 438 297 441 
rect 294 441 297 444 
rect 294 444 297 447 
rect 294 447 297 450 
rect 294 450 297 453 
rect 294 453 297 456 
rect 294 456 297 459 
rect 294 459 297 462 
rect 294 462 297 465 
rect 294 465 297 468 
rect 294 468 297 471 
rect 294 471 297 474 
rect 294 474 297 477 
rect 294 477 297 480 
rect 294 480 297 483 
rect 294 483 297 486 
rect 294 486 297 489 
rect 294 489 297 492 
rect 294 492 297 495 
rect 294 495 297 498 
rect 294 498 297 501 
rect 294 501 297 504 
rect 294 504 297 507 
rect 294 507 297 510 
rect 297 0 300 3 
rect 297 3 300 6 
rect 297 6 300 9 
rect 297 9 300 12 
rect 297 12 300 15 
rect 297 15 300 18 
rect 297 18 300 21 
rect 297 21 300 24 
rect 297 24 300 27 
rect 297 27 300 30 
rect 297 30 300 33 
rect 297 33 300 36 
rect 297 36 300 39 
rect 297 39 300 42 
rect 297 42 300 45 
rect 297 45 300 48 
rect 297 48 300 51 
rect 297 51 300 54 
rect 297 54 300 57 
rect 297 57 300 60 
rect 297 60 300 63 
rect 297 63 300 66 
rect 297 66 300 69 
rect 297 69 300 72 
rect 297 72 300 75 
rect 297 75 300 78 
rect 297 78 300 81 
rect 297 81 300 84 
rect 297 84 300 87 
rect 297 87 300 90 
rect 297 90 300 93 
rect 297 93 300 96 
rect 297 96 300 99 
rect 297 99 300 102 
rect 297 102 300 105 
rect 297 105 300 108 
rect 297 108 300 111 
rect 297 111 300 114 
rect 297 114 300 117 
rect 297 117 300 120 
rect 297 120 300 123 
rect 297 123 300 126 
rect 297 126 300 129 
rect 297 129 300 132 
rect 297 132 300 135 
rect 297 135 300 138 
rect 297 138 300 141 
rect 297 141 300 144 
rect 297 144 300 147 
rect 297 147 300 150 
rect 297 150 300 153 
rect 297 153 300 156 
rect 297 156 300 159 
rect 297 159 300 162 
rect 297 162 300 165 
rect 297 165 300 168 
rect 297 168 300 171 
rect 297 171 300 174 
rect 297 174 300 177 
rect 297 177 300 180 
rect 297 180 300 183 
rect 297 183 300 186 
rect 297 186 300 189 
rect 297 189 300 192 
rect 297 192 300 195 
rect 297 195 300 198 
rect 297 198 300 201 
rect 297 201 300 204 
rect 297 204 300 207 
rect 297 207 300 210 
rect 297 210 300 213 
rect 297 213 300 216 
rect 297 216 300 219 
rect 297 219 300 222 
rect 297 222 300 225 
rect 297 225 300 228 
rect 297 228 300 231 
rect 297 231 300 234 
rect 297 234 300 237 
rect 297 237 300 240 
rect 297 240 300 243 
rect 297 243 300 246 
rect 297 246 300 249 
rect 297 249 300 252 
rect 297 252 300 255 
rect 297 255 300 258 
rect 297 258 300 261 
rect 297 261 300 264 
rect 297 264 300 267 
rect 297 267 300 270 
rect 297 270 300 273 
rect 297 273 300 276 
rect 297 276 300 279 
rect 297 279 300 282 
rect 297 282 300 285 
rect 297 285 300 288 
rect 297 288 300 291 
rect 297 291 300 294 
rect 297 294 300 297 
rect 297 297 300 300 
rect 297 300 300 303 
rect 297 303 300 306 
rect 297 306 300 309 
rect 297 309 300 312 
rect 297 312 300 315 
rect 297 315 300 318 
rect 297 318 300 321 
rect 297 321 300 324 
rect 297 324 300 327 
rect 297 327 300 330 
rect 297 330 300 333 
rect 297 333 300 336 
rect 297 336 300 339 
rect 297 339 300 342 
rect 297 342 300 345 
rect 297 345 300 348 
rect 297 348 300 351 
rect 297 351 300 354 
rect 297 354 300 357 
rect 297 357 300 360 
rect 297 360 300 363 
rect 297 363 300 366 
rect 297 366 300 369 
rect 297 369 300 372 
rect 297 372 300 375 
rect 297 375 300 378 
rect 297 378 300 381 
rect 297 381 300 384 
rect 297 384 300 387 
rect 297 387 300 390 
rect 297 390 300 393 
rect 297 393 300 396 
rect 297 396 300 399 
rect 297 399 300 402 
rect 297 402 300 405 
rect 297 405 300 408 
rect 297 408 300 411 
rect 297 411 300 414 
rect 297 414 300 417 
rect 297 417 300 420 
rect 297 420 300 423 
rect 297 423 300 426 
rect 297 426 300 429 
rect 297 429 300 432 
rect 297 432 300 435 
rect 297 435 300 438 
rect 297 438 300 441 
rect 297 441 300 444 
rect 297 444 300 447 
rect 297 447 300 450 
rect 297 450 300 453 
rect 297 453 300 456 
rect 297 456 300 459 
rect 297 459 300 462 
rect 297 462 300 465 
rect 297 465 300 468 
rect 297 468 300 471 
rect 297 471 300 474 
rect 297 474 300 477 
rect 297 477 300 480 
rect 297 480 300 483 
rect 297 483 300 486 
rect 297 486 300 489 
rect 297 489 300 492 
rect 297 492 300 495 
rect 297 495 300 498 
rect 297 498 300 501 
rect 297 501 300 504 
rect 297 504 300 507 
rect 297 507 300 510 
rect 300 0 303 3 
rect 300 3 303 6 
rect 300 6 303 9 
rect 300 9 303 12 
rect 300 12 303 15 
rect 300 15 303 18 
rect 300 18 303 21 
rect 300 21 303 24 
rect 300 24 303 27 
rect 300 27 303 30 
rect 300 30 303 33 
rect 300 33 303 36 
rect 300 36 303 39 
rect 300 39 303 42 
rect 300 42 303 45 
rect 300 45 303 48 
rect 300 48 303 51 
rect 300 51 303 54 
rect 300 54 303 57 
rect 300 57 303 60 
rect 300 60 303 63 
rect 300 63 303 66 
rect 300 66 303 69 
rect 300 69 303 72 
rect 300 72 303 75 
rect 300 75 303 78 
rect 300 78 303 81 
rect 300 81 303 84 
rect 300 84 303 87 
rect 300 87 303 90 
rect 300 90 303 93 
rect 300 93 303 96 
rect 300 96 303 99 
rect 300 99 303 102 
rect 300 102 303 105 
rect 300 105 303 108 
rect 300 108 303 111 
rect 300 111 303 114 
rect 300 114 303 117 
rect 300 117 303 120 
rect 300 120 303 123 
rect 300 123 303 126 
rect 300 126 303 129 
rect 300 129 303 132 
rect 300 132 303 135 
rect 300 135 303 138 
rect 300 138 303 141 
rect 300 141 303 144 
rect 300 144 303 147 
rect 300 147 303 150 
rect 300 150 303 153 
rect 300 153 303 156 
rect 300 156 303 159 
rect 300 159 303 162 
rect 300 162 303 165 
rect 300 165 303 168 
rect 300 168 303 171 
rect 300 171 303 174 
rect 300 174 303 177 
rect 300 177 303 180 
rect 300 180 303 183 
rect 300 183 303 186 
rect 300 186 303 189 
rect 300 189 303 192 
rect 300 192 303 195 
rect 300 195 303 198 
rect 300 198 303 201 
rect 300 201 303 204 
rect 300 204 303 207 
rect 300 207 303 210 
rect 300 210 303 213 
rect 300 213 303 216 
rect 300 216 303 219 
rect 300 219 303 222 
rect 300 222 303 225 
rect 300 225 303 228 
rect 300 228 303 231 
rect 300 231 303 234 
rect 300 234 303 237 
rect 300 237 303 240 
rect 300 240 303 243 
rect 300 243 303 246 
rect 300 246 303 249 
rect 300 249 303 252 
rect 300 252 303 255 
rect 300 255 303 258 
rect 300 258 303 261 
rect 300 261 303 264 
rect 300 264 303 267 
rect 300 267 303 270 
rect 300 270 303 273 
rect 300 273 303 276 
rect 300 276 303 279 
rect 300 279 303 282 
rect 300 282 303 285 
rect 300 285 303 288 
rect 300 288 303 291 
rect 300 291 303 294 
rect 300 294 303 297 
rect 300 297 303 300 
rect 300 300 303 303 
rect 300 303 303 306 
rect 300 306 303 309 
rect 300 309 303 312 
rect 300 312 303 315 
rect 300 315 303 318 
rect 300 318 303 321 
rect 300 321 303 324 
rect 300 324 303 327 
rect 300 327 303 330 
rect 300 330 303 333 
rect 300 333 303 336 
rect 300 336 303 339 
rect 300 339 303 342 
rect 300 342 303 345 
rect 300 345 303 348 
rect 300 348 303 351 
rect 300 351 303 354 
rect 300 354 303 357 
rect 300 357 303 360 
rect 300 360 303 363 
rect 300 363 303 366 
rect 300 366 303 369 
rect 300 369 303 372 
rect 300 372 303 375 
rect 300 375 303 378 
rect 300 378 303 381 
rect 300 381 303 384 
rect 300 384 303 387 
rect 300 387 303 390 
rect 300 390 303 393 
rect 300 393 303 396 
rect 300 396 303 399 
rect 300 399 303 402 
rect 300 402 303 405 
rect 300 405 303 408 
rect 300 408 303 411 
rect 300 411 303 414 
rect 300 414 303 417 
rect 300 417 303 420 
rect 300 420 303 423 
rect 300 423 303 426 
rect 300 426 303 429 
rect 300 429 303 432 
rect 300 432 303 435 
rect 300 435 303 438 
rect 300 438 303 441 
rect 300 441 303 444 
rect 300 444 303 447 
rect 300 447 303 450 
rect 300 450 303 453 
rect 300 453 303 456 
rect 300 456 303 459 
rect 300 459 303 462 
rect 300 462 303 465 
rect 300 465 303 468 
rect 300 468 303 471 
rect 300 471 303 474 
rect 300 474 303 477 
rect 300 477 303 480 
rect 300 480 303 483 
rect 300 483 303 486 
rect 300 486 303 489 
rect 300 489 303 492 
rect 300 492 303 495 
rect 300 495 303 498 
rect 300 498 303 501 
rect 300 501 303 504 
rect 300 504 303 507 
rect 300 507 303 510 
rect 303 0 306 3 
rect 303 3 306 6 
rect 303 6 306 9 
rect 303 9 306 12 
rect 303 12 306 15 
rect 303 15 306 18 
rect 303 18 306 21 
rect 303 21 306 24 
rect 303 24 306 27 
rect 303 27 306 30 
rect 303 30 306 33 
rect 303 33 306 36 
rect 303 36 306 39 
rect 303 39 306 42 
rect 303 42 306 45 
rect 303 45 306 48 
rect 303 48 306 51 
rect 303 51 306 54 
rect 303 54 306 57 
rect 303 57 306 60 
rect 303 60 306 63 
rect 303 63 306 66 
rect 303 66 306 69 
rect 303 69 306 72 
rect 303 72 306 75 
rect 303 75 306 78 
rect 303 78 306 81 
rect 303 81 306 84 
rect 303 84 306 87 
rect 303 87 306 90 
rect 303 90 306 93 
rect 303 93 306 96 
rect 303 96 306 99 
rect 303 99 306 102 
rect 303 102 306 105 
rect 303 105 306 108 
rect 303 108 306 111 
rect 303 111 306 114 
rect 303 114 306 117 
rect 303 117 306 120 
rect 303 120 306 123 
rect 303 123 306 126 
rect 303 126 306 129 
rect 303 129 306 132 
rect 303 132 306 135 
rect 303 135 306 138 
rect 303 138 306 141 
rect 303 141 306 144 
rect 303 144 306 147 
rect 303 147 306 150 
rect 303 150 306 153 
rect 303 153 306 156 
rect 303 156 306 159 
rect 303 159 306 162 
rect 303 162 306 165 
rect 303 165 306 168 
rect 303 168 306 171 
rect 303 171 306 174 
rect 303 174 306 177 
rect 303 177 306 180 
rect 303 180 306 183 
rect 303 183 306 186 
rect 303 186 306 189 
rect 303 189 306 192 
rect 303 192 306 195 
rect 303 195 306 198 
rect 303 198 306 201 
rect 303 201 306 204 
rect 303 204 306 207 
rect 303 207 306 210 
rect 303 210 306 213 
rect 303 213 306 216 
rect 303 216 306 219 
rect 303 219 306 222 
rect 303 222 306 225 
rect 303 225 306 228 
rect 303 228 306 231 
rect 303 231 306 234 
rect 303 234 306 237 
rect 303 237 306 240 
rect 303 240 306 243 
rect 303 243 306 246 
rect 303 246 306 249 
rect 303 249 306 252 
rect 303 252 306 255 
rect 303 255 306 258 
rect 303 258 306 261 
rect 303 261 306 264 
rect 303 264 306 267 
rect 303 267 306 270 
rect 303 270 306 273 
rect 303 273 306 276 
rect 303 276 306 279 
rect 303 279 306 282 
rect 303 282 306 285 
rect 303 285 306 288 
rect 303 288 306 291 
rect 303 291 306 294 
rect 303 294 306 297 
rect 303 297 306 300 
rect 303 300 306 303 
rect 303 303 306 306 
rect 303 306 306 309 
rect 303 309 306 312 
rect 303 312 306 315 
rect 303 315 306 318 
rect 303 318 306 321 
rect 303 321 306 324 
rect 303 324 306 327 
rect 303 327 306 330 
rect 303 330 306 333 
rect 303 333 306 336 
rect 303 336 306 339 
rect 303 339 306 342 
rect 303 342 306 345 
rect 303 345 306 348 
rect 303 348 306 351 
rect 303 351 306 354 
rect 303 354 306 357 
rect 303 357 306 360 
rect 303 360 306 363 
rect 303 363 306 366 
rect 303 366 306 369 
rect 303 369 306 372 
rect 303 372 306 375 
rect 303 375 306 378 
rect 303 378 306 381 
rect 303 381 306 384 
rect 303 384 306 387 
rect 303 387 306 390 
rect 303 390 306 393 
rect 303 393 306 396 
rect 303 396 306 399 
rect 303 399 306 402 
rect 303 402 306 405 
rect 303 405 306 408 
rect 303 408 306 411 
rect 303 411 306 414 
rect 303 414 306 417 
rect 303 417 306 420 
rect 303 420 306 423 
rect 303 423 306 426 
rect 303 426 306 429 
rect 303 429 306 432 
rect 303 432 306 435 
rect 303 435 306 438 
rect 303 438 306 441 
rect 303 441 306 444 
rect 303 444 306 447 
rect 303 447 306 450 
rect 303 450 306 453 
rect 303 453 306 456 
rect 303 456 306 459 
rect 303 459 306 462 
rect 303 462 306 465 
rect 303 465 306 468 
rect 303 468 306 471 
rect 303 471 306 474 
rect 303 474 306 477 
rect 303 477 306 480 
rect 303 480 306 483 
rect 303 483 306 486 
rect 303 486 306 489 
rect 303 489 306 492 
rect 303 492 306 495 
rect 303 495 306 498 
rect 303 498 306 501 
rect 303 501 306 504 
rect 303 504 306 507 
rect 303 507 306 510 
rect 306 0 309 3 
rect 306 3 309 6 
rect 306 6 309 9 
rect 306 9 309 12 
rect 306 12 309 15 
rect 306 15 309 18 
rect 306 18 309 21 
rect 306 21 309 24 
rect 306 24 309 27 
rect 306 27 309 30 
rect 306 30 309 33 
rect 306 33 309 36 
rect 306 36 309 39 
rect 306 39 309 42 
rect 306 42 309 45 
rect 306 45 309 48 
rect 306 48 309 51 
rect 306 51 309 54 
rect 306 54 309 57 
rect 306 57 309 60 
rect 306 60 309 63 
rect 306 63 309 66 
rect 306 66 309 69 
rect 306 69 309 72 
rect 306 72 309 75 
rect 306 75 309 78 
rect 306 78 309 81 
rect 306 81 309 84 
rect 306 84 309 87 
rect 306 87 309 90 
rect 306 90 309 93 
rect 306 93 309 96 
rect 306 96 309 99 
rect 306 99 309 102 
rect 306 102 309 105 
rect 306 105 309 108 
rect 306 108 309 111 
rect 306 111 309 114 
rect 306 114 309 117 
rect 306 117 309 120 
rect 306 120 309 123 
rect 306 123 309 126 
rect 306 126 309 129 
rect 306 129 309 132 
rect 306 132 309 135 
rect 306 135 309 138 
rect 306 138 309 141 
rect 306 141 309 144 
rect 306 144 309 147 
rect 306 147 309 150 
rect 306 150 309 153 
rect 306 153 309 156 
rect 306 156 309 159 
rect 306 159 309 162 
rect 306 162 309 165 
rect 306 165 309 168 
rect 306 168 309 171 
rect 306 171 309 174 
rect 306 174 309 177 
rect 306 177 309 180 
rect 306 180 309 183 
rect 306 183 309 186 
rect 306 186 309 189 
rect 306 189 309 192 
rect 306 192 309 195 
rect 306 195 309 198 
rect 306 198 309 201 
rect 306 201 309 204 
rect 306 204 309 207 
rect 306 207 309 210 
rect 306 210 309 213 
rect 306 213 309 216 
rect 306 216 309 219 
rect 306 219 309 222 
rect 306 222 309 225 
rect 306 225 309 228 
rect 306 228 309 231 
rect 306 231 309 234 
rect 306 234 309 237 
rect 306 237 309 240 
rect 306 240 309 243 
rect 306 243 309 246 
rect 306 246 309 249 
rect 306 249 309 252 
rect 306 252 309 255 
rect 306 255 309 258 
rect 306 258 309 261 
rect 306 261 309 264 
rect 306 264 309 267 
rect 306 267 309 270 
rect 306 270 309 273 
rect 306 273 309 276 
rect 306 276 309 279 
rect 306 279 309 282 
rect 306 282 309 285 
rect 306 285 309 288 
rect 306 288 309 291 
rect 306 291 309 294 
rect 306 294 309 297 
rect 306 297 309 300 
rect 306 300 309 303 
rect 306 303 309 306 
rect 306 306 309 309 
rect 306 309 309 312 
rect 306 312 309 315 
rect 306 315 309 318 
rect 306 318 309 321 
rect 306 321 309 324 
rect 306 324 309 327 
rect 306 327 309 330 
rect 306 330 309 333 
rect 306 333 309 336 
rect 306 336 309 339 
rect 306 339 309 342 
rect 306 342 309 345 
rect 306 345 309 348 
rect 306 348 309 351 
rect 306 351 309 354 
rect 306 354 309 357 
rect 306 357 309 360 
rect 306 360 309 363 
rect 306 363 309 366 
rect 306 366 309 369 
rect 306 369 309 372 
rect 306 372 309 375 
rect 306 375 309 378 
rect 306 378 309 381 
rect 306 381 309 384 
rect 306 384 309 387 
rect 306 387 309 390 
rect 306 390 309 393 
rect 306 393 309 396 
rect 306 396 309 399 
rect 306 399 309 402 
rect 306 402 309 405 
rect 306 405 309 408 
rect 306 408 309 411 
rect 306 411 309 414 
rect 306 414 309 417 
rect 306 417 309 420 
rect 306 420 309 423 
rect 306 423 309 426 
rect 306 426 309 429 
rect 306 429 309 432 
rect 306 432 309 435 
rect 306 435 309 438 
rect 306 438 309 441 
rect 306 441 309 444 
rect 306 444 309 447 
rect 306 447 309 450 
rect 306 450 309 453 
rect 306 453 309 456 
rect 306 456 309 459 
rect 306 459 309 462 
rect 306 462 309 465 
rect 306 465 309 468 
rect 306 468 309 471 
rect 306 471 309 474 
rect 306 474 309 477 
rect 306 477 309 480 
rect 306 480 309 483 
rect 306 483 309 486 
rect 306 486 309 489 
rect 306 489 309 492 
rect 306 492 309 495 
rect 306 495 309 498 
rect 306 498 309 501 
rect 306 501 309 504 
rect 306 504 309 507 
rect 306 507 309 510 
rect 309 0 312 3 
rect 309 3 312 6 
rect 309 6 312 9 
rect 309 9 312 12 
rect 309 12 312 15 
rect 309 15 312 18 
rect 309 18 312 21 
rect 309 21 312 24 
rect 309 24 312 27 
rect 309 27 312 30 
rect 309 30 312 33 
rect 309 33 312 36 
rect 309 36 312 39 
rect 309 39 312 42 
rect 309 42 312 45 
rect 309 45 312 48 
rect 309 48 312 51 
rect 309 51 312 54 
rect 309 54 312 57 
rect 309 57 312 60 
rect 309 60 312 63 
rect 309 63 312 66 
rect 309 66 312 69 
rect 309 69 312 72 
rect 309 72 312 75 
rect 309 75 312 78 
rect 309 78 312 81 
rect 309 81 312 84 
rect 309 84 312 87 
rect 309 87 312 90 
rect 309 90 312 93 
rect 309 93 312 96 
rect 309 96 312 99 
rect 309 99 312 102 
rect 309 102 312 105 
rect 309 105 312 108 
rect 309 108 312 111 
rect 309 111 312 114 
rect 309 114 312 117 
rect 309 117 312 120 
rect 309 120 312 123 
rect 309 123 312 126 
rect 309 126 312 129 
rect 309 129 312 132 
rect 309 132 312 135 
rect 309 135 312 138 
rect 309 138 312 141 
rect 309 141 312 144 
rect 309 144 312 147 
rect 309 147 312 150 
rect 309 150 312 153 
rect 309 153 312 156 
rect 309 156 312 159 
rect 309 159 312 162 
rect 309 162 312 165 
rect 309 165 312 168 
rect 309 168 312 171 
rect 309 171 312 174 
rect 309 174 312 177 
rect 309 177 312 180 
rect 309 180 312 183 
rect 309 183 312 186 
rect 309 186 312 189 
rect 309 189 312 192 
rect 309 192 312 195 
rect 309 195 312 198 
rect 309 198 312 201 
rect 309 201 312 204 
rect 309 204 312 207 
rect 309 207 312 210 
rect 309 210 312 213 
rect 309 213 312 216 
rect 309 216 312 219 
rect 309 219 312 222 
rect 309 222 312 225 
rect 309 225 312 228 
rect 309 228 312 231 
rect 309 231 312 234 
rect 309 234 312 237 
rect 309 237 312 240 
rect 309 240 312 243 
rect 309 243 312 246 
rect 309 246 312 249 
rect 309 249 312 252 
rect 309 252 312 255 
rect 309 255 312 258 
rect 309 258 312 261 
rect 309 261 312 264 
rect 309 264 312 267 
rect 309 267 312 270 
rect 309 270 312 273 
rect 309 273 312 276 
rect 309 276 312 279 
rect 309 279 312 282 
rect 309 282 312 285 
rect 309 285 312 288 
rect 309 288 312 291 
rect 309 291 312 294 
rect 309 294 312 297 
rect 309 297 312 300 
rect 309 300 312 303 
rect 309 303 312 306 
rect 309 306 312 309 
rect 309 309 312 312 
rect 309 312 312 315 
rect 309 315 312 318 
rect 309 318 312 321 
rect 309 321 312 324 
rect 309 324 312 327 
rect 309 327 312 330 
rect 309 330 312 333 
rect 309 333 312 336 
rect 309 336 312 339 
rect 309 339 312 342 
rect 309 342 312 345 
rect 309 345 312 348 
rect 309 348 312 351 
rect 309 351 312 354 
rect 309 354 312 357 
rect 309 357 312 360 
rect 309 360 312 363 
rect 309 363 312 366 
rect 309 366 312 369 
rect 309 369 312 372 
rect 309 372 312 375 
rect 309 375 312 378 
rect 309 378 312 381 
rect 309 381 312 384 
rect 309 384 312 387 
rect 309 387 312 390 
rect 309 390 312 393 
rect 309 393 312 396 
rect 309 396 312 399 
rect 309 399 312 402 
rect 309 402 312 405 
rect 309 405 312 408 
rect 309 408 312 411 
rect 309 411 312 414 
rect 309 414 312 417 
rect 309 417 312 420 
rect 309 420 312 423 
rect 309 423 312 426 
rect 309 426 312 429 
rect 309 429 312 432 
rect 309 432 312 435 
rect 309 435 312 438 
rect 309 438 312 441 
rect 309 441 312 444 
rect 309 444 312 447 
rect 309 447 312 450 
rect 309 450 312 453 
rect 309 453 312 456 
rect 309 456 312 459 
rect 309 459 312 462 
rect 309 462 312 465 
rect 309 465 312 468 
rect 309 468 312 471 
rect 309 471 312 474 
rect 309 474 312 477 
rect 309 477 312 480 
rect 309 480 312 483 
rect 309 483 312 486 
rect 309 486 312 489 
rect 309 489 312 492 
rect 309 492 312 495 
rect 309 495 312 498 
rect 309 498 312 501 
rect 309 501 312 504 
rect 309 504 312 507 
rect 309 507 312 510 
rect 312 0 315 3 
rect 312 3 315 6 
rect 312 6 315 9 
rect 312 9 315 12 
rect 312 12 315 15 
rect 312 15 315 18 
rect 312 18 315 21 
rect 312 21 315 24 
rect 312 24 315 27 
rect 312 27 315 30 
rect 312 30 315 33 
rect 312 33 315 36 
rect 312 36 315 39 
rect 312 39 315 42 
rect 312 42 315 45 
rect 312 45 315 48 
rect 312 48 315 51 
rect 312 51 315 54 
rect 312 54 315 57 
rect 312 57 315 60 
rect 312 60 315 63 
rect 312 63 315 66 
rect 312 66 315 69 
rect 312 69 315 72 
rect 312 72 315 75 
rect 312 75 315 78 
rect 312 78 315 81 
rect 312 81 315 84 
rect 312 84 315 87 
rect 312 87 315 90 
rect 312 90 315 93 
rect 312 93 315 96 
rect 312 96 315 99 
rect 312 99 315 102 
rect 312 102 315 105 
rect 312 105 315 108 
rect 312 108 315 111 
rect 312 111 315 114 
rect 312 114 315 117 
rect 312 117 315 120 
rect 312 120 315 123 
rect 312 123 315 126 
rect 312 126 315 129 
rect 312 129 315 132 
rect 312 132 315 135 
rect 312 135 315 138 
rect 312 138 315 141 
rect 312 141 315 144 
rect 312 144 315 147 
rect 312 147 315 150 
rect 312 150 315 153 
rect 312 153 315 156 
rect 312 156 315 159 
rect 312 159 315 162 
rect 312 162 315 165 
rect 312 165 315 168 
rect 312 168 315 171 
rect 312 171 315 174 
rect 312 174 315 177 
rect 312 177 315 180 
rect 312 180 315 183 
rect 312 183 315 186 
rect 312 186 315 189 
rect 312 189 315 192 
rect 312 192 315 195 
rect 312 195 315 198 
rect 312 198 315 201 
rect 312 201 315 204 
rect 312 204 315 207 
rect 312 207 315 210 
rect 312 210 315 213 
rect 312 213 315 216 
rect 312 216 315 219 
rect 312 219 315 222 
rect 312 222 315 225 
rect 312 225 315 228 
rect 312 228 315 231 
rect 312 231 315 234 
rect 312 234 315 237 
rect 312 237 315 240 
rect 312 240 315 243 
rect 312 243 315 246 
rect 312 246 315 249 
rect 312 249 315 252 
rect 312 252 315 255 
rect 312 255 315 258 
rect 312 258 315 261 
rect 312 261 315 264 
rect 312 264 315 267 
rect 312 267 315 270 
rect 312 270 315 273 
rect 312 273 315 276 
rect 312 276 315 279 
rect 312 279 315 282 
rect 312 282 315 285 
rect 312 285 315 288 
rect 312 288 315 291 
rect 312 291 315 294 
rect 312 294 315 297 
rect 312 297 315 300 
rect 312 300 315 303 
rect 312 303 315 306 
rect 312 306 315 309 
rect 312 309 315 312 
rect 312 312 315 315 
rect 312 315 315 318 
rect 312 318 315 321 
rect 312 321 315 324 
rect 312 324 315 327 
rect 312 327 315 330 
rect 312 330 315 333 
rect 312 333 315 336 
rect 312 336 315 339 
rect 312 339 315 342 
rect 312 342 315 345 
rect 312 345 315 348 
rect 312 348 315 351 
rect 312 351 315 354 
rect 312 354 315 357 
rect 312 357 315 360 
rect 312 360 315 363 
rect 312 363 315 366 
rect 312 366 315 369 
rect 312 369 315 372 
rect 312 372 315 375 
rect 312 375 315 378 
rect 312 378 315 381 
rect 312 381 315 384 
rect 312 384 315 387 
rect 312 387 315 390 
rect 312 390 315 393 
rect 312 393 315 396 
rect 312 396 315 399 
rect 312 399 315 402 
rect 312 402 315 405 
rect 312 405 315 408 
rect 312 408 315 411 
rect 312 411 315 414 
rect 312 414 315 417 
rect 312 417 315 420 
rect 312 420 315 423 
rect 312 423 315 426 
rect 312 426 315 429 
rect 312 429 315 432 
rect 312 432 315 435 
rect 312 435 315 438 
rect 312 438 315 441 
rect 312 441 315 444 
rect 312 444 315 447 
rect 312 447 315 450 
rect 312 450 315 453 
rect 312 453 315 456 
rect 312 456 315 459 
rect 312 459 315 462 
rect 312 462 315 465 
rect 312 465 315 468 
rect 312 468 315 471 
rect 312 471 315 474 
rect 312 474 315 477 
rect 312 477 315 480 
rect 312 480 315 483 
rect 312 483 315 486 
rect 312 486 315 489 
rect 312 489 315 492 
rect 312 492 315 495 
rect 312 495 315 498 
rect 312 498 315 501 
rect 312 501 315 504 
rect 312 504 315 507 
rect 312 507 315 510 
rect 315 0 318 3 
rect 315 3 318 6 
rect 315 6 318 9 
rect 315 9 318 12 
rect 315 12 318 15 
rect 315 15 318 18 
rect 315 18 318 21 
rect 315 21 318 24 
rect 315 24 318 27 
rect 315 27 318 30 
rect 315 30 318 33 
rect 315 33 318 36 
rect 315 36 318 39 
rect 315 39 318 42 
rect 315 42 318 45 
rect 315 45 318 48 
rect 315 48 318 51 
rect 315 51 318 54 
rect 315 54 318 57 
rect 315 57 318 60 
rect 315 60 318 63 
rect 315 63 318 66 
rect 315 66 318 69 
rect 315 69 318 72 
rect 315 72 318 75 
rect 315 75 318 78 
rect 315 78 318 81 
rect 315 81 318 84 
rect 315 84 318 87 
rect 315 87 318 90 
rect 315 90 318 93 
rect 315 93 318 96 
rect 315 96 318 99 
rect 315 99 318 102 
rect 315 102 318 105 
rect 315 105 318 108 
rect 315 108 318 111 
rect 315 111 318 114 
rect 315 114 318 117 
rect 315 117 318 120 
rect 315 120 318 123 
rect 315 123 318 126 
rect 315 126 318 129 
rect 315 129 318 132 
rect 315 132 318 135 
rect 315 135 318 138 
rect 315 138 318 141 
rect 315 141 318 144 
rect 315 144 318 147 
rect 315 147 318 150 
rect 315 150 318 153 
rect 315 153 318 156 
rect 315 156 318 159 
rect 315 159 318 162 
rect 315 162 318 165 
rect 315 165 318 168 
rect 315 168 318 171 
rect 315 171 318 174 
rect 315 174 318 177 
rect 315 177 318 180 
rect 315 180 318 183 
rect 315 183 318 186 
rect 315 186 318 189 
rect 315 189 318 192 
rect 315 192 318 195 
rect 315 195 318 198 
rect 315 198 318 201 
rect 315 201 318 204 
rect 315 204 318 207 
rect 315 207 318 210 
rect 315 210 318 213 
rect 315 213 318 216 
rect 315 216 318 219 
rect 315 219 318 222 
rect 315 222 318 225 
rect 315 225 318 228 
rect 315 228 318 231 
rect 315 231 318 234 
rect 315 234 318 237 
rect 315 237 318 240 
rect 315 240 318 243 
rect 315 243 318 246 
rect 315 246 318 249 
rect 315 249 318 252 
rect 315 252 318 255 
rect 315 255 318 258 
rect 315 258 318 261 
rect 315 261 318 264 
rect 315 264 318 267 
rect 315 267 318 270 
rect 315 270 318 273 
rect 315 273 318 276 
rect 315 276 318 279 
rect 315 279 318 282 
rect 315 282 318 285 
rect 315 285 318 288 
rect 315 288 318 291 
rect 315 291 318 294 
rect 315 294 318 297 
rect 315 297 318 300 
rect 315 300 318 303 
rect 315 303 318 306 
rect 315 306 318 309 
rect 315 309 318 312 
rect 315 312 318 315 
rect 315 315 318 318 
rect 315 318 318 321 
rect 315 321 318 324 
rect 315 324 318 327 
rect 315 327 318 330 
rect 315 330 318 333 
rect 315 333 318 336 
rect 315 336 318 339 
rect 315 339 318 342 
rect 315 342 318 345 
rect 315 345 318 348 
rect 315 348 318 351 
rect 315 351 318 354 
rect 315 354 318 357 
rect 315 357 318 360 
rect 315 360 318 363 
rect 315 363 318 366 
rect 315 366 318 369 
rect 315 369 318 372 
rect 315 372 318 375 
rect 315 375 318 378 
rect 315 378 318 381 
rect 315 381 318 384 
rect 315 384 318 387 
rect 315 387 318 390 
rect 315 390 318 393 
rect 315 393 318 396 
rect 315 396 318 399 
rect 315 399 318 402 
rect 315 402 318 405 
rect 315 405 318 408 
rect 315 408 318 411 
rect 315 411 318 414 
rect 315 414 318 417 
rect 315 417 318 420 
rect 315 420 318 423 
rect 315 423 318 426 
rect 315 426 318 429 
rect 315 429 318 432 
rect 315 432 318 435 
rect 315 435 318 438 
rect 315 438 318 441 
rect 315 441 318 444 
rect 315 444 318 447 
rect 315 447 318 450 
rect 315 450 318 453 
rect 315 453 318 456 
rect 315 456 318 459 
rect 315 459 318 462 
rect 315 462 318 465 
rect 315 465 318 468 
rect 315 468 318 471 
rect 315 471 318 474 
rect 315 474 318 477 
rect 315 477 318 480 
rect 315 480 318 483 
rect 315 483 318 486 
rect 315 486 318 489 
rect 315 489 318 492 
rect 315 492 318 495 
rect 315 495 318 498 
rect 315 498 318 501 
rect 315 501 318 504 
rect 315 504 318 507 
rect 315 507 318 510 
rect 318 0 321 3 
rect 318 3 321 6 
rect 318 6 321 9 
rect 318 9 321 12 
rect 318 12 321 15 
rect 318 15 321 18 
rect 318 18 321 21 
rect 318 21 321 24 
rect 318 24 321 27 
rect 318 27 321 30 
rect 318 30 321 33 
rect 318 33 321 36 
rect 318 36 321 39 
rect 318 39 321 42 
rect 318 42 321 45 
rect 318 45 321 48 
rect 318 48 321 51 
rect 318 51 321 54 
rect 318 54 321 57 
rect 318 57 321 60 
rect 318 60 321 63 
rect 318 63 321 66 
rect 318 66 321 69 
rect 318 69 321 72 
rect 318 72 321 75 
rect 318 75 321 78 
rect 318 78 321 81 
rect 318 81 321 84 
rect 318 84 321 87 
rect 318 87 321 90 
rect 318 90 321 93 
rect 318 93 321 96 
rect 318 96 321 99 
rect 318 99 321 102 
rect 318 102 321 105 
rect 318 105 321 108 
rect 318 108 321 111 
rect 318 111 321 114 
rect 318 114 321 117 
rect 318 117 321 120 
rect 318 120 321 123 
rect 318 123 321 126 
rect 318 126 321 129 
rect 318 129 321 132 
rect 318 132 321 135 
rect 318 135 321 138 
rect 318 138 321 141 
rect 318 141 321 144 
rect 318 144 321 147 
rect 318 147 321 150 
rect 318 150 321 153 
rect 318 153 321 156 
rect 318 156 321 159 
rect 318 159 321 162 
rect 318 162 321 165 
rect 318 165 321 168 
rect 318 168 321 171 
rect 318 171 321 174 
rect 318 174 321 177 
rect 318 177 321 180 
rect 318 180 321 183 
rect 318 183 321 186 
rect 318 189 321 192 
rect 318 192 321 195 
rect 318 195 321 198 
rect 318 198 321 201 
rect 318 201 321 204 
rect 318 204 321 207 
rect 318 207 321 210 
rect 318 210 321 213 
rect 318 213 321 216 
rect 318 216 321 219 
rect 318 219 321 222 
rect 318 222 321 225 
rect 318 225 321 228 
rect 318 228 321 231 
rect 318 231 321 234 
rect 318 237 321 240 
rect 318 240 321 243 
rect 318 243 321 246 
rect 318 246 321 249 
rect 318 249 321 252 
rect 318 252 321 255 
rect 318 255 321 258 
rect 318 258 321 261 
rect 318 261 321 264 
rect 318 264 321 267 
rect 318 267 321 270 
rect 318 270 321 273 
rect 318 273 321 276 
rect 318 276 321 279 
rect 318 279 321 282 
rect 318 282 321 285 
rect 318 285 321 288 
rect 318 288 321 291 
rect 318 291 321 294 
rect 318 294 321 297 
rect 318 297 321 300 
rect 318 300 321 303 
rect 318 303 321 306 
rect 318 306 321 309 
rect 318 309 321 312 
rect 318 312 321 315 
rect 318 315 321 318 
rect 318 318 321 321 
rect 318 321 321 324 
rect 318 324 321 327 
rect 318 327 321 330 
rect 318 333 321 336 
rect 318 336 321 339 
rect 318 339 321 342 
rect 318 342 321 345 
rect 318 345 321 348 
rect 318 348 321 351 
rect 318 351 321 354 
rect 318 354 321 357 
rect 318 357 321 360 
rect 318 360 321 363 
rect 318 363 321 366 
rect 318 366 321 369 
rect 318 372 321 375 
rect 318 375 321 378 
rect 318 381 321 384 
rect 318 384 321 387 
rect 318 387 321 390 
rect 318 390 321 393 
rect 318 393 321 396 
rect 318 396 321 399 
rect 318 399 321 402 
rect 318 402 321 405 
rect 318 405 321 408 
rect 318 408 321 411 
rect 318 411 321 414 
rect 318 414 321 417 
rect 318 417 321 420 
rect 318 420 321 423 
rect 318 423 321 426 
rect 318 426 321 429 
rect 318 429 321 432 
rect 318 432 321 435 
rect 318 435 321 438 
rect 318 438 321 441 
rect 318 441 321 444 
rect 318 444 321 447 
rect 318 447 321 450 
rect 318 450 321 453 
rect 318 453 321 456 
rect 318 456 321 459 
rect 318 459 321 462 
rect 318 462 321 465 
rect 318 465 321 468 
rect 318 468 321 471 
rect 318 471 321 474 
rect 318 474 321 477 
rect 318 477 321 480 
rect 318 480 321 483 
rect 318 483 321 486 
rect 318 486 321 489 
rect 318 489 321 492 
rect 318 492 321 495 
rect 318 495 321 498 
rect 318 498 321 501 
rect 318 501 321 504 
rect 318 504 321 507 
rect 318 507 321 510 
rect 321 0 324 3 
rect 321 3 324 6 
rect 321 6 324 9 
rect 321 9 324 12 
rect 321 12 324 15 
rect 321 15 324 18 
rect 321 18 324 21 
rect 321 21 324 24 
rect 321 24 324 27 
rect 321 27 324 30 
rect 321 30 324 33 
rect 321 33 324 36 
rect 321 36 324 39 
rect 321 39 324 42 
rect 321 42 324 45 
rect 321 45 324 48 
rect 321 48 324 51 
rect 321 51 324 54 
rect 321 54 324 57 
rect 321 57 324 60 
rect 321 60 324 63 
rect 321 63 324 66 
rect 321 66 324 69 
rect 321 69 324 72 
rect 321 72 324 75 
rect 321 75 324 78 
rect 321 78 324 81 
rect 321 81 324 84 
rect 321 84 324 87 
rect 321 87 324 90 
rect 321 90 324 93 
rect 321 93 324 96 
rect 321 96 324 99 
rect 321 99 324 102 
rect 321 102 324 105 
rect 321 105 324 108 
rect 321 108 324 111 
rect 321 111 324 114 
rect 321 114 324 117 
rect 321 117 324 120 
rect 321 120 324 123 
rect 321 123 324 126 
rect 321 126 324 129 
rect 321 129 324 132 
rect 321 132 324 135 
rect 321 135 324 138 
rect 321 138 324 141 
rect 321 141 324 144 
rect 321 144 324 147 
rect 321 147 324 150 
rect 321 150 324 153 
rect 321 153 324 156 
rect 321 156 324 159 
rect 321 159 324 162 
rect 321 162 324 165 
rect 321 165 324 168 
rect 321 168 324 171 
rect 321 171 324 174 
rect 321 174 324 177 
rect 321 177 324 180 
rect 321 180 324 183 
rect 321 183 324 186 
rect 321 186 324 189 
rect 321 189 324 192 
rect 321 192 324 195 
rect 321 195 324 198 
rect 321 198 324 201 
rect 321 201 324 204 
rect 321 204 324 207 
rect 321 207 324 210 
rect 321 210 324 213 
rect 321 213 324 216 
rect 321 216 324 219 
rect 321 219 324 222 
rect 321 222 324 225 
rect 321 225 324 228 
rect 321 228 324 231 
rect 321 231 324 234 
rect 321 234 324 237 
rect 321 237 324 240 
rect 321 240 324 243 
rect 321 243 324 246 
rect 321 246 324 249 
rect 321 249 324 252 
rect 321 252 324 255 
rect 321 255 324 258 
rect 321 258 324 261 
rect 321 261 324 264 
rect 321 264 324 267 
rect 321 267 324 270 
rect 321 270 324 273 
rect 321 273 324 276 
rect 321 276 324 279 
rect 321 279 324 282 
rect 321 282 324 285 
rect 321 285 324 288 
rect 321 288 324 291 
rect 321 291 324 294 
rect 321 294 324 297 
rect 321 297 324 300 
rect 321 300 324 303 
rect 321 303 324 306 
rect 321 306 324 309 
rect 321 309 324 312 
rect 321 312 324 315 
rect 321 315 324 318 
rect 321 318 324 321 
rect 321 321 324 324 
rect 321 324 324 327 
rect 321 327 324 330 
rect 321 330 324 333 
rect 321 333 324 336 
rect 321 336 324 339 
rect 321 339 324 342 
rect 321 342 324 345 
rect 321 345 324 348 
rect 321 348 324 351 
rect 321 351 324 354 
rect 321 354 324 357 
rect 321 357 324 360 
rect 321 360 324 363 
rect 321 363 324 366 
rect 321 366 324 369 
rect 321 369 324 372 
rect 321 372 324 375 
rect 321 375 324 378 
rect 321 378 324 381 
rect 321 381 324 384 
rect 321 384 324 387 
rect 321 387 324 390 
rect 321 390 324 393 
rect 321 393 324 396 
rect 321 396 324 399 
rect 321 399 324 402 
rect 321 402 324 405 
rect 321 405 324 408 
rect 321 408 324 411 
rect 321 411 324 414 
rect 321 414 324 417 
rect 321 417 324 420 
rect 321 420 324 423 
rect 321 423 324 426 
rect 321 426 324 429 
rect 321 429 324 432 
rect 321 432 324 435 
rect 321 435 324 438 
rect 321 438 324 441 
rect 321 441 324 444 
rect 321 444 324 447 
rect 321 447 324 450 
rect 321 450 324 453 
rect 321 453 324 456 
rect 321 456 324 459 
rect 321 459 324 462 
rect 321 462 324 465 
rect 321 465 324 468 
rect 321 468 324 471 
rect 321 471 324 474 
rect 321 474 324 477 
rect 321 477 324 480 
rect 321 480 324 483 
rect 321 483 324 486 
rect 321 486 324 489 
rect 321 489 324 492 
rect 321 492 324 495 
rect 321 495 324 498 
rect 321 498 324 501 
rect 321 501 324 504 
rect 321 504 324 507 
rect 321 507 324 510 
rect 324 0 327 3 
rect 324 3 327 6 
rect 324 6 327 9 
rect 324 9 327 12 
rect 324 12 327 15 
rect 324 15 327 18 
rect 324 18 327 21 
rect 324 21 327 24 
rect 324 24 327 27 
rect 324 27 327 30 
rect 324 30 327 33 
rect 324 33 327 36 
rect 324 36 327 39 
rect 324 39 327 42 
rect 324 42 327 45 
rect 324 45 327 48 
rect 324 48 327 51 
rect 324 51 327 54 
rect 324 54 327 57 
rect 324 57 327 60 
rect 324 60 327 63 
rect 324 63 327 66 
rect 324 66 327 69 
rect 324 69 327 72 
rect 324 72 327 75 
rect 324 75 327 78 
rect 324 78 327 81 
rect 324 81 327 84 
rect 324 84 327 87 
rect 324 87 327 90 
rect 324 90 327 93 
rect 324 93 327 96 
rect 324 96 327 99 
rect 324 99 327 102 
rect 324 102 327 105 
rect 324 105 327 108 
rect 324 108 327 111 
rect 324 111 327 114 
rect 324 114 327 117 
rect 324 117 327 120 
rect 324 120 327 123 
rect 324 123 327 126 
rect 324 126 327 129 
rect 324 129 327 132 
rect 324 132 327 135 
rect 324 135 327 138 
rect 324 138 327 141 
rect 324 141 327 144 
rect 324 144 327 147 
rect 324 147 327 150 
rect 324 150 327 153 
rect 324 153 327 156 
rect 324 156 327 159 
rect 324 159 327 162 
rect 324 162 327 165 
rect 324 165 327 168 
rect 324 168 327 171 
rect 324 171 327 174 
rect 324 174 327 177 
rect 324 177 327 180 
rect 324 180 327 183 
rect 324 183 327 186 
rect 324 186 327 189 
rect 324 189 327 192 
rect 324 192 327 195 
rect 324 195 327 198 
rect 324 198 327 201 
rect 324 201 327 204 
rect 324 204 327 207 
rect 324 207 327 210 
rect 324 210 327 213 
rect 324 213 327 216 
rect 324 216 327 219 
rect 324 219 327 222 
rect 324 222 327 225 
rect 324 225 327 228 
rect 324 228 327 231 
rect 324 231 327 234 
rect 324 234 327 237 
rect 324 237 327 240 
rect 324 240 327 243 
rect 324 243 327 246 
rect 324 246 327 249 
rect 324 249 327 252 
rect 324 252 327 255 
rect 324 255 327 258 
rect 324 258 327 261 
rect 324 261 327 264 
rect 324 264 327 267 
rect 324 267 327 270 
rect 324 270 327 273 
rect 324 273 327 276 
rect 324 276 327 279 
rect 324 279 327 282 
rect 324 282 327 285 
rect 324 285 327 288 
rect 324 288 327 291 
rect 324 291 327 294 
rect 324 294 327 297 
rect 324 297 327 300 
rect 324 300 327 303 
rect 324 303 327 306 
rect 324 306 327 309 
rect 324 309 327 312 
rect 324 312 327 315 
rect 324 315 327 318 
rect 324 318 327 321 
rect 324 321 327 324 
rect 324 324 327 327 
rect 324 327 327 330 
rect 324 330 327 333 
rect 324 333 327 336 
rect 324 336 327 339 
rect 324 339 327 342 
rect 324 342 327 345 
rect 324 345 327 348 
rect 324 348 327 351 
rect 324 351 327 354 
rect 324 354 327 357 
rect 324 357 327 360 
rect 324 360 327 363 
rect 324 363 327 366 
rect 324 366 327 369 
rect 324 369 327 372 
rect 324 372 327 375 
rect 324 375 327 378 
rect 324 378 327 381 
rect 324 381 327 384 
rect 324 384 327 387 
rect 324 387 327 390 
rect 324 390 327 393 
rect 324 393 327 396 
rect 324 396 327 399 
rect 324 399 327 402 
rect 324 402 327 405 
rect 324 405 327 408 
rect 324 408 327 411 
rect 324 411 327 414 
rect 324 414 327 417 
rect 324 417 327 420 
rect 324 420 327 423 
rect 324 423 327 426 
rect 324 426 327 429 
rect 324 429 327 432 
rect 324 432 327 435 
rect 324 435 327 438 
rect 324 438 327 441 
rect 324 441 327 444 
rect 324 444 327 447 
rect 324 447 327 450 
rect 324 450 327 453 
rect 324 453 327 456 
rect 324 456 327 459 
rect 324 459 327 462 
rect 324 462 327 465 
rect 324 465 327 468 
rect 324 468 327 471 
rect 324 471 327 474 
rect 324 474 327 477 
rect 324 477 327 480 
rect 324 480 327 483 
rect 324 483 327 486 
rect 324 486 327 489 
rect 324 489 327 492 
rect 324 492 327 495 
rect 324 495 327 498 
rect 324 498 327 501 
rect 324 501 327 504 
rect 324 504 327 507 
rect 324 507 327 510 
rect 327 0 330 3 
rect 327 3 330 6 
rect 327 6 330 9 
rect 327 9 330 12 
rect 327 12 330 15 
rect 327 15 330 18 
rect 327 18 330 21 
rect 327 21 330 24 
rect 327 24 330 27 
rect 327 27 330 30 
rect 327 30 330 33 
rect 327 33 330 36 
rect 327 36 330 39 
rect 327 39 330 42 
rect 327 42 330 45 
rect 327 45 330 48 
rect 327 48 330 51 
rect 327 51 330 54 
rect 327 54 330 57 
rect 327 57 330 60 
rect 327 60 330 63 
rect 327 63 330 66 
rect 327 66 330 69 
rect 327 69 330 72 
rect 327 72 330 75 
rect 327 75 330 78 
rect 327 78 330 81 
rect 327 81 330 84 
rect 327 84 330 87 
rect 327 87 330 90 
rect 327 90 330 93 
rect 327 93 330 96 
rect 327 96 330 99 
rect 327 99 330 102 
rect 327 102 330 105 
rect 327 105 330 108 
rect 327 108 330 111 
rect 327 111 330 114 
rect 327 114 330 117 
rect 327 117 330 120 
rect 327 120 330 123 
rect 327 123 330 126 
rect 327 126 330 129 
rect 327 129 330 132 
rect 327 132 330 135 
rect 327 135 330 138 
rect 327 138 330 141 
rect 327 141 330 144 
rect 327 144 330 147 
rect 327 147 330 150 
rect 327 150 330 153 
rect 327 153 330 156 
rect 327 156 330 159 
rect 327 159 330 162 
rect 327 162 330 165 
rect 327 165 330 168 
rect 327 168 330 171 
rect 327 171 330 174 
rect 327 174 330 177 
rect 327 177 330 180 
rect 327 180 330 183 
rect 327 183 330 186 
rect 327 186 330 189 
rect 327 189 330 192 
rect 327 192 330 195 
rect 327 195 330 198 
rect 327 198 330 201 
rect 327 201 330 204 
rect 327 204 330 207 
rect 327 207 330 210 
rect 327 210 330 213 
rect 327 213 330 216 
rect 327 216 330 219 
rect 327 219 330 222 
rect 327 222 330 225 
rect 327 225 330 228 
rect 327 228 330 231 
rect 327 231 330 234 
rect 327 234 330 237 
rect 327 237 330 240 
rect 327 240 330 243 
rect 327 243 330 246 
rect 327 246 330 249 
rect 327 249 330 252 
rect 327 252 330 255 
rect 327 255 330 258 
rect 327 258 330 261 
rect 327 261 330 264 
rect 327 264 330 267 
rect 327 267 330 270 
rect 327 270 330 273 
rect 327 273 330 276 
rect 327 276 330 279 
rect 327 279 330 282 
rect 327 282 330 285 
rect 327 285 330 288 
rect 327 288 330 291 
rect 327 291 330 294 
rect 327 294 330 297 
rect 327 297 330 300 
rect 327 300 330 303 
rect 327 303 330 306 
rect 327 306 330 309 
rect 327 309 330 312 
rect 327 312 330 315 
rect 327 315 330 318 
rect 327 318 330 321 
rect 327 321 330 324 
rect 327 324 330 327 
rect 327 327 330 330 
rect 327 330 330 333 
rect 327 333 330 336 
rect 327 336 330 339 
rect 327 339 330 342 
rect 327 342 330 345 
rect 327 345 330 348 
rect 327 348 330 351 
rect 327 351 330 354 
rect 327 354 330 357 
rect 327 357 330 360 
rect 327 360 330 363 
rect 327 363 330 366 
rect 327 366 330 369 
rect 327 369 330 372 
rect 327 372 330 375 
rect 327 375 330 378 
rect 327 378 330 381 
rect 327 381 330 384 
rect 327 384 330 387 
rect 327 387 330 390 
rect 327 390 330 393 
rect 327 393 330 396 
rect 327 396 330 399 
rect 327 399 330 402 
rect 327 402 330 405 
rect 327 405 330 408 
rect 327 408 330 411 
rect 327 411 330 414 
rect 327 414 330 417 
rect 327 417 330 420 
rect 327 420 330 423 
rect 327 423 330 426 
rect 327 426 330 429 
rect 327 429 330 432 
rect 327 432 330 435 
rect 327 435 330 438 
rect 327 438 330 441 
rect 327 441 330 444 
rect 327 444 330 447 
rect 327 447 330 450 
rect 327 450 330 453 
rect 327 453 330 456 
rect 327 456 330 459 
rect 327 459 330 462 
rect 327 462 330 465 
rect 327 465 330 468 
rect 327 468 330 471 
rect 327 471 330 474 
rect 327 474 330 477 
rect 327 477 330 480 
rect 327 480 330 483 
rect 327 483 330 486 
rect 327 486 330 489 
rect 327 489 330 492 
rect 327 492 330 495 
rect 327 495 330 498 
rect 327 498 330 501 
rect 327 501 330 504 
rect 327 504 330 507 
rect 327 507 330 510 
rect 330 0 333 3 
rect 330 3 333 6 
rect 330 6 333 9 
rect 330 9 333 12 
rect 330 12 333 15 
rect 330 15 333 18 
rect 330 18 333 21 
rect 330 21 333 24 
rect 330 24 333 27 
rect 330 27 333 30 
rect 330 30 333 33 
rect 330 33 333 36 
rect 330 36 333 39 
rect 330 39 333 42 
rect 330 42 333 45 
rect 330 45 333 48 
rect 330 48 333 51 
rect 330 51 333 54 
rect 330 54 333 57 
rect 330 57 333 60 
rect 330 60 333 63 
rect 330 63 333 66 
rect 330 66 333 69 
rect 330 69 333 72 
rect 330 72 333 75 
rect 330 75 333 78 
rect 330 78 333 81 
rect 330 81 333 84 
rect 330 84 333 87 
rect 330 87 333 90 
rect 330 90 333 93 
rect 330 93 333 96 
rect 330 96 333 99 
rect 330 99 333 102 
rect 330 102 333 105 
rect 330 105 333 108 
rect 330 108 333 111 
rect 330 111 333 114 
rect 330 114 333 117 
rect 330 117 333 120 
rect 330 120 333 123 
rect 330 123 333 126 
rect 330 126 333 129 
rect 330 129 333 132 
rect 330 132 333 135 
rect 330 135 333 138 
rect 330 138 333 141 
rect 330 141 333 144 
rect 330 144 333 147 
rect 330 147 333 150 
rect 330 150 333 153 
rect 330 153 333 156 
rect 330 156 333 159 
rect 330 159 333 162 
rect 330 162 333 165 
rect 330 165 333 168 
rect 330 168 333 171 
rect 330 171 333 174 
rect 330 174 333 177 
rect 330 177 333 180 
rect 330 180 333 183 
rect 330 183 333 186 
rect 330 186 333 189 
rect 330 189 333 192 
rect 330 192 333 195 
rect 330 195 333 198 
rect 330 198 333 201 
rect 330 201 333 204 
rect 330 204 333 207 
rect 330 207 333 210 
rect 330 210 333 213 
rect 330 213 333 216 
rect 330 216 333 219 
rect 330 219 333 222 
rect 330 222 333 225 
rect 330 225 333 228 
rect 330 228 333 231 
rect 330 231 333 234 
rect 330 234 333 237 
rect 330 237 333 240 
rect 330 240 333 243 
rect 330 243 333 246 
rect 330 246 333 249 
rect 330 249 333 252 
rect 330 252 333 255 
rect 330 255 333 258 
rect 330 258 333 261 
rect 330 261 333 264 
rect 330 264 333 267 
rect 330 267 333 270 
rect 330 270 333 273 
rect 330 273 333 276 
rect 330 276 333 279 
rect 330 279 333 282 
rect 330 282 333 285 
rect 330 285 333 288 
rect 330 288 333 291 
rect 330 291 333 294 
rect 330 294 333 297 
rect 330 297 333 300 
rect 330 300 333 303 
rect 330 303 333 306 
rect 330 306 333 309 
rect 330 309 333 312 
rect 330 312 333 315 
rect 330 315 333 318 
rect 330 318 333 321 
rect 330 321 333 324 
rect 330 324 333 327 
rect 330 327 333 330 
rect 330 330 333 333 
rect 330 333 333 336 
rect 330 336 333 339 
rect 330 339 333 342 
rect 330 342 333 345 
rect 330 345 333 348 
rect 330 348 333 351 
rect 330 351 333 354 
rect 330 354 333 357 
rect 330 357 333 360 
rect 330 360 333 363 
rect 330 363 333 366 
rect 330 366 333 369 
rect 330 369 333 372 
rect 330 372 333 375 
rect 330 375 333 378 
rect 330 378 333 381 
rect 330 381 333 384 
rect 330 384 333 387 
rect 330 387 333 390 
rect 330 390 333 393 
rect 330 393 333 396 
rect 330 396 333 399 
rect 330 399 333 402 
rect 330 402 333 405 
rect 330 405 333 408 
rect 330 408 333 411 
rect 330 411 333 414 
rect 330 414 333 417 
rect 330 417 333 420 
rect 330 420 333 423 
rect 330 423 333 426 
rect 330 426 333 429 
rect 330 429 333 432 
rect 330 432 333 435 
rect 330 435 333 438 
rect 330 438 333 441 
rect 330 441 333 444 
rect 330 444 333 447 
rect 330 447 333 450 
rect 330 450 333 453 
rect 330 453 333 456 
rect 330 456 333 459 
rect 330 459 333 462 
rect 330 462 333 465 
rect 330 465 333 468 
rect 330 468 333 471 
rect 330 471 333 474 
rect 330 474 333 477 
rect 330 477 333 480 
rect 330 480 333 483 
rect 330 483 333 486 
rect 330 486 333 489 
rect 330 489 333 492 
rect 330 492 333 495 
rect 330 495 333 498 
rect 330 498 333 501 
rect 330 501 333 504 
rect 330 504 333 507 
rect 330 507 333 510 
rect 333 0 336 3 
rect 333 3 336 6 
rect 333 6 336 9 
rect 333 9 336 12 
rect 333 12 336 15 
rect 333 15 336 18 
rect 333 18 336 21 
rect 333 21 336 24 
rect 333 24 336 27 
rect 333 27 336 30 
rect 333 30 336 33 
rect 333 33 336 36 
rect 333 36 336 39 
rect 333 39 336 42 
rect 333 42 336 45 
rect 333 45 336 48 
rect 333 48 336 51 
rect 333 51 336 54 
rect 333 54 336 57 
rect 333 57 336 60 
rect 333 60 336 63 
rect 333 63 336 66 
rect 333 66 336 69 
rect 333 69 336 72 
rect 333 72 336 75 
rect 333 75 336 78 
rect 333 78 336 81 
rect 333 81 336 84 
rect 333 84 336 87 
rect 333 87 336 90 
rect 333 90 336 93 
rect 333 93 336 96 
rect 333 96 336 99 
rect 333 99 336 102 
rect 333 102 336 105 
rect 333 105 336 108 
rect 333 108 336 111 
rect 333 111 336 114 
rect 333 114 336 117 
rect 333 117 336 120 
rect 333 120 336 123 
rect 333 123 336 126 
rect 333 126 336 129 
rect 333 129 336 132 
rect 333 132 336 135 
rect 333 135 336 138 
rect 333 138 336 141 
rect 333 141 336 144 
rect 333 144 336 147 
rect 333 147 336 150 
rect 333 150 336 153 
rect 333 153 336 156 
rect 333 156 336 159 
rect 333 159 336 162 
rect 333 162 336 165 
rect 333 165 336 168 
rect 333 168 336 171 
rect 333 171 336 174 
rect 333 174 336 177 
rect 333 177 336 180 
rect 333 180 336 183 
rect 333 183 336 186 
rect 333 186 336 189 
rect 333 189 336 192 
rect 333 192 336 195 
rect 333 195 336 198 
rect 333 198 336 201 
rect 333 201 336 204 
rect 333 204 336 207 
rect 333 207 336 210 
rect 333 210 336 213 
rect 333 213 336 216 
rect 333 216 336 219 
rect 333 219 336 222 
rect 333 222 336 225 
rect 333 225 336 228 
rect 333 228 336 231 
rect 333 231 336 234 
rect 333 234 336 237 
rect 333 237 336 240 
rect 333 240 336 243 
rect 333 243 336 246 
rect 333 246 336 249 
rect 333 249 336 252 
rect 333 252 336 255 
rect 333 255 336 258 
rect 333 258 336 261 
rect 333 261 336 264 
rect 333 264 336 267 
rect 333 267 336 270 
rect 333 270 336 273 
rect 333 273 336 276 
rect 333 276 336 279 
rect 333 279 336 282 
rect 333 282 336 285 
rect 333 285 336 288 
rect 333 288 336 291 
rect 333 291 336 294 
rect 333 294 336 297 
rect 333 297 336 300 
rect 333 300 336 303 
rect 333 303 336 306 
rect 333 306 336 309 
rect 333 309 336 312 
rect 333 312 336 315 
rect 333 315 336 318 
rect 333 318 336 321 
rect 333 324 336 327 
rect 333 327 336 330 
rect 333 330 336 333 
rect 333 333 336 336 
rect 333 336 336 339 
rect 333 339 336 342 
rect 333 342 336 345 
rect 333 345 336 348 
rect 333 348 336 351 
rect 333 351 336 354 
rect 333 354 336 357 
rect 333 357 336 360 
rect 333 360 336 363 
rect 333 363 336 366 
rect 333 366 336 369 
rect 333 372 336 375 
rect 333 375 336 378 
rect 333 381 336 384 
rect 333 384 336 387 
rect 333 387 336 390 
rect 333 390 336 393 
rect 333 393 336 396 
rect 333 396 336 399 
rect 333 399 336 402 
rect 333 402 336 405 
rect 333 405 336 408 
rect 333 408 336 411 
rect 333 411 336 414 
rect 333 414 336 417 
rect 333 417 336 420 
rect 333 420 336 423 
rect 333 423 336 426 
rect 333 426 336 429 
rect 333 429 336 432 
rect 333 432 336 435 
rect 333 435 336 438 
rect 333 438 336 441 
rect 333 441 336 444 
rect 333 444 336 447 
rect 333 447 336 450 
rect 333 450 336 453 
rect 333 453 336 456 
rect 333 456 336 459 
rect 333 459 336 462 
rect 333 462 336 465 
rect 333 465 336 468 
rect 333 468 336 471 
rect 333 471 336 474 
rect 333 474 336 477 
rect 333 477 336 480 
rect 333 480 336 483 
rect 333 483 336 486 
rect 333 486 336 489 
rect 333 489 336 492 
rect 333 492 336 495 
rect 333 495 336 498 
rect 333 498 336 501 
rect 333 501 336 504 
rect 333 504 336 507 
rect 333 507 336 510 
rect 336 0 339 3 
rect 336 3 339 6 
rect 336 6 339 9 
rect 336 9 339 12 
rect 336 12 339 15 
rect 336 15 339 18 
rect 336 18 339 21 
rect 336 21 339 24 
rect 336 24 339 27 
rect 336 27 339 30 
rect 336 30 339 33 
rect 336 33 339 36 
rect 336 36 339 39 
rect 336 39 339 42 
rect 336 42 339 45 
rect 336 45 339 48 
rect 336 48 339 51 
rect 336 51 339 54 
rect 336 54 339 57 
rect 336 57 339 60 
rect 336 60 339 63 
rect 336 63 339 66 
rect 336 66 339 69 
rect 336 69 339 72 
rect 336 72 339 75 
rect 336 75 339 78 
rect 336 78 339 81 
rect 336 81 339 84 
rect 336 84 339 87 
rect 336 87 339 90 
rect 336 90 339 93 
rect 336 93 339 96 
rect 336 96 339 99 
rect 336 99 339 102 
rect 336 102 339 105 
rect 336 105 339 108 
rect 336 108 339 111 
rect 336 111 339 114 
rect 336 114 339 117 
rect 336 117 339 120 
rect 336 120 339 123 
rect 336 123 339 126 
rect 336 126 339 129 
rect 336 129 339 132 
rect 336 132 339 135 
rect 336 135 339 138 
rect 336 138 339 141 
rect 336 141 339 144 
rect 336 144 339 147 
rect 336 147 339 150 
rect 336 150 339 153 
rect 336 153 339 156 
rect 336 156 339 159 
rect 336 159 339 162 
rect 336 162 339 165 
rect 336 165 339 168 
rect 336 168 339 171 
rect 336 171 339 174 
rect 336 174 339 177 
rect 336 177 339 180 
rect 336 180 339 183 
rect 336 183 339 186 
rect 336 186 339 189 
rect 336 189 339 192 
rect 336 192 339 195 
rect 336 195 339 198 
rect 336 198 339 201 
rect 336 201 339 204 
rect 336 204 339 207 
rect 336 207 339 210 
rect 336 210 339 213 
rect 336 213 339 216 
rect 336 216 339 219 
rect 336 219 339 222 
rect 336 222 339 225 
rect 336 225 339 228 
rect 336 228 339 231 
rect 336 231 339 234 
rect 336 234 339 237 
rect 336 237 339 240 
rect 336 240 339 243 
rect 336 243 339 246 
rect 336 246 339 249 
rect 336 249 339 252 
rect 336 252 339 255 
rect 336 255 339 258 
rect 336 258 339 261 
rect 336 261 339 264 
rect 336 264 339 267 
rect 336 267 339 270 
rect 336 270 339 273 
rect 336 273 339 276 
rect 336 276 339 279 
rect 336 279 339 282 
rect 336 282 339 285 
rect 336 285 339 288 
rect 336 288 339 291 
rect 336 291 339 294 
rect 336 294 339 297 
rect 336 297 339 300 
rect 336 300 339 303 
rect 336 303 339 306 
rect 336 306 339 309 
rect 336 309 339 312 
rect 336 312 339 315 
rect 336 315 339 318 
rect 336 318 339 321 
rect 336 321 339 324 
rect 336 324 339 327 
rect 336 327 339 330 
rect 336 330 339 333 
rect 336 333 339 336 
rect 336 336 339 339 
rect 336 339 339 342 
rect 336 342 339 345 
rect 336 345 339 348 
rect 336 348 339 351 
rect 336 351 339 354 
rect 336 354 339 357 
rect 336 357 339 360 
rect 336 360 339 363 
rect 336 363 339 366 
rect 336 366 339 369 
rect 336 369 339 372 
rect 336 372 339 375 
rect 336 375 339 378 
rect 336 378 339 381 
rect 336 381 339 384 
rect 336 384 339 387 
rect 336 387 339 390 
rect 336 390 339 393 
rect 336 393 339 396 
rect 336 396 339 399 
rect 336 399 339 402 
rect 336 402 339 405 
rect 336 405 339 408 
rect 336 408 339 411 
rect 336 411 339 414 
rect 336 414 339 417 
rect 336 417 339 420 
rect 336 420 339 423 
rect 336 423 339 426 
rect 336 426 339 429 
rect 336 429 339 432 
rect 336 432 339 435 
rect 336 435 339 438 
rect 336 438 339 441 
rect 336 441 339 444 
rect 336 444 339 447 
rect 336 447 339 450 
rect 336 450 339 453 
rect 336 453 339 456 
rect 336 456 339 459 
rect 336 459 339 462 
rect 336 462 339 465 
rect 336 465 339 468 
rect 336 468 339 471 
rect 336 471 339 474 
rect 336 474 339 477 
rect 336 477 339 480 
rect 336 480 339 483 
rect 336 483 339 486 
rect 336 486 339 489 
rect 336 489 339 492 
rect 336 492 339 495 
rect 336 495 339 498 
rect 336 498 339 501 
rect 336 501 339 504 
rect 336 504 339 507 
rect 336 507 339 510 
rect 339 0 342 3 
rect 339 3 342 6 
rect 339 6 342 9 
rect 339 9 342 12 
rect 339 12 342 15 
rect 339 15 342 18 
rect 339 18 342 21 
rect 339 21 342 24 
rect 339 24 342 27 
rect 339 27 342 30 
rect 339 30 342 33 
rect 339 33 342 36 
rect 339 36 342 39 
rect 339 39 342 42 
rect 339 42 342 45 
rect 339 45 342 48 
rect 339 48 342 51 
rect 339 51 342 54 
rect 339 54 342 57 
rect 339 57 342 60 
rect 339 60 342 63 
rect 339 63 342 66 
rect 339 66 342 69 
rect 339 69 342 72 
rect 339 72 342 75 
rect 339 75 342 78 
rect 339 78 342 81 
rect 339 81 342 84 
rect 339 84 342 87 
rect 339 87 342 90 
rect 339 90 342 93 
rect 339 93 342 96 
rect 339 96 342 99 
rect 339 99 342 102 
rect 339 102 342 105 
rect 339 105 342 108 
rect 339 108 342 111 
rect 339 111 342 114 
rect 339 114 342 117 
rect 339 117 342 120 
rect 339 120 342 123 
rect 339 123 342 126 
rect 339 126 342 129 
rect 339 129 342 132 
rect 339 132 342 135 
rect 339 135 342 138 
rect 339 138 342 141 
rect 339 141 342 144 
rect 339 144 342 147 
rect 339 147 342 150 
rect 339 150 342 153 
rect 339 153 342 156 
rect 339 156 342 159 
rect 339 159 342 162 
rect 339 162 342 165 
rect 339 165 342 168 
rect 339 168 342 171 
rect 339 171 342 174 
rect 339 174 342 177 
rect 339 177 342 180 
rect 339 180 342 183 
rect 339 183 342 186 
rect 339 186 342 189 
rect 339 189 342 192 
rect 339 192 342 195 
rect 339 195 342 198 
rect 339 198 342 201 
rect 339 201 342 204 
rect 339 204 342 207 
rect 339 207 342 210 
rect 339 210 342 213 
rect 339 213 342 216 
rect 339 216 342 219 
rect 339 219 342 222 
rect 339 222 342 225 
rect 339 225 342 228 
rect 339 228 342 231 
rect 339 231 342 234 
rect 339 234 342 237 
rect 339 237 342 240 
rect 339 240 342 243 
rect 339 243 342 246 
rect 339 246 342 249 
rect 339 249 342 252 
rect 339 252 342 255 
rect 339 255 342 258 
rect 339 258 342 261 
rect 339 261 342 264 
rect 339 264 342 267 
rect 339 267 342 270 
rect 339 270 342 273 
rect 339 273 342 276 
rect 339 276 342 279 
rect 339 279 342 282 
rect 339 282 342 285 
rect 339 285 342 288 
rect 339 288 342 291 
rect 339 291 342 294 
rect 339 294 342 297 
rect 339 297 342 300 
rect 339 300 342 303 
rect 339 303 342 306 
rect 339 306 342 309 
rect 339 309 342 312 
rect 339 312 342 315 
rect 339 315 342 318 
rect 339 318 342 321 
rect 339 321 342 324 
rect 339 324 342 327 
rect 339 327 342 330 
rect 339 330 342 333 
rect 339 333 342 336 
rect 339 336 342 339 
rect 339 339 342 342 
rect 339 342 342 345 
rect 339 345 342 348 
rect 339 348 342 351 
rect 339 351 342 354 
rect 339 354 342 357 
rect 339 357 342 360 
rect 339 360 342 363 
rect 339 363 342 366 
rect 339 366 342 369 
rect 339 369 342 372 
rect 339 372 342 375 
rect 339 375 342 378 
rect 339 378 342 381 
rect 339 381 342 384 
rect 339 384 342 387 
rect 339 387 342 390 
rect 339 390 342 393 
rect 339 393 342 396 
rect 339 396 342 399 
rect 339 399 342 402 
rect 339 402 342 405 
rect 339 405 342 408 
rect 339 408 342 411 
rect 339 411 342 414 
rect 339 414 342 417 
rect 339 417 342 420 
rect 339 420 342 423 
rect 339 423 342 426 
rect 339 426 342 429 
rect 339 429 342 432 
rect 339 432 342 435 
rect 339 435 342 438 
rect 339 438 342 441 
rect 339 441 342 444 
rect 339 444 342 447 
rect 339 447 342 450 
rect 339 450 342 453 
rect 339 453 342 456 
rect 339 456 342 459 
rect 339 459 342 462 
rect 339 462 342 465 
rect 339 465 342 468 
rect 339 468 342 471 
rect 339 471 342 474 
rect 339 474 342 477 
rect 339 477 342 480 
rect 339 480 342 483 
rect 339 483 342 486 
rect 339 486 342 489 
rect 339 489 342 492 
rect 339 492 342 495 
rect 339 495 342 498 
rect 339 498 342 501 
rect 339 501 342 504 
rect 339 504 342 507 
rect 339 507 342 510 
rect 342 0 345 3 
rect 342 3 345 6 
rect 342 6 345 9 
rect 342 9 345 12 
rect 342 12 345 15 
rect 342 15 345 18 
rect 342 18 345 21 
rect 342 21 345 24 
rect 342 24 345 27 
rect 342 27 345 30 
rect 342 30 345 33 
rect 342 33 345 36 
rect 342 36 345 39 
rect 342 39 345 42 
rect 342 42 345 45 
rect 342 45 345 48 
rect 342 48 345 51 
rect 342 51 345 54 
rect 342 54 345 57 
rect 342 57 345 60 
rect 342 60 345 63 
rect 342 63 345 66 
rect 342 66 345 69 
rect 342 69 345 72 
rect 342 72 345 75 
rect 342 75 345 78 
rect 342 78 345 81 
rect 342 81 345 84 
rect 342 84 345 87 
rect 342 87 345 90 
rect 342 90 345 93 
rect 342 93 345 96 
rect 342 96 345 99 
rect 342 99 345 102 
rect 342 102 345 105 
rect 342 105 345 108 
rect 342 108 345 111 
rect 342 111 345 114 
rect 342 114 345 117 
rect 342 117 345 120 
rect 342 120 345 123 
rect 342 123 345 126 
rect 342 126 345 129 
rect 342 129 345 132 
rect 342 132 345 135 
rect 342 135 345 138 
rect 342 138 345 141 
rect 342 141 345 144 
rect 342 144 345 147 
rect 342 147 345 150 
rect 342 150 345 153 
rect 342 153 345 156 
rect 342 156 345 159 
rect 342 159 345 162 
rect 342 162 345 165 
rect 342 165 345 168 
rect 342 168 345 171 
rect 342 171 345 174 
rect 342 174 345 177 
rect 342 177 345 180 
rect 342 180 345 183 
rect 342 183 345 186 
rect 342 186 345 189 
rect 342 189 345 192 
rect 342 192 345 195 
rect 342 195 345 198 
rect 342 198 345 201 
rect 342 201 345 204 
rect 342 204 345 207 
rect 342 207 345 210 
rect 342 210 345 213 
rect 342 213 345 216 
rect 342 216 345 219 
rect 342 219 345 222 
rect 342 222 345 225 
rect 342 225 345 228 
rect 342 228 345 231 
rect 342 231 345 234 
rect 342 234 345 237 
rect 342 237 345 240 
rect 342 240 345 243 
rect 342 243 345 246 
rect 342 246 345 249 
rect 342 249 345 252 
rect 342 252 345 255 
rect 342 255 345 258 
rect 342 258 345 261 
rect 342 261 345 264 
rect 342 264 345 267 
rect 342 267 345 270 
rect 342 270 345 273 
rect 342 273 345 276 
rect 342 276 345 279 
rect 342 279 345 282 
rect 342 282 345 285 
rect 342 285 345 288 
rect 342 288 345 291 
rect 342 291 345 294 
rect 342 294 345 297 
rect 342 297 345 300 
rect 342 300 345 303 
rect 342 303 345 306 
rect 342 306 345 309 
rect 342 309 345 312 
rect 342 312 345 315 
rect 342 315 345 318 
rect 342 318 345 321 
rect 342 321 345 324 
rect 342 324 345 327 
rect 342 327 345 330 
rect 342 330 345 333 
rect 342 333 345 336 
rect 342 336 345 339 
rect 342 339 345 342 
rect 342 342 345 345 
rect 342 345 345 348 
rect 342 348 345 351 
rect 342 351 345 354 
rect 342 354 345 357 
rect 342 357 345 360 
rect 342 360 345 363 
rect 342 363 345 366 
rect 342 366 345 369 
rect 342 369 345 372 
rect 342 372 345 375 
rect 342 375 345 378 
rect 342 378 345 381 
rect 342 381 345 384 
rect 342 384 345 387 
rect 342 387 345 390 
rect 342 390 345 393 
rect 342 393 345 396 
rect 342 396 345 399 
rect 342 399 345 402 
rect 342 402 345 405 
rect 342 405 345 408 
rect 342 408 345 411 
rect 342 411 345 414 
rect 342 414 345 417 
rect 342 417 345 420 
rect 342 420 345 423 
rect 342 423 345 426 
rect 342 426 345 429 
rect 342 429 345 432 
rect 342 432 345 435 
rect 342 435 345 438 
rect 342 438 345 441 
rect 342 441 345 444 
rect 342 444 345 447 
rect 342 447 345 450 
rect 342 450 345 453 
rect 342 453 345 456 
rect 342 456 345 459 
rect 342 459 345 462 
rect 342 462 345 465 
rect 342 465 345 468 
rect 342 468 345 471 
rect 342 471 345 474 
rect 342 474 345 477 
rect 342 477 345 480 
rect 342 480 345 483 
rect 342 483 345 486 
rect 342 486 345 489 
rect 342 489 345 492 
rect 342 492 345 495 
rect 342 495 345 498 
rect 342 498 345 501 
rect 342 501 345 504 
rect 342 504 345 507 
rect 342 507 345 510 
rect 345 0 348 3 
rect 345 3 348 6 
rect 345 6 348 9 
rect 345 9 348 12 
rect 345 12 348 15 
rect 345 15 348 18 
rect 345 18 348 21 
rect 345 21 348 24 
rect 345 24 348 27 
rect 345 27 348 30 
rect 345 30 348 33 
rect 345 33 348 36 
rect 345 36 348 39 
rect 345 39 348 42 
rect 345 42 348 45 
rect 345 45 348 48 
rect 345 48 348 51 
rect 345 51 348 54 
rect 345 54 348 57 
rect 345 57 348 60 
rect 345 60 348 63 
rect 345 63 348 66 
rect 345 66 348 69 
rect 345 69 348 72 
rect 345 72 348 75 
rect 345 75 348 78 
rect 345 78 348 81 
rect 345 81 348 84 
rect 345 84 348 87 
rect 345 87 348 90 
rect 345 90 348 93 
rect 345 93 348 96 
rect 345 96 348 99 
rect 345 99 348 102 
rect 345 102 348 105 
rect 345 105 348 108 
rect 345 108 348 111 
rect 345 111 348 114 
rect 345 114 348 117 
rect 345 117 348 120 
rect 345 120 348 123 
rect 345 123 348 126 
rect 345 126 348 129 
rect 345 129 348 132 
rect 345 132 348 135 
rect 345 135 348 138 
rect 345 138 348 141 
rect 345 141 348 144 
rect 345 144 348 147 
rect 345 147 348 150 
rect 345 150 348 153 
rect 345 153 348 156 
rect 345 156 348 159 
rect 345 159 348 162 
rect 345 162 348 165 
rect 345 165 348 168 
rect 345 168 348 171 
rect 345 171 348 174 
rect 345 174 348 177 
rect 345 177 348 180 
rect 345 180 348 183 
rect 345 183 348 186 
rect 345 186 348 189 
rect 345 189 348 192 
rect 345 192 348 195 
rect 345 195 348 198 
rect 345 198 348 201 
rect 345 201 348 204 
rect 345 204 348 207 
rect 345 207 348 210 
rect 345 210 348 213 
rect 345 213 348 216 
rect 345 216 348 219 
rect 345 219 348 222 
rect 345 222 348 225 
rect 345 225 348 228 
rect 345 228 348 231 
rect 345 231 348 234 
rect 345 234 348 237 
rect 345 237 348 240 
rect 345 240 348 243 
rect 345 243 348 246 
rect 345 246 348 249 
rect 345 249 348 252 
rect 345 252 348 255 
rect 345 255 348 258 
rect 345 258 348 261 
rect 345 261 348 264 
rect 345 264 348 267 
rect 345 267 348 270 
rect 345 270 348 273 
rect 345 273 348 276 
rect 345 276 348 279 
rect 345 279 348 282 
rect 345 282 348 285 
rect 345 285 348 288 
rect 345 288 348 291 
rect 345 291 348 294 
rect 345 294 348 297 
rect 345 297 348 300 
rect 345 300 348 303 
rect 345 303 348 306 
rect 345 306 348 309 
rect 345 309 348 312 
rect 345 312 348 315 
rect 345 315 348 318 
rect 345 318 348 321 
rect 345 321 348 324 
rect 345 324 348 327 
rect 345 327 348 330 
rect 345 330 348 333 
rect 345 333 348 336 
rect 345 336 348 339 
rect 345 339 348 342 
rect 345 342 348 345 
rect 345 345 348 348 
rect 345 348 348 351 
rect 345 351 348 354 
rect 345 354 348 357 
rect 345 357 348 360 
rect 345 360 348 363 
rect 345 363 348 366 
rect 345 366 348 369 
rect 345 369 348 372 
rect 345 372 348 375 
rect 345 375 348 378 
rect 345 378 348 381 
rect 345 381 348 384 
rect 345 384 348 387 
rect 345 387 348 390 
rect 345 390 348 393 
rect 345 393 348 396 
rect 345 396 348 399 
rect 345 399 348 402 
rect 345 402 348 405 
rect 345 405 348 408 
rect 345 408 348 411 
rect 345 411 348 414 
rect 345 414 348 417 
rect 345 417 348 420 
rect 345 420 348 423 
rect 345 423 348 426 
rect 345 426 348 429 
rect 345 429 348 432 
rect 345 432 348 435 
rect 345 435 348 438 
rect 345 438 348 441 
rect 345 441 348 444 
rect 345 444 348 447 
rect 345 447 348 450 
rect 345 450 348 453 
rect 345 453 348 456 
rect 345 456 348 459 
rect 345 459 348 462 
rect 345 462 348 465 
rect 345 465 348 468 
rect 345 468 348 471 
rect 345 471 348 474 
rect 345 474 348 477 
rect 345 477 348 480 
rect 345 480 348 483 
rect 345 483 348 486 
rect 345 486 348 489 
rect 345 489 348 492 
rect 345 492 348 495 
rect 345 495 348 498 
rect 345 498 348 501 
rect 345 501 348 504 
rect 345 504 348 507 
rect 345 507 348 510 
rect 348 0 351 3 
rect 348 3 351 6 
rect 348 6 351 9 
rect 348 9 351 12 
rect 348 12 351 15 
rect 348 15 351 18 
rect 348 18 351 21 
rect 348 21 351 24 
rect 348 24 351 27 
rect 348 27 351 30 
rect 348 30 351 33 
rect 348 33 351 36 
rect 348 36 351 39 
rect 348 39 351 42 
rect 348 42 351 45 
rect 348 45 351 48 
rect 348 48 351 51 
rect 348 51 351 54 
rect 348 54 351 57 
rect 348 57 351 60 
rect 348 60 351 63 
rect 348 63 351 66 
rect 348 66 351 69 
rect 348 69 351 72 
rect 348 72 351 75 
rect 348 75 351 78 
rect 348 78 351 81 
rect 348 81 351 84 
rect 348 84 351 87 
rect 348 87 351 90 
rect 348 90 351 93 
rect 348 93 351 96 
rect 348 96 351 99 
rect 348 99 351 102 
rect 348 102 351 105 
rect 348 105 351 108 
rect 348 108 351 111 
rect 348 111 351 114 
rect 348 114 351 117 
rect 348 117 351 120 
rect 348 120 351 123 
rect 348 123 351 126 
rect 348 126 351 129 
rect 348 129 351 132 
rect 348 132 351 135 
rect 348 135 351 138 
rect 348 138 351 141 
rect 348 141 351 144 
rect 348 144 351 147 
rect 348 147 351 150 
rect 348 150 351 153 
rect 348 153 351 156 
rect 348 156 351 159 
rect 348 159 351 162 
rect 348 162 351 165 
rect 348 165 351 168 
rect 348 168 351 171 
rect 348 171 351 174 
rect 348 174 351 177 
rect 348 177 351 180 
rect 348 180 351 183 
rect 348 183 351 186 
rect 348 186 351 189 
rect 348 189 351 192 
rect 348 192 351 195 
rect 348 195 351 198 
rect 348 198 351 201 
rect 348 201 351 204 
rect 348 204 351 207 
rect 348 207 351 210 
rect 348 210 351 213 
rect 348 213 351 216 
rect 348 216 351 219 
rect 348 219 351 222 
rect 348 222 351 225 
rect 348 225 351 228 
rect 348 228 351 231 
rect 348 231 351 234 
rect 348 234 351 237 
rect 348 237 351 240 
rect 348 240 351 243 
rect 348 243 351 246 
rect 348 246 351 249 
rect 348 249 351 252 
rect 348 252 351 255 
rect 348 255 351 258 
rect 348 258 351 261 
rect 348 261 351 264 
rect 348 264 351 267 
rect 348 267 351 270 
rect 348 270 351 273 
rect 348 273 351 276 
rect 348 276 351 279 
rect 348 279 351 282 
rect 348 282 351 285 
rect 348 285 351 288 
rect 348 288 351 291 
rect 348 291 351 294 
rect 348 294 351 297 
rect 348 297 351 300 
rect 348 300 351 303 
rect 348 303 351 306 
rect 348 306 351 309 
rect 348 309 351 312 
rect 348 312 351 315 
rect 348 315 351 318 
rect 348 318 351 321 
rect 348 321 351 324 
rect 348 324 351 327 
rect 348 327 351 330 
rect 348 330 351 333 
rect 348 333 351 336 
rect 348 336 351 339 
rect 348 339 351 342 
rect 348 342 351 345 
rect 348 345 351 348 
rect 348 348 351 351 
rect 348 351 351 354 
rect 348 354 351 357 
rect 348 357 351 360 
rect 348 360 351 363 
rect 348 363 351 366 
rect 348 366 351 369 
rect 348 369 351 372 
rect 348 372 351 375 
rect 348 375 351 378 
rect 348 378 351 381 
rect 348 381 351 384 
rect 348 384 351 387 
rect 348 387 351 390 
rect 348 390 351 393 
rect 348 393 351 396 
rect 348 396 351 399 
rect 348 399 351 402 
rect 348 402 351 405 
rect 348 405 351 408 
rect 348 408 351 411 
rect 348 411 351 414 
rect 348 414 351 417 
rect 348 417 351 420 
rect 348 420 351 423 
rect 348 423 351 426 
rect 348 426 351 429 
rect 348 429 351 432 
rect 348 432 351 435 
rect 348 435 351 438 
rect 348 438 351 441 
rect 348 441 351 444 
rect 348 444 351 447 
rect 348 447 351 450 
rect 348 450 351 453 
rect 348 453 351 456 
rect 348 456 351 459 
rect 348 459 351 462 
rect 348 462 351 465 
rect 348 465 351 468 
rect 348 468 351 471 
rect 348 471 351 474 
rect 348 474 351 477 
rect 348 477 351 480 
rect 348 480 351 483 
rect 348 483 351 486 
rect 348 486 351 489 
rect 348 489 351 492 
rect 348 492 351 495 
rect 348 495 351 498 
rect 348 498 351 501 
rect 348 501 351 504 
rect 348 504 351 507 
rect 348 507 351 510 
rect 351 0 354 3 
rect 351 3 354 6 
rect 351 6 354 9 
rect 351 9 354 12 
rect 351 12 354 15 
rect 351 15 354 18 
rect 351 18 354 21 
rect 351 21 354 24 
rect 351 24 354 27 
rect 351 27 354 30 
rect 351 30 354 33 
rect 351 33 354 36 
rect 351 36 354 39 
rect 351 39 354 42 
rect 351 42 354 45 
rect 351 45 354 48 
rect 351 48 354 51 
rect 351 51 354 54 
rect 351 54 354 57 
rect 351 57 354 60 
rect 351 60 354 63 
rect 351 63 354 66 
rect 351 66 354 69 
rect 351 69 354 72 
rect 351 72 354 75 
rect 351 75 354 78 
rect 351 78 354 81 
rect 351 81 354 84 
rect 351 84 354 87 
rect 351 87 354 90 
rect 351 90 354 93 
rect 351 93 354 96 
rect 351 96 354 99 
rect 351 99 354 102 
rect 351 102 354 105 
rect 351 105 354 108 
rect 351 108 354 111 
rect 351 111 354 114 
rect 351 114 354 117 
rect 351 117 354 120 
rect 351 120 354 123 
rect 351 123 354 126 
rect 351 126 354 129 
rect 351 129 354 132 
rect 351 132 354 135 
rect 351 135 354 138 
rect 351 138 354 141 
rect 351 141 354 144 
rect 351 144 354 147 
rect 351 147 354 150 
rect 351 150 354 153 
rect 351 153 354 156 
rect 351 156 354 159 
rect 351 159 354 162 
rect 351 162 354 165 
rect 351 165 354 168 
rect 351 168 354 171 
rect 351 171 354 174 
rect 351 174 354 177 
rect 351 177 354 180 
rect 351 180 354 183 
rect 351 183 354 186 
rect 351 186 354 189 
rect 351 189 354 192 
rect 351 192 354 195 
rect 351 195 354 198 
rect 351 198 354 201 
rect 351 201 354 204 
rect 351 204 354 207 
rect 351 207 354 210 
rect 351 210 354 213 
rect 351 213 354 216 
rect 351 216 354 219 
rect 351 219 354 222 
rect 351 222 354 225 
rect 351 225 354 228 
rect 351 228 354 231 
rect 351 231 354 234 
rect 351 234 354 237 
rect 351 237 354 240 
rect 351 240 354 243 
rect 351 243 354 246 
rect 351 246 354 249 
rect 351 249 354 252 
rect 351 252 354 255 
rect 351 255 354 258 
rect 351 258 354 261 
rect 351 261 354 264 
rect 351 264 354 267 
rect 351 267 354 270 
rect 351 270 354 273 
rect 351 273 354 276 
rect 351 276 354 279 
rect 351 279 354 282 
rect 351 282 354 285 
rect 351 285 354 288 
rect 351 288 354 291 
rect 351 291 354 294 
rect 351 294 354 297 
rect 351 297 354 300 
rect 351 300 354 303 
rect 351 303 354 306 
rect 351 306 354 309 
rect 351 309 354 312 
rect 351 312 354 315 
rect 351 315 354 318 
rect 351 318 354 321 
rect 351 321 354 324 
rect 351 324 354 327 
rect 351 327 354 330 
rect 351 330 354 333 
rect 351 333 354 336 
rect 351 336 354 339 
rect 351 339 354 342 
rect 351 342 354 345 
rect 351 345 354 348 
rect 351 348 354 351 
rect 351 351 354 354 
rect 351 354 354 357 
rect 351 357 354 360 
rect 351 360 354 363 
rect 351 363 354 366 
rect 351 366 354 369 
rect 351 369 354 372 
rect 351 372 354 375 
rect 351 375 354 378 
rect 351 378 354 381 
rect 351 381 354 384 
rect 351 384 354 387 
rect 351 387 354 390 
rect 351 390 354 393 
rect 351 393 354 396 
rect 351 396 354 399 
rect 351 399 354 402 
rect 351 402 354 405 
rect 351 405 354 408 
rect 351 408 354 411 
rect 351 411 354 414 
rect 351 414 354 417 
rect 351 417 354 420 
rect 351 420 354 423 
rect 351 423 354 426 
rect 351 426 354 429 
rect 351 429 354 432 
rect 351 432 354 435 
rect 351 435 354 438 
rect 351 438 354 441 
rect 351 441 354 444 
rect 351 444 354 447 
rect 351 447 354 450 
rect 351 450 354 453 
rect 351 453 354 456 
rect 351 456 354 459 
rect 351 459 354 462 
rect 351 462 354 465 
rect 351 465 354 468 
rect 351 468 354 471 
rect 351 471 354 474 
rect 351 474 354 477 
rect 351 477 354 480 
rect 351 480 354 483 
rect 351 483 354 486 
rect 351 486 354 489 
rect 351 489 354 492 
rect 351 492 354 495 
rect 351 495 354 498 
rect 351 498 354 501 
rect 351 501 354 504 
rect 351 504 354 507 
rect 351 507 354 510 
rect 354 0 357 3 
rect 354 3 357 6 
rect 354 6 357 9 
rect 354 9 357 12 
rect 354 12 357 15 
rect 354 15 357 18 
rect 354 18 357 21 
rect 354 21 357 24 
rect 354 24 357 27 
rect 354 27 357 30 
rect 354 30 357 33 
rect 354 33 357 36 
rect 354 36 357 39 
rect 354 39 357 42 
rect 354 42 357 45 
rect 354 45 357 48 
rect 354 48 357 51 
rect 354 51 357 54 
rect 354 54 357 57 
rect 354 57 357 60 
rect 354 60 357 63 
rect 354 63 357 66 
rect 354 66 357 69 
rect 354 69 357 72 
rect 354 72 357 75 
rect 354 75 357 78 
rect 354 78 357 81 
rect 354 81 357 84 
rect 354 84 357 87 
rect 354 87 357 90 
rect 354 90 357 93 
rect 354 93 357 96 
rect 354 96 357 99 
rect 354 99 357 102 
rect 354 102 357 105 
rect 354 105 357 108 
rect 354 108 357 111 
rect 354 111 357 114 
rect 354 114 357 117 
rect 354 117 357 120 
rect 354 120 357 123 
rect 354 123 357 126 
rect 354 126 357 129 
rect 354 129 357 132 
rect 354 132 357 135 
rect 354 135 357 138 
rect 354 138 357 141 
rect 354 141 357 144 
rect 354 144 357 147 
rect 354 147 357 150 
rect 354 150 357 153 
rect 354 153 357 156 
rect 354 156 357 159 
rect 354 159 357 162 
rect 354 162 357 165 
rect 354 165 357 168 
rect 354 168 357 171 
rect 354 171 357 174 
rect 354 174 357 177 
rect 354 177 357 180 
rect 354 180 357 183 
rect 354 183 357 186 
rect 354 186 357 189 
rect 354 189 357 192 
rect 354 192 357 195 
rect 354 195 357 198 
rect 354 198 357 201 
rect 354 201 357 204 
rect 354 204 357 207 
rect 354 207 357 210 
rect 354 210 357 213 
rect 354 213 357 216 
rect 354 216 357 219 
rect 354 219 357 222 
rect 354 222 357 225 
rect 354 225 357 228 
rect 354 228 357 231 
rect 354 231 357 234 
rect 354 234 357 237 
rect 354 237 357 240 
rect 354 240 357 243 
rect 354 243 357 246 
rect 354 246 357 249 
rect 354 249 357 252 
rect 354 252 357 255 
rect 354 255 357 258 
rect 354 258 357 261 
rect 354 261 357 264 
rect 354 264 357 267 
rect 354 267 357 270 
rect 354 270 357 273 
rect 354 273 357 276 
rect 354 276 357 279 
rect 354 279 357 282 
rect 354 282 357 285 
rect 354 285 357 288 
rect 354 288 357 291 
rect 354 291 357 294 
rect 354 294 357 297 
rect 354 297 357 300 
rect 354 300 357 303 
rect 354 303 357 306 
rect 354 306 357 309 
rect 354 309 357 312 
rect 354 312 357 315 
rect 354 315 357 318 
rect 354 318 357 321 
rect 354 321 357 324 
rect 354 324 357 327 
rect 354 327 357 330 
rect 354 330 357 333 
rect 354 333 357 336 
rect 354 336 357 339 
rect 354 339 357 342 
rect 354 342 357 345 
rect 354 345 357 348 
rect 354 348 357 351 
rect 354 351 357 354 
rect 354 354 357 357 
rect 354 357 357 360 
rect 354 360 357 363 
rect 354 363 357 366 
rect 354 366 357 369 
rect 354 369 357 372 
rect 354 372 357 375 
rect 354 375 357 378 
rect 354 378 357 381 
rect 354 381 357 384 
rect 354 384 357 387 
rect 354 387 357 390 
rect 354 390 357 393 
rect 354 393 357 396 
rect 354 396 357 399 
rect 354 399 357 402 
rect 354 402 357 405 
rect 354 405 357 408 
rect 354 408 357 411 
rect 354 411 357 414 
rect 354 414 357 417 
rect 354 417 357 420 
rect 354 420 357 423 
rect 354 423 357 426 
rect 354 426 357 429 
rect 354 429 357 432 
rect 354 432 357 435 
rect 354 435 357 438 
rect 354 438 357 441 
rect 354 441 357 444 
rect 354 444 357 447 
rect 354 447 357 450 
rect 354 450 357 453 
rect 354 453 357 456 
rect 354 456 357 459 
rect 354 459 357 462 
rect 354 462 357 465 
rect 354 465 357 468 
rect 354 468 357 471 
rect 354 471 357 474 
rect 354 474 357 477 
rect 354 477 357 480 
rect 354 480 357 483 
rect 354 483 357 486 
rect 354 486 357 489 
rect 354 489 357 492 
rect 354 492 357 495 
rect 354 495 357 498 
rect 354 498 357 501 
rect 354 501 357 504 
rect 354 504 357 507 
rect 354 507 357 510 
rect 357 0 360 3 
rect 357 3 360 6 
rect 357 6 360 9 
rect 357 9 360 12 
rect 357 12 360 15 
rect 357 15 360 18 
rect 357 18 360 21 
rect 357 21 360 24 
rect 357 24 360 27 
rect 357 27 360 30 
rect 357 30 360 33 
rect 357 33 360 36 
rect 357 36 360 39 
rect 357 39 360 42 
rect 357 42 360 45 
rect 357 45 360 48 
rect 357 48 360 51 
rect 357 51 360 54 
rect 357 54 360 57 
rect 357 57 360 60 
rect 357 60 360 63 
rect 357 63 360 66 
rect 357 66 360 69 
rect 357 69 360 72 
rect 357 72 360 75 
rect 357 75 360 78 
rect 357 78 360 81 
rect 357 81 360 84 
rect 357 84 360 87 
rect 357 87 360 90 
rect 357 90 360 93 
rect 357 93 360 96 
rect 357 96 360 99 
rect 357 99 360 102 
rect 357 102 360 105 
rect 357 105 360 108 
rect 357 108 360 111 
rect 357 111 360 114 
rect 357 114 360 117 
rect 357 117 360 120 
rect 357 120 360 123 
rect 357 123 360 126 
rect 357 126 360 129 
rect 357 129 360 132 
rect 357 132 360 135 
rect 357 135 360 138 
rect 357 138 360 141 
rect 357 141 360 144 
rect 357 144 360 147 
rect 357 147 360 150 
rect 357 150 360 153 
rect 357 153 360 156 
rect 357 156 360 159 
rect 357 159 360 162 
rect 357 162 360 165 
rect 357 165 360 168 
rect 357 168 360 171 
rect 357 171 360 174 
rect 357 174 360 177 
rect 357 177 360 180 
rect 357 180 360 183 
rect 357 183 360 186 
rect 357 186 360 189 
rect 357 189 360 192 
rect 357 192 360 195 
rect 357 195 360 198 
rect 357 198 360 201 
rect 357 201 360 204 
rect 357 204 360 207 
rect 357 207 360 210 
rect 357 210 360 213 
rect 357 213 360 216 
rect 357 216 360 219 
rect 357 219 360 222 
rect 357 222 360 225 
rect 357 225 360 228 
rect 357 228 360 231 
rect 357 231 360 234 
rect 357 234 360 237 
rect 357 237 360 240 
rect 357 240 360 243 
rect 357 243 360 246 
rect 357 246 360 249 
rect 357 249 360 252 
rect 357 252 360 255 
rect 357 255 360 258 
rect 357 258 360 261 
rect 357 261 360 264 
rect 357 264 360 267 
rect 357 267 360 270 
rect 357 270 360 273 
rect 357 273 360 276 
rect 357 276 360 279 
rect 357 279 360 282 
rect 357 282 360 285 
rect 357 285 360 288 
rect 357 288 360 291 
rect 357 291 360 294 
rect 357 294 360 297 
rect 357 297 360 300 
rect 357 300 360 303 
rect 357 303 360 306 
rect 357 306 360 309 
rect 357 309 360 312 
rect 357 312 360 315 
rect 357 315 360 318 
rect 357 318 360 321 
rect 357 321 360 324 
rect 357 324 360 327 
rect 357 327 360 330 
rect 357 330 360 333 
rect 357 333 360 336 
rect 357 336 360 339 
rect 357 339 360 342 
rect 357 342 360 345 
rect 357 345 360 348 
rect 357 348 360 351 
rect 357 351 360 354 
rect 357 354 360 357 
rect 357 357 360 360 
rect 357 360 360 363 
rect 357 363 360 366 
rect 357 366 360 369 
rect 357 369 360 372 
rect 357 372 360 375 
rect 357 375 360 378 
rect 357 378 360 381 
rect 357 381 360 384 
rect 357 384 360 387 
rect 357 387 360 390 
rect 357 390 360 393 
rect 357 393 360 396 
rect 357 396 360 399 
rect 357 399 360 402 
rect 357 402 360 405 
rect 357 405 360 408 
rect 357 408 360 411 
rect 357 411 360 414 
rect 357 414 360 417 
rect 357 417 360 420 
rect 357 420 360 423 
rect 357 423 360 426 
rect 357 426 360 429 
rect 357 429 360 432 
rect 357 432 360 435 
rect 357 435 360 438 
rect 357 438 360 441 
rect 357 441 360 444 
rect 357 444 360 447 
rect 357 447 360 450 
rect 357 450 360 453 
rect 357 453 360 456 
rect 357 456 360 459 
rect 357 459 360 462 
rect 357 462 360 465 
rect 357 465 360 468 
rect 357 468 360 471 
rect 357 471 360 474 
rect 357 474 360 477 
rect 357 477 360 480 
rect 357 480 360 483 
rect 357 483 360 486 
rect 357 486 360 489 
rect 357 489 360 492 
rect 357 492 360 495 
rect 357 495 360 498 
rect 357 498 360 501 
rect 357 501 360 504 
rect 357 504 360 507 
rect 357 507 360 510 
rect 360 0 363 3 
rect 360 3 363 6 
rect 360 6 363 9 
rect 360 9 363 12 
rect 360 12 363 15 
rect 360 15 363 18 
rect 360 18 363 21 
rect 360 21 363 24 
rect 360 24 363 27 
rect 360 27 363 30 
rect 360 30 363 33 
rect 360 33 363 36 
rect 360 36 363 39 
rect 360 39 363 42 
rect 360 42 363 45 
rect 360 45 363 48 
rect 360 48 363 51 
rect 360 51 363 54 
rect 360 54 363 57 
rect 360 57 363 60 
rect 360 60 363 63 
rect 360 63 363 66 
rect 360 66 363 69 
rect 360 69 363 72 
rect 360 72 363 75 
rect 360 75 363 78 
rect 360 78 363 81 
rect 360 81 363 84 
rect 360 84 363 87 
rect 360 87 363 90 
rect 360 90 363 93 
rect 360 93 363 96 
rect 360 96 363 99 
rect 360 99 363 102 
rect 360 102 363 105 
rect 360 105 363 108 
rect 360 108 363 111 
rect 360 111 363 114 
rect 360 114 363 117 
rect 360 117 363 120 
rect 360 120 363 123 
rect 360 123 363 126 
rect 360 126 363 129 
rect 360 129 363 132 
rect 360 132 363 135 
rect 360 135 363 138 
rect 360 138 363 141 
rect 360 141 363 144 
rect 360 144 363 147 
rect 360 147 363 150 
rect 360 150 363 153 
rect 360 153 363 156 
rect 360 156 363 159 
rect 360 159 363 162 
rect 360 162 363 165 
rect 360 165 363 168 
rect 360 168 363 171 
rect 360 171 363 174 
rect 360 174 363 177 
rect 360 177 363 180 
rect 360 180 363 183 
rect 360 183 363 186 
rect 360 186 363 189 
rect 360 189 363 192 
rect 360 192 363 195 
rect 360 195 363 198 
rect 360 198 363 201 
rect 360 201 363 204 
rect 360 204 363 207 
rect 360 207 363 210 
rect 360 210 363 213 
rect 360 213 363 216 
rect 360 216 363 219 
rect 360 219 363 222 
rect 360 222 363 225 
rect 360 225 363 228 
rect 360 228 363 231 
rect 360 231 363 234 
rect 360 234 363 237 
rect 360 237 363 240 
rect 360 240 363 243 
rect 360 243 363 246 
rect 360 246 363 249 
rect 360 249 363 252 
rect 360 252 363 255 
rect 360 255 363 258 
rect 360 258 363 261 
rect 360 261 363 264 
rect 360 264 363 267 
rect 360 267 363 270 
rect 360 270 363 273 
rect 360 273 363 276 
rect 360 276 363 279 
rect 360 279 363 282 
rect 360 282 363 285 
rect 360 285 363 288 
rect 360 288 363 291 
rect 360 291 363 294 
rect 360 294 363 297 
rect 360 297 363 300 
rect 360 300 363 303 
rect 360 303 363 306 
rect 360 306 363 309 
rect 360 309 363 312 
rect 360 312 363 315 
rect 360 315 363 318 
rect 360 318 363 321 
rect 360 321 363 324 
rect 360 324 363 327 
rect 360 327 363 330 
rect 360 330 363 333 
rect 360 333 363 336 
rect 360 336 363 339 
rect 360 339 363 342 
rect 360 342 363 345 
rect 360 345 363 348 
rect 360 348 363 351 
rect 360 351 363 354 
rect 360 354 363 357 
rect 360 357 363 360 
rect 360 360 363 363 
rect 360 363 363 366 
rect 360 366 363 369 
rect 360 369 363 372 
rect 360 372 363 375 
rect 360 375 363 378 
rect 360 378 363 381 
rect 360 381 363 384 
rect 360 384 363 387 
rect 360 387 363 390 
rect 360 390 363 393 
rect 360 393 363 396 
rect 360 396 363 399 
rect 360 399 363 402 
rect 360 402 363 405 
rect 360 405 363 408 
rect 360 408 363 411 
rect 360 411 363 414 
rect 360 414 363 417 
rect 360 417 363 420 
rect 360 420 363 423 
rect 360 423 363 426 
rect 360 426 363 429 
rect 360 429 363 432 
rect 360 432 363 435 
rect 360 435 363 438 
rect 360 438 363 441 
rect 360 441 363 444 
rect 360 444 363 447 
rect 360 447 363 450 
rect 360 450 363 453 
rect 360 453 363 456 
rect 360 456 363 459 
rect 360 459 363 462 
rect 360 462 363 465 
rect 360 465 363 468 
rect 360 468 363 471 
rect 360 471 363 474 
rect 360 474 363 477 
rect 360 477 363 480 
rect 360 480 363 483 
rect 360 483 363 486 
rect 360 486 363 489 
rect 360 489 363 492 
rect 360 492 363 495 
rect 360 495 363 498 
rect 360 498 363 501 
rect 360 501 363 504 
rect 360 504 363 507 
rect 360 507 363 510 
rect 363 0 366 3 
rect 363 3 366 6 
rect 363 6 366 9 
rect 363 9 366 12 
rect 363 12 366 15 
rect 363 15 366 18 
rect 363 18 366 21 
rect 363 21 366 24 
rect 363 24 366 27 
rect 363 27 366 30 
rect 363 30 366 33 
rect 363 33 366 36 
rect 363 36 366 39 
rect 363 39 366 42 
rect 363 42 366 45 
rect 363 45 366 48 
rect 363 48 366 51 
rect 363 51 366 54 
rect 363 54 366 57 
rect 363 57 366 60 
rect 363 60 366 63 
rect 363 63 366 66 
rect 363 66 366 69 
rect 363 69 366 72 
rect 363 72 366 75 
rect 363 75 366 78 
rect 363 78 366 81 
rect 363 81 366 84 
rect 363 84 366 87 
rect 363 87 366 90 
rect 363 90 366 93 
rect 363 93 366 96 
rect 363 96 366 99 
rect 363 99 366 102 
rect 363 102 366 105 
rect 363 105 366 108 
rect 363 108 366 111 
rect 363 111 366 114 
rect 363 114 366 117 
rect 363 117 366 120 
rect 363 120 366 123 
rect 363 123 366 126 
rect 363 126 366 129 
rect 363 129 366 132 
rect 363 132 366 135 
rect 363 135 366 138 
rect 363 138 366 141 
rect 363 141 366 144 
rect 363 144 366 147 
rect 363 147 366 150 
rect 363 150 366 153 
rect 363 153 366 156 
rect 363 156 366 159 
rect 363 159 366 162 
rect 363 162 366 165 
rect 363 165 366 168 
rect 363 168 366 171 
rect 363 171 366 174 
rect 363 174 366 177 
rect 363 177 366 180 
rect 363 180 366 183 
rect 363 183 366 186 
rect 363 186 366 189 
rect 363 189 366 192 
rect 363 192 366 195 
rect 363 195 366 198 
rect 363 198 366 201 
rect 363 201 366 204 
rect 363 204 366 207 
rect 363 207 366 210 
rect 363 210 366 213 
rect 363 213 366 216 
rect 363 216 366 219 
rect 363 219 366 222 
rect 363 222 366 225 
rect 363 225 366 228 
rect 363 228 366 231 
rect 363 231 366 234 
rect 363 234 366 237 
rect 363 237 366 240 
rect 363 240 366 243 
rect 363 243 366 246 
rect 363 246 366 249 
rect 363 249 366 252 
rect 363 252 366 255 
rect 363 255 366 258 
rect 363 258 366 261 
rect 363 261 366 264 
rect 363 264 366 267 
rect 363 267 366 270 
rect 363 270 366 273 
rect 363 273 366 276 
rect 363 276 366 279 
rect 363 279 366 282 
rect 363 282 366 285 
rect 363 285 366 288 
rect 363 288 366 291 
rect 363 291 366 294 
rect 363 294 366 297 
rect 363 297 366 300 
rect 363 300 366 303 
rect 363 303 366 306 
rect 363 306 366 309 
rect 363 309 366 312 
rect 363 312 366 315 
rect 363 315 366 318 
rect 363 318 366 321 
rect 363 321 366 324 
rect 363 324 366 327 
rect 363 327 366 330 
rect 363 330 366 333 
rect 363 333 366 336 
rect 363 336 366 339 
rect 363 339 366 342 
rect 363 342 366 345 
rect 363 345 366 348 
rect 363 348 366 351 
rect 363 351 366 354 
rect 363 354 366 357 
rect 363 357 366 360 
rect 363 360 366 363 
rect 363 363 366 366 
rect 363 366 366 369 
rect 363 369 366 372 
rect 363 372 366 375 
rect 363 375 366 378 
rect 363 378 366 381 
rect 363 381 366 384 
rect 363 384 366 387 
rect 363 387 366 390 
rect 363 390 366 393 
rect 363 393 366 396 
rect 363 396 366 399 
rect 363 399 366 402 
rect 363 402 366 405 
rect 363 405 366 408 
rect 363 408 366 411 
rect 363 411 366 414 
rect 363 414 366 417 
rect 363 417 366 420 
rect 363 420 366 423 
rect 363 423 366 426 
rect 363 426 366 429 
rect 363 429 366 432 
rect 363 432 366 435 
rect 363 435 366 438 
rect 363 438 366 441 
rect 363 441 366 444 
rect 363 444 366 447 
rect 363 447 366 450 
rect 363 450 366 453 
rect 363 453 366 456 
rect 363 456 366 459 
rect 363 459 366 462 
rect 363 462 366 465 
rect 363 465 366 468 
rect 363 468 366 471 
rect 363 471 366 474 
rect 363 474 366 477 
rect 363 477 366 480 
rect 363 480 366 483 
rect 363 483 366 486 
rect 363 486 366 489 
rect 363 489 366 492 
rect 363 492 366 495 
rect 363 495 366 498 
rect 363 498 366 501 
rect 363 501 366 504 
rect 363 504 366 507 
rect 363 507 366 510 
rect 366 0 369 3 
rect 366 3 369 6 
rect 366 6 369 9 
rect 366 9 369 12 
rect 366 12 369 15 
rect 366 15 369 18 
rect 366 18 369 21 
rect 366 21 369 24 
rect 366 24 369 27 
rect 366 27 369 30 
rect 366 30 369 33 
rect 366 33 369 36 
rect 366 36 369 39 
rect 366 39 369 42 
rect 366 42 369 45 
rect 366 45 369 48 
rect 366 48 369 51 
rect 366 51 369 54 
rect 366 54 369 57 
rect 366 57 369 60 
rect 366 60 369 63 
rect 366 63 369 66 
rect 366 66 369 69 
rect 366 69 369 72 
rect 366 72 369 75 
rect 366 75 369 78 
rect 366 78 369 81 
rect 366 81 369 84 
rect 366 84 369 87 
rect 366 87 369 90 
rect 366 93 369 96 
rect 366 96 369 99 
rect 366 99 369 102 
rect 366 102 369 105 
rect 366 105 369 108 
rect 366 108 369 111 
rect 366 111 369 114 
rect 366 114 369 117 
rect 366 117 369 120 
rect 366 120 369 123 
rect 366 123 369 126 
rect 366 126 369 129 
rect 366 129 369 132 
rect 366 132 369 135 
rect 366 135 369 138 
rect 366 138 369 141 
rect 366 141 369 144 
rect 366 144 369 147 
rect 366 147 369 150 
rect 366 150 369 153 
rect 366 153 369 156 
rect 366 156 369 159 
rect 366 159 369 162 
rect 366 162 369 165 
rect 366 165 369 168 
rect 366 168 369 171 
rect 366 171 369 174 
rect 366 174 369 177 
rect 366 180 369 183 
rect 366 183 369 186 
rect 366 189 369 192 
rect 366 192 369 195 
rect 366 195 369 198 
rect 366 198 369 201 
rect 366 201 369 204 
rect 366 204 369 207 
rect 366 207 369 210 
rect 366 210 369 213 
rect 366 213 369 216 
rect 366 216 369 219 
rect 366 219 369 222 
rect 366 222 369 225 
rect 366 225 369 228 
rect 366 228 369 231 
rect 366 231 369 234 
rect 366 237 369 240 
rect 366 240 369 243 
rect 366 243 369 246 
rect 366 246 369 249 
rect 366 249 369 252 
rect 366 252 369 255 
rect 366 255 369 258 
rect 366 258 369 261 
rect 366 261 369 264 
rect 366 264 369 267 
rect 366 267 369 270 
rect 366 270 369 273 
rect 366 273 369 276 
rect 366 276 369 279 
rect 366 279 369 282 
rect 366 282 369 285 
rect 366 285 369 288 
rect 366 288 369 291 
rect 366 291 369 294 
rect 366 294 369 297 
rect 366 297 369 300 
rect 366 300 369 303 
rect 366 303 369 306 
rect 366 306 369 309 
rect 366 309 369 312 
rect 366 312 369 315 
rect 366 315 369 318 
rect 366 318 369 321 
rect 366 321 369 324 
rect 366 324 369 327 
rect 366 327 369 330 
rect 366 330 369 333 
rect 366 333 369 336 
rect 366 336 369 339 
rect 366 339 369 342 
rect 366 342 369 345 
rect 366 345 369 348 
rect 366 348 369 351 
rect 366 351 369 354 
rect 366 354 369 357 
rect 366 357 369 360 
rect 366 360 369 363 
rect 366 363 369 366 
rect 366 366 369 369 
rect 366 372 369 375 
rect 366 375 369 378 
rect 366 378 369 381 
rect 366 381 369 384 
rect 366 384 369 387 
rect 366 387 369 390 
rect 366 390 369 393 
rect 366 393 369 396 
rect 366 396 369 399 
rect 366 399 369 402 
rect 366 402 369 405 
rect 366 405 369 408 
rect 366 408 369 411 
rect 366 411 369 414 
rect 366 414 369 417 
rect 366 417 369 420 
rect 366 420 369 423 
rect 366 423 369 426 
rect 366 426 369 429 
rect 366 429 369 432 
rect 366 432 369 435 
rect 366 435 369 438 
rect 366 438 369 441 
rect 366 441 369 444 
rect 366 444 369 447 
rect 366 447 369 450 
rect 366 450 369 453 
rect 366 453 369 456 
rect 366 456 369 459 
rect 366 459 369 462 
rect 366 462 369 465 
rect 366 468 369 471 
rect 366 471 369 474 
rect 366 474 369 477 
rect 366 477 369 480 
rect 366 480 369 483 
rect 366 483 369 486 
rect 366 486 369 489 
rect 366 489 369 492 
rect 366 492 369 495 
rect 366 495 369 498 
rect 366 498 369 501 
rect 366 501 369 504 
rect 366 504 369 507 
rect 366 507 369 510 
rect 369 0 372 3 
rect 369 3 372 6 
rect 369 6 372 9 
rect 369 9 372 12 
rect 369 12 372 15 
rect 369 15 372 18 
rect 369 18 372 21 
rect 369 21 372 24 
rect 369 24 372 27 
rect 369 27 372 30 
rect 369 30 372 33 
rect 369 33 372 36 
rect 369 36 372 39 
rect 369 39 372 42 
rect 369 42 372 45 
rect 369 45 372 48 
rect 369 48 372 51 
rect 369 51 372 54 
rect 369 54 372 57 
rect 369 57 372 60 
rect 369 60 372 63 
rect 369 63 372 66 
rect 369 66 372 69 
rect 369 69 372 72 
rect 369 72 372 75 
rect 369 75 372 78 
rect 369 78 372 81 
rect 369 81 372 84 
rect 369 84 372 87 
rect 369 87 372 90 
rect 369 90 372 93 
rect 369 93 372 96 
rect 369 96 372 99 
rect 369 99 372 102 
rect 369 102 372 105 
rect 369 105 372 108 
rect 369 108 372 111 
rect 369 111 372 114 
rect 369 114 372 117 
rect 369 117 372 120 
rect 369 120 372 123 
rect 369 123 372 126 
rect 369 126 372 129 
rect 369 129 372 132 
rect 369 132 372 135 
rect 369 135 372 138 
rect 369 138 372 141 
rect 369 141 372 144 
rect 369 144 372 147 
rect 369 147 372 150 
rect 369 150 372 153 
rect 369 153 372 156 
rect 369 156 372 159 
rect 369 159 372 162 
rect 369 162 372 165 
rect 369 165 372 168 
rect 369 168 372 171 
rect 369 171 372 174 
rect 369 174 372 177 
rect 369 177 372 180 
rect 369 180 372 183 
rect 369 183 372 186 
rect 369 186 372 189 
rect 369 189 372 192 
rect 369 192 372 195 
rect 369 195 372 198 
rect 369 198 372 201 
rect 369 201 372 204 
rect 369 204 372 207 
rect 369 207 372 210 
rect 369 210 372 213 
rect 369 213 372 216 
rect 369 216 372 219 
rect 369 219 372 222 
rect 369 222 372 225 
rect 369 225 372 228 
rect 369 228 372 231 
rect 369 231 372 234 
rect 369 234 372 237 
rect 369 237 372 240 
rect 369 240 372 243 
rect 369 243 372 246 
rect 369 246 372 249 
rect 369 249 372 252 
rect 369 252 372 255 
rect 369 255 372 258 
rect 369 258 372 261 
rect 369 261 372 264 
rect 369 264 372 267 
rect 369 267 372 270 
rect 369 270 372 273 
rect 369 273 372 276 
rect 369 276 372 279 
rect 369 279 372 282 
rect 369 282 372 285 
rect 369 285 372 288 
rect 369 288 372 291 
rect 369 291 372 294 
rect 369 294 372 297 
rect 369 297 372 300 
rect 369 300 372 303 
rect 369 303 372 306 
rect 369 306 372 309 
rect 369 309 372 312 
rect 369 312 372 315 
rect 369 315 372 318 
rect 369 318 372 321 
rect 369 321 372 324 
rect 369 324 372 327 
rect 369 327 372 330 
rect 369 330 372 333 
rect 369 333 372 336 
rect 369 336 372 339 
rect 369 339 372 342 
rect 369 342 372 345 
rect 369 345 372 348 
rect 369 348 372 351 
rect 369 351 372 354 
rect 369 354 372 357 
rect 369 357 372 360 
rect 369 360 372 363 
rect 369 363 372 366 
rect 369 366 372 369 
rect 369 369 372 372 
rect 369 372 372 375 
rect 369 375 372 378 
rect 369 378 372 381 
rect 369 381 372 384 
rect 369 384 372 387 
rect 369 387 372 390 
rect 369 390 372 393 
rect 369 393 372 396 
rect 369 396 372 399 
rect 369 399 372 402 
rect 369 402 372 405 
rect 369 405 372 408 
rect 369 408 372 411 
rect 369 411 372 414 
rect 369 414 372 417 
rect 369 417 372 420 
rect 369 420 372 423 
rect 369 423 372 426 
rect 369 426 372 429 
rect 369 429 372 432 
rect 369 432 372 435 
rect 369 435 372 438 
rect 369 438 372 441 
rect 369 441 372 444 
rect 369 444 372 447 
rect 369 447 372 450 
rect 369 450 372 453 
rect 369 453 372 456 
rect 369 456 372 459 
rect 369 459 372 462 
rect 369 462 372 465 
rect 369 465 372 468 
rect 369 468 372 471 
rect 369 471 372 474 
rect 369 474 372 477 
rect 369 477 372 480 
rect 369 480 372 483 
rect 369 483 372 486 
rect 369 486 372 489 
rect 369 489 372 492 
rect 369 492 372 495 
rect 369 495 372 498 
rect 369 498 372 501 
rect 369 501 372 504 
rect 369 504 372 507 
rect 369 507 372 510 
rect 372 0 375 3 
rect 372 3 375 6 
rect 372 6 375 9 
rect 372 9 375 12 
rect 372 12 375 15 
rect 372 15 375 18 
rect 372 18 375 21 
rect 372 21 375 24 
rect 372 24 375 27 
rect 372 27 375 30 
rect 372 30 375 33 
rect 372 33 375 36 
rect 372 36 375 39 
rect 372 39 375 42 
rect 372 42 375 45 
rect 372 45 375 48 
rect 372 48 375 51 
rect 372 51 375 54 
rect 372 54 375 57 
rect 372 57 375 60 
rect 372 60 375 63 
rect 372 63 375 66 
rect 372 66 375 69 
rect 372 69 375 72 
rect 372 72 375 75 
rect 372 75 375 78 
rect 372 78 375 81 
rect 372 81 375 84 
rect 372 84 375 87 
rect 372 87 375 90 
rect 372 90 375 93 
rect 372 93 375 96 
rect 372 96 375 99 
rect 372 99 375 102 
rect 372 102 375 105 
rect 372 105 375 108 
rect 372 108 375 111 
rect 372 111 375 114 
rect 372 114 375 117 
rect 372 117 375 120 
rect 372 120 375 123 
rect 372 123 375 126 
rect 372 126 375 129 
rect 372 129 375 132 
rect 372 132 375 135 
rect 372 135 375 138 
rect 372 138 375 141 
rect 372 141 375 144 
rect 372 144 375 147 
rect 372 147 375 150 
rect 372 150 375 153 
rect 372 153 375 156 
rect 372 156 375 159 
rect 372 159 375 162 
rect 372 162 375 165 
rect 372 165 375 168 
rect 372 168 375 171 
rect 372 171 375 174 
rect 372 174 375 177 
rect 372 177 375 180 
rect 372 180 375 183 
rect 372 183 375 186 
rect 372 186 375 189 
rect 372 189 375 192 
rect 372 192 375 195 
rect 372 195 375 198 
rect 372 198 375 201 
rect 372 201 375 204 
rect 372 204 375 207 
rect 372 207 375 210 
rect 372 210 375 213 
rect 372 213 375 216 
rect 372 216 375 219 
rect 372 219 375 222 
rect 372 222 375 225 
rect 372 225 375 228 
rect 372 228 375 231 
rect 372 231 375 234 
rect 372 234 375 237 
rect 372 237 375 240 
rect 372 240 375 243 
rect 372 243 375 246 
rect 372 246 375 249 
rect 372 249 375 252 
rect 372 252 375 255 
rect 372 255 375 258 
rect 372 258 375 261 
rect 372 261 375 264 
rect 372 264 375 267 
rect 372 267 375 270 
rect 372 270 375 273 
rect 372 273 375 276 
rect 372 276 375 279 
rect 372 279 375 282 
rect 372 282 375 285 
rect 372 285 375 288 
rect 372 288 375 291 
rect 372 291 375 294 
rect 372 294 375 297 
rect 372 297 375 300 
rect 372 300 375 303 
rect 372 303 375 306 
rect 372 306 375 309 
rect 372 309 375 312 
rect 372 312 375 315 
rect 372 315 375 318 
rect 372 318 375 321 
rect 372 321 375 324 
rect 372 324 375 327 
rect 372 327 375 330 
rect 372 330 375 333 
rect 372 333 375 336 
rect 372 336 375 339 
rect 372 339 375 342 
rect 372 342 375 345 
rect 372 345 375 348 
rect 372 348 375 351 
rect 372 351 375 354 
rect 372 354 375 357 
rect 372 357 375 360 
rect 372 360 375 363 
rect 372 363 375 366 
rect 372 366 375 369 
rect 372 369 375 372 
rect 372 372 375 375 
rect 372 375 375 378 
rect 372 378 375 381 
rect 372 381 375 384 
rect 372 384 375 387 
rect 372 387 375 390 
rect 372 390 375 393 
rect 372 393 375 396 
rect 372 396 375 399 
rect 372 399 375 402 
rect 372 402 375 405 
rect 372 405 375 408 
rect 372 408 375 411 
rect 372 411 375 414 
rect 372 414 375 417 
rect 372 417 375 420 
rect 372 420 375 423 
rect 372 423 375 426 
rect 372 426 375 429 
rect 372 429 375 432 
rect 372 432 375 435 
rect 372 435 375 438 
rect 372 438 375 441 
rect 372 441 375 444 
rect 372 444 375 447 
rect 372 447 375 450 
rect 372 450 375 453 
rect 372 453 375 456 
rect 372 456 375 459 
rect 372 459 375 462 
rect 372 462 375 465 
rect 372 465 375 468 
rect 372 468 375 471 
rect 372 471 375 474 
rect 372 474 375 477 
rect 372 477 375 480 
rect 372 480 375 483 
rect 372 483 375 486 
rect 372 486 375 489 
rect 372 489 375 492 
rect 372 492 375 495 
rect 372 495 375 498 
rect 372 498 375 501 
rect 372 501 375 504 
rect 372 504 375 507 
rect 372 507 375 510 
rect 375 0 378 3 
rect 375 3 378 6 
rect 375 6 378 9 
rect 375 9 378 12 
rect 375 12 378 15 
rect 375 15 378 18 
rect 375 18 378 21 
rect 375 21 378 24 
rect 375 24 378 27 
rect 375 27 378 30 
rect 375 30 378 33 
rect 375 33 378 36 
rect 375 36 378 39 
rect 375 39 378 42 
rect 375 42 378 45 
rect 375 45 378 48 
rect 375 48 378 51 
rect 375 51 378 54 
rect 375 54 378 57 
rect 375 57 378 60 
rect 375 60 378 63 
rect 375 63 378 66 
rect 375 66 378 69 
rect 375 69 378 72 
rect 375 72 378 75 
rect 375 75 378 78 
rect 375 78 378 81 
rect 375 81 378 84 
rect 375 84 378 87 
rect 375 87 378 90 
rect 375 90 378 93 
rect 375 93 378 96 
rect 375 96 378 99 
rect 375 99 378 102 
rect 375 102 378 105 
rect 375 105 378 108 
rect 375 108 378 111 
rect 375 111 378 114 
rect 375 114 378 117 
rect 375 117 378 120 
rect 375 120 378 123 
rect 375 123 378 126 
rect 375 126 378 129 
rect 375 129 378 132 
rect 375 132 378 135 
rect 375 135 378 138 
rect 375 138 378 141 
rect 375 141 378 144 
rect 375 144 378 147 
rect 375 147 378 150 
rect 375 150 378 153 
rect 375 153 378 156 
rect 375 156 378 159 
rect 375 159 378 162 
rect 375 162 378 165 
rect 375 165 378 168 
rect 375 168 378 171 
rect 375 171 378 174 
rect 375 174 378 177 
rect 375 177 378 180 
rect 375 180 378 183 
rect 375 183 378 186 
rect 375 186 378 189 
rect 375 189 378 192 
rect 375 192 378 195 
rect 375 195 378 198 
rect 375 198 378 201 
rect 375 201 378 204 
rect 375 204 378 207 
rect 375 207 378 210 
rect 375 210 378 213 
rect 375 213 378 216 
rect 375 216 378 219 
rect 375 219 378 222 
rect 375 222 378 225 
rect 375 225 378 228 
rect 375 228 378 231 
rect 375 231 378 234 
rect 375 234 378 237 
rect 375 237 378 240 
rect 375 240 378 243 
rect 375 243 378 246 
rect 375 246 378 249 
rect 375 249 378 252 
rect 375 252 378 255 
rect 375 255 378 258 
rect 375 258 378 261 
rect 375 261 378 264 
rect 375 264 378 267 
rect 375 267 378 270 
rect 375 270 378 273 
rect 375 273 378 276 
rect 375 276 378 279 
rect 375 279 378 282 
rect 375 282 378 285 
rect 375 285 378 288 
rect 375 288 378 291 
rect 375 291 378 294 
rect 375 294 378 297 
rect 375 297 378 300 
rect 375 300 378 303 
rect 375 303 378 306 
rect 375 306 378 309 
rect 375 309 378 312 
rect 375 312 378 315 
rect 375 315 378 318 
rect 375 318 378 321 
rect 375 321 378 324 
rect 375 324 378 327 
rect 375 327 378 330 
rect 375 330 378 333 
rect 375 333 378 336 
rect 375 336 378 339 
rect 375 339 378 342 
rect 375 342 378 345 
rect 375 345 378 348 
rect 375 348 378 351 
rect 375 351 378 354 
rect 375 354 378 357 
rect 375 357 378 360 
rect 375 360 378 363 
rect 375 363 378 366 
rect 375 366 378 369 
rect 375 369 378 372 
rect 375 372 378 375 
rect 375 375 378 378 
rect 375 378 378 381 
rect 375 381 378 384 
rect 375 384 378 387 
rect 375 387 378 390 
rect 375 390 378 393 
rect 375 393 378 396 
rect 375 396 378 399 
rect 375 399 378 402 
rect 375 402 378 405 
rect 375 405 378 408 
rect 375 408 378 411 
rect 375 411 378 414 
rect 375 414 378 417 
rect 375 417 378 420 
rect 375 420 378 423 
rect 375 423 378 426 
rect 375 426 378 429 
rect 375 429 378 432 
rect 375 432 378 435 
rect 375 435 378 438 
rect 375 438 378 441 
rect 375 441 378 444 
rect 375 444 378 447 
rect 375 447 378 450 
rect 375 450 378 453 
rect 375 453 378 456 
rect 375 456 378 459 
rect 375 459 378 462 
rect 375 462 378 465 
rect 375 465 378 468 
rect 375 468 378 471 
rect 375 471 378 474 
rect 375 474 378 477 
rect 375 477 378 480 
rect 375 480 378 483 
rect 375 483 378 486 
rect 375 486 378 489 
rect 375 489 378 492 
rect 375 492 378 495 
rect 375 495 378 498 
rect 375 498 378 501 
rect 375 501 378 504 
rect 375 504 378 507 
rect 375 507 378 510 
rect 378 0 381 3 
rect 378 3 381 6 
rect 378 6 381 9 
rect 378 9 381 12 
rect 378 12 381 15 
rect 378 15 381 18 
rect 378 18 381 21 
rect 378 21 381 24 
rect 378 24 381 27 
rect 378 27 381 30 
rect 378 30 381 33 
rect 378 33 381 36 
rect 378 36 381 39 
rect 378 39 381 42 
rect 378 42 381 45 
rect 378 45 381 48 
rect 378 48 381 51 
rect 378 51 381 54 
rect 378 54 381 57 
rect 378 57 381 60 
rect 378 60 381 63 
rect 378 63 381 66 
rect 378 66 381 69 
rect 378 69 381 72 
rect 378 72 381 75 
rect 378 75 381 78 
rect 378 78 381 81 
rect 378 81 381 84 
rect 378 84 381 87 
rect 378 87 381 90 
rect 378 90 381 93 
rect 378 93 381 96 
rect 378 96 381 99 
rect 378 99 381 102 
rect 378 102 381 105 
rect 378 105 381 108 
rect 378 108 381 111 
rect 378 111 381 114 
rect 378 114 381 117 
rect 378 117 381 120 
rect 378 120 381 123 
rect 378 123 381 126 
rect 378 126 381 129 
rect 378 129 381 132 
rect 378 132 381 135 
rect 378 135 381 138 
rect 378 138 381 141 
rect 378 141 381 144 
rect 378 144 381 147 
rect 378 147 381 150 
rect 378 150 381 153 
rect 378 153 381 156 
rect 378 156 381 159 
rect 378 159 381 162 
rect 378 162 381 165 
rect 378 165 381 168 
rect 378 168 381 171 
rect 378 171 381 174 
rect 378 174 381 177 
rect 378 177 381 180 
rect 378 180 381 183 
rect 378 183 381 186 
rect 378 186 381 189 
rect 378 189 381 192 
rect 378 192 381 195 
rect 378 195 381 198 
rect 378 198 381 201 
rect 378 201 381 204 
rect 378 204 381 207 
rect 378 207 381 210 
rect 378 210 381 213 
rect 378 213 381 216 
rect 378 216 381 219 
rect 378 219 381 222 
rect 378 222 381 225 
rect 378 225 381 228 
rect 378 228 381 231 
rect 378 231 381 234 
rect 378 234 381 237 
rect 378 237 381 240 
rect 378 240 381 243 
rect 378 243 381 246 
rect 378 246 381 249 
rect 378 249 381 252 
rect 378 252 381 255 
rect 378 255 381 258 
rect 378 258 381 261 
rect 378 261 381 264 
rect 378 264 381 267 
rect 378 267 381 270 
rect 378 270 381 273 
rect 378 273 381 276 
rect 378 276 381 279 
rect 378 279 381 282 
rect 378 282 381 285 
rect 378 285 381 288 
rect 378 288 381 291 
rect 378 291 381 294 
rect 378 294 381 297 
rect 378 297 381 300 
rect 378 300 381 303 
rect 378 303 381 306 
rect 378 306 381 309 
rect 378 309 381 312 
rect 378 312 381 315 
rect 378 315 381 318 
rect 378 318 381 321 
rect 378 321 381 324 
rect 378 324 381 327 
rect 378 327 381 330 
rect 378 330 381 333 
rect 378 333 381 336 
rect 378 336 381 339 
rect 378 339 381 342 
rect 378 342 381 345 
rect 378 345 381 348 
rect 378 348 381 351 
rect 378 351 381 354 
rect 378 354 381 357 
rect 378 357 381 360 
rect 378 360 381 363 
rect 378 363 381 366 
rect 378 366 381 369 
rect 378 369 381 372 
rect 378 372 381 375 
rect 378 375 381 378 
rect 378 378 381 381 
rect 378 381 381 384 
rect 378 384 381 387 
rect 378 387 381 390 
rect 378 390 381 393 
rect 378 393 381 396 
rect 378 396 381 399 
rect 378 399 381 402 
rect 378 402 381 405 
rect 378 405 381 408 
rect 378 408 381 411 
rect 378 411 381 414 
rect 378 414 381 417 
rect 378 417 381 420 
rect 378 420 381 423 
rect 378 423 381 426 
rect 378 426 381 429 
rect 378 429 381 432 
rect 378 432 381 435 
rect 378 435 381 438 
rect 378 438 381 441 
rect 378 441 381 444 
rect 378 444 381 447 
rect 378 447 381 450 
rect 378 450 381 453 
rect 378 453 381 456 
rect 378 456 381 459 
rect 378 459 381 462 
rect 378 462 381 465 
rect 378 465 381 468 
rect 378 468 381 471 
rect 378 471 381 474 
rect 378 474 381 477 
rect 378 477 381 480 
rect 378 480 381 483 
rect 378 483 381 486 
rect 378 486 381 489 
rect 378 489 381 492 
rect 378 492 381 495 
rect 378 495 381 498 
rect 378 498 381 501 
rect 378 501 381 504 
rect 378 504 381 507 
rect 378 507 381 510 
rect 381 0 384 3 
rect 381 3 384 6 
rect 381 6 384 9 
rect 381 9 384 12 
rect 381 12 384 15 
rect 381 15 384 18 
rect 381 18 384 21 
rect 381 21 384 24 
rect 381 24 384 27 
rect 381 27 384 30 
rect 381 30 384 33 
rect 381 33 384 36 
rect 381 36 384 39 
rect 381 39 384 42 
rect 381 42 384 45 
rect 381 45 384 48 
rect 381 48 384 51 
rect 381 51 384 54 
rect 381 54 384 57 
rect 381 57 384 60 
rect 381 60 384 63 
rect 381 63 384 66 
rect 381 66 384 69 
rect 381 69 384 72 
rect 381 72 384 75 
rect 381 75 384 78 
rect 381 78 384 81 
rect 381 81 384 84 
rect 381 84 384 87 
rect 381 87 384 90 
rect 381 90 384 93 
rect 381 93 384 96 
rect 381 96 384 99 
rect 381 99 384 102 
rect 381 102 384 105 
rect 381 105 384 108 
rect 381 108 384 111 
rect 381 111 384 114 
rect 381 114 384 117 
rect 381 117 384 120 
rect 381 120 384 123 
rect 381 123 384 126 
rect 381 126 384 129 
rect 381 132 384 135 
rect 381 135 384 138 
rect 381 138 384 141 
rect 381 141 384 144 
rect 381 144 384 147 
rect 381 147 384 150 
rect 381 150 384 153 
rect 381 153 384 156 
rect 381 156 384 159 
rect 381 159 384 162 
rect 381 162 384 165 
rect 381 165 384 168 
rect 381 168 384 171 
rect 381 171 384 174 
rect 381 174 384 177 
rect 381 177 384 180 
rect 381 180 384 183 
rect 381 183 384 186 
rect 381 189 384 192 
rect 381 192 384 195 
rect 381 195 384 198 
rect 381 198 384 201 
rect 381 201 384 204 
rect 381 204 384 207 
rect 381 207 384 210 
rect 381 210 384 213 
rect 381 213 384 216 
rect 381 216 384 219 
rect 381 219 384 222 
rect 381 222 384 225 
rect 381 228 384 231 
rect 381 231 384 234 
rect 381 234 384 237 
rect 381 237 384 240 
rect 381 240 384 243 
rect 381 243 384 246 
rect 381 246 384 249 
rect 381 249 384 252 
rect 381 252 384 255 
rect 381 255 384 258 
rect 381 258 384 261 
rect 381 261 384 264 
rect 381 264 384 267 
rect 381 267 384 270 
rect 381 270 384 273 
rect 381 276 384 279 
rect 381 279 384 282 
rect 381 285 384 288 
rect 381 288 384 291 
rect 381 291 384 294 
rect 381 294 384 297 
rect 381 297 384 300 
rect 381 300 384 303 
rect 381 303 384 306 
rect 381 306 384 309 
rect 381 309 384 312 
rect 381 312 384 315 
rect 381 315 384 318 
rect 381 318 384 321 
rect 381 321 384 324 
rect 381 324 384 327 
rect 381 327 384 330 
rect 381 330 384 333 
rect 381 333 384 336 
rect 381 336 384 339 
rect 381 339 384 342 
rect 381 342 384 345 
rect 381 345 384 348 
rect 381 348 384 351 
rect 381 351 384 354 
rect 381 354 384 357 
rect 381 357 384 360 
rect 381 360 384 363 
rect 381 363 384 366 
rect 381 366 384 369 
rect 381 369 384 372 
rect 381 372 384 375 
rect 381 375 384 378 
rect 381 381 384 384 
rect 381 384 384 387 
rect 381 387 384 390 
rect 381 390 384 393 
rect 381 393 384 396 
rect 381 396 384 399 
rect 381 399 384 402 
rect 381 402 384 405 
rect 381 405 384 408 
rect 381 408 384 411 
rect 381 411 384 414 
rect 381 414 384 417 
rect 381 417 384 420 
rect 381 420 384 423 
rect 381 423 384 426 
rect 381 426 384 429 
rect 381 429 384 432 
rect 381 432 384 435 
rect 381 435 384 438 
rect 381 438 384 441 
rect 381 441 384 444 
rect 381 444 384 447 
rect 381 447 384 450 
rect 381 450 384 453 
rect 381 453 384 456 
rect 381 456 384 459 
rect 381 459 384 462 
rect 381 462 384 465 
rect 381 465 384 468 
rect 381 468 384 471 
rect 381 471 384 474 
rect 381 474 384 477 
rect 381 477 384 480 
rect 381 480 384 483 
rect 381 483 384 486 
rect 381 486 384 489 
rect 381 489 384 492 
rect 381 492 384 495 
rect 381 495 384 498 
rect 381 498 384 501 
rect 381 501 384 504 
rect 381 504 384 507 
rect 381 507 384 510 
rect 384 0 387 3 
rect 384 3 387 6 
rect 384 6 387 9 
rect 384 9 387 12 
rect 384 12 387 15 
rect 384 15 387 18 
rect 384 18 387 21 
rect 384 21 387 24 
rect 384 24 387 27 
rect 384 27 387 30 
rect 384 30 387 33 
rect 384 33 387 36 
rect 384 36 387 39 
rect 384 39 387 42 
rect 384 42 387 45 
rect 384 45 387 48 
rect 384 48 387 51 
rect 384 51 387 54 
rect 384 54 387 57 
rect 384 57 387 60 
rect 384 60 387 63 
rect 384 63 387 66 
rect 384 66 387 69 
rect 384 69 387 72 
rect 384 72 387 75 
rect 384 75 387 78 
rect 384 78 387 81 
rect 384 81 387 84 
rect 384 84 387 87 
rect 384 87 387 90 
rect 384 90 387 93 
rect 384 93 387 96 
rect 384 96 387 99 
rect 384 99 387 102 
rect 384 102 387 105 
rect 384 105 387 108 
rect 384 108 387 111 
rect 384 111 387 114 
rect 384 114 387 117 
rect 384 117 387 120 
rect 384 120 387 123 
rect 384 123 387 126 
rect 384 126 387 129 
rect 384 129 387 132 
rect 384 132 387 135 
rect 384 135 387 138 
rect 384 138 387 141 
rect 384 141 387 144 
rect 384 144 387 147 
rect 384 147 387 150 
rect 384 150 387 153 
rect 384 153 387 156 
rect 384 156 387 159 
rect 384 159 387 162 
rect 384 162 387 165 
rect 384 165 387 168 
rect 384 168 387 171 
rect 384 171 387 174 
rect 384 174 387 177 
rect 384 177 387 180 
rect 384 180 387 183 
rect 384 183 387 186 
rect 384 186 387 189 
rect 384 189 387 192 
rect 384 192 387 195 
rect 384 195 387 198 
rect 384 198 387 201 
rect 384 201 387 204 
rect 384 204 387 207 
rect 384 207 387 210 
rect 384 210 387 213 
rect 384 213 387 216 
rect 384 216 387 219 
rect 384 219 387 222 
rect 384 222 387 225 
rect 384 225 387 228 
rect 384 228 387 231 
rect 384 231 387 234 
rect 384 234 387 237 
rect 384 237 387 240 
rect 384 240 387 243 
rect 384 243 387 246 
rect 384 246 387 249 
rect 384 249 387 252 
rect 384 252 387 255 
rect 384 255 387 258 
rect 384 258 387 261 
rect 384 261 387 264 
rect 384 264 387 267 
rect 384 267 387 270 
rect 384 270 387 273 
rect 384 273 387 276 
rect 384 276 387 279 
rect 384 279 387 282 
rect 384 282 387 285 
rect 384 285 387 288 
rect 384 288 387 291 
rect 384 291 387 294 
rect 384 294 387 297 
rect 384 297 387 300 
rect 384 300 387 303 
rect 384 303 387 306 
rect 384 306 387 309 
rect 384 309 387 312 
rect 384 312 387 315 
rect 384 315 387 318 
rect 384 318 387 321 
rect 384 321 387 324 
rect 384 324 387 327 
rect 384 327 387 330 
rect 384 330 387 333 
rect 384 333 387 336 
rect 384 336 387 339 
rect 384 339 387 342 
rect 384 342 387 345 
rect 384 345 387 348 
rect 384 348 387 351 
rect 384 351 387 354 
rect 384 354 387 357 
rect 384 357 387 360 
rect 384 360 387 363 
rect 384 363 387 366 
rect 384 366 387 369 
rect 384 369 387 372 
rect 384 372 387 375 
rect 384 375 387 378 
rect 384 378 387 381 
rect 384 381 387 384 
rect 384 384 387 387 
rect 384 387 387 390 
rect 384 390 387 393 
rect 384 393 387 396 
rect 384 396 387 399 
rect 384 399 387 402 
rect 384 402 387 405 
rect 384 405 387 408 
rect 384 408 387 411 
rect 384 411 387 414 
rect 384 414 387 417 
rect 384 417 387 420 
rect 384 420 387 423 
rect 384 423 387 426 
rect 384 426 387 429 
rect 384 429 387 432 
rect 384 432 387 435 
rect 384 435 387 438 
rect 384 438 387 441 
rect 384 441 387 444 
rect 384 444 387 447 
rect 384 447 387 450 
rect 384 450 387 453 
rect 384 453 387 456 
rect 384 456 387 459 
rect 384 459 387 462 
rect 384 462 387 465 
rect 384 465 387 468 
rect 384 468 387 471 
rect 384 471 387 474 
rect 384 474 387 477 
rect 384 477 387 480 
rect 384 480 387 483 
rect 384 483 387 486 
rect 384 486 387 489 
rect 384 489 387 492 
rect 384 492 387 495 
rect 384 495 387 498 
rect 384 498 387 501 
rect 384 501 387 504 
rect 384 504 387 507 
rect 384 507 387 510 
rect 387 0 390 3 
rect 387 3 390 6 
rect 387 6 390 9 
rect 387 9 390 12 
rect 387 12 390 15 
rect 387 15 390 18 
rect 387 18 390 21 
rect 387 21 390 24 
rect 387 24 390 27 
rect 387 27 390 30 
rect 387 30 390 33 
rect 387 33 390 36 
rect 387 36 390 39 
rect 387 39 390 42 
rect 387 42 390 45 
rect 387 45 390 48 
rect 387 48 390 51 
rect 387 51 390 54 
rect 387 54 390 57 
rect 387 57 390 60 
rect 387 60 390 63 
rect 387 63 390 66 
rect 387 66 390 69 
rect 387 69 390 72 
rect 387 72 390 75 
rect 387 75 390 78 
rect 387 78 390 81 
rect 387 81 390 84 
rect 387 84 390 87 
rect 387 87 390 90 
rect 387 90 390 93 
rect 387 93 390 96 
rect 387 96 390 99 
rect 387 99 390 102 
rect 387 102 390 105 
rect 387 105 390 108 
rect 387 108 390 111 
rect 387 111 390 114 
rect 387 114 390 117 
rect 387 117 390 120 
rect 387 120 390 123 
rect 387 123 390 126 
rect 387 126 390 129 
rect 387 129 390 132 
rect 387 132 390 135 
rect 387 135 390 138 
rect 387 138 390 141 
rect 387 141 390 144 
rect 387 144 390 147 
rect 387 147 390 150 
rect 387 150 390 153 
rect 387 153 390 156 
rect 387 156 390 159 
rect 387 159 390 162 
rect 387 162 390 165 
rect 387 165 390 168 
rect 387 168 390 171 
rect 387 171 390 174 
rect 387 174 390 177 
rect 387 177 390 180 
rect 387 180 390 183 
rect 387 183 390 186 
rect 387 186 390 189 
rect 387 189 390 192 
rect 387 192 390 195 
rect 387 195 390 198 
rect 387 198 390 201 
rect 387 201 390 204 
rect 387 204 390 207 
rect 387 207 390 210 
rect 387 210 390 213 
rect 387 213 390 216 
rect 387 216 390 219 
rect 387 219 390 222 
rect 387 222 390 225 
rect 387 225 390 228 
rect 387 228 390 231 
rect 387 231 390 234 
rect 387 234 390 237 
rect 387 237 390 240 
rect 387 240 390 243 
rect 387 243 390 246 
rect 387 246 390 249 
rect 387 249 390 252 
rect 387 252 390 255 
rect 387 255 390 258 
rect 387 258 390 261 
rect 387 261 390 264 
rect 387 264 390 267 
rect 387 267 390 270 
rect 387 270 390 273 
rect 387 273 390 276 
rect 387 276 390 279 
rect 387 279 390 282 
rect 387 282 390 285 
rect 387 285 390 288 
rect 387 288 390 291 
rect 387 291 390 294 
rect 387 294 390 297 
rect 387 297 390 300 
rect 387 300 390 303 
rect 387 303 390 306 
rect 387 306 390 309 
rect 387 309 390 312 
rect 387 312 390 315 
rect 387 315 390 318 
rect 387 318 390 321 
rect 387 321 390 324 
rect 387 324 390 327 
rect 387 327 390 330 
rect 387 330 390 333 
rect 387 333 390 336 
rect 387 336 390 339 
rect 387 339 390 342 
rect 387 342 390 345 
rect 387 345 390 348 
rect 387 348 390 351 
rect 387 351 390 354 
rect 387 354 390 357 
rect 387 357 390 360 
rect 387 360 390 363 
rect 387 363 390 366 
rect 387 366 390 369 
rect 387 369 390 372 
rect 387 372 390 375 
rect 387 375 390 378 
rect 387 378 390 381 
rect 387 381 390 384 
rect 387 384 390 387 
rect 387 387 390 390 
rect 387 390 390 393 
rect 387 393 390 396 
rect 387 396 390 399 
rect 387 399 390 402 
rect 387 402 390 405 
rect 387 405 390 408 
rect 387 408 390 411 
rect 387 411 390 414 
rect 387 414 390 417 
rect 387 417 390 420 
rect 387 420 390 423 
rect 387 423 390 426 
rect 387 426 390 429 
rect 387 429 390 432 
rect 387 432 390 435 
rect 387 435 390 438 
rect 387 438 390 441 
rect 387 441 390 444 
rect 387 444 390 447 
rect 387 447 390 450 
rect 387 450 390 453 
rect 387 453 390 456 
rect 387 456 390 459 
rect 387 459 390 462 
rect 387 462 390 465 
rect 387 465 390 468 
rect 387 468 390 471 
rect 387 471 390 474 
rect 387 474 390 477 
rect 387 477 390 480 
rect 387 480 390 483 
rect 387 483 390 486 
rect 387 486 390 489 
rect 387 489 390 492 
rect 387 492 390 495 
rect 387 495 390 498 
rect 387 498 390 501 
rect 387 501 390 504 
rect 387 504 390 507 
rect 387 507 390 510 
rect 390 0 393 3 
rect 390 3 393 6 
rect 390 6 393 9 
rect 390 9 393 12 
rect 390 12 393 15 
rect 390 15 393 18 
rect 390 18 393 21 
rect 390 21 393 24 
rect 390 24 393 27 
rect 390 27 393 30 
rect 390 30 393 33 
rect 390 33 393 36 
rect 390 36 393 39 
rect 390 39 393 42 
rect 390 42 393 45 
rect 390 45 393 48 
rect 390 48 393 51 
rect 390 51 393 54 
rect 390 54 393 57 
rect 390 57 393 60 
rect 390 60 393 63 
rect 390 63 393 66 
rect 390 66 393 69 
rect 390 69 393 72 
rect 390 72 393 75 
rect 390 75 393 78 
rect 390 78 393 81 
rect 390 81 393 84 
rect 390 84 393 87 
rect 390 87 393 90 
rect 390 90 393 93 
rect 390 93 393 96 
rect 390 96 393 99 
rect 390 99 393 102 
rect 390 102 393 105 
rect 390 105 393 108 
rect 390 108 393 111 
rect 390 111 393 114 
rect 390 114 393 117 
rect 390 117 393 120 
rect 390 120 393 123 
rect 390 123 393 126 
rect 390 126 393 129 
rect 390 129 393 132 
rect 390 132 393 135 
rect 390 135 393 138 
rect 390 138 393 141 
rect 390 141 393 144 
rect 390 144 393 147 
rect 390 147 393 150 
rect 390 150 393 153 
rect 390 153 393 156 
rect 390 156 393 159 
rect 390 159 393 162 
rect 390 162 393 165 
rect 390 165 393 168 
rect 390 168 393 171 
rect 390 171 393 174 
rect 390 174 393 177 
rect 390 177 393 180 
rect 390 180 393 183 
rect 390 183 393 186 
rect 390 186 393 189 
rect 390 189 393 192 
rect 390 192 393 195 
rect 390 195 393 198 
rect 390 198 393 201 
rect 390 201 393 204 
rect 390 204 393 207 
rect 390 207 393 210 
rect 390 210 393 213 
rect 390 213 393 216 
rect 390 216 393 219 
rect 390 219 393 222 
rect 390 222 393 225 
rect 390 225 393 228 
rect 390 228 393 231 
rect 390 231 393 234 
rect 390 234 393 237 
rect 390 237 393 240 
rect 390 240 393 243 
rect 390 243 393 246 
rect 390 246 393 249 
rect 390 249 393 252 
rect 390 252 393 255 
rect 390 255 393 258 
rect 390 258 393 261 
rect 390 261 393 264 
rect 390 264 393 267 
rect 390 267 393 270 
rect 390 270 393 273 
rect 390 273 393 276 
rect 390 276 393 279 
rect 390 279 393 282 
rect 390 282 393 285 
rect 390 285 393 288 
rect 390 288 393 291 
rect 390 291 393 294 
rect 390 294 393 297 
rect 390 297 393 300 
rect 390 300 393 303 
rect 390 303 393 306 
rect 390 306 393 309 
rect 390 309 393 312 
rect 390 312 393 315 
rect 390 315 393 318 
rect 390 318 393 321 
rect 390 321 393 324 
rect 390 324 393 327 
rect 390 327 393 330 
rect 390 330 393 333 
rect 390 333 393 336 
rect 390 336 393 339 
rect 390 339 393 342 
rect 390 342 393 345 
rect 390 345 393 348 
rect 390 348 393 351 
rect 390 351 393 354 
rect 390 354 393 357 
rect 390 357 393 360 
rect 390 360 393 363 
rect 390 363 393 366 
rect 390 366 393 369 
rect 390 369 393 372 
rect 390 372 393 375 
rect 390 375 393 378 
rect 390 378 393 381 
rect 390 381 393 384 
rect 390 384 393 387 
rect 390 387 393 390 
rect 390 390 393 393 
rect 390 393 393 396 
rect 390 396 393 399 
rect 390 399 393 402 
rect 390 402 393 405 
rect 390 405 393 408 
rect 390 408 393 411 
rect 390 411 393 414 
rect 390 414 393 417 
rect 390 417 393 420 
rect 390 420 393 423 
rect 390 423 393 426 
rect 390 426 393 429 
rect 390 429 393 432 
rect 390 432 393 435 
rect 390 435 393 438 
rect 390 438 393 441 
rect 390 441 393 444 
rect 390 444 393 447 
rect 390 447 393 450 
rect 390 450 393 453 
rect 390 453 393 456 
rect 390 456 393 459 
rect 390 459 393 462 
rect 390 462 393 465 
rect 390 465 393 468 
rect 390 468 393 471 
rect 390 471 393 474 
rect 390 474 393 477 
rect 390 477 393 480 
rect 390 480 393 483 
rect 390 483 393 486 
rect 390 486 393 489 
rect 390 489 393 492 
rect 390 492 393 495 
rect 390 495 393 498 
rect 390 498 393 501 
rect 390 501 393 504 
rect 390 504 393 507 
rect 390 507 393 510 
rect 393 0 396 3 
rect 393 3 396 6 
rect 393 6 396 9 
rect 393 9 396 12 
rect 393 12 396 15 
rect 393 15 396 18 
rect 393 18 396 21 
rect 393 21 396 24 
rect 393 24 396 27 
rect 393 27 396 30 
rect 393 30 396 33 
rect 393 33 396 36 
rect 393 36 396 39 
rect 393 39 396 42 
rect 393 42 396 45 
rect 393 45 396 48 
rect 393 48 396 51 
rect 393 51 396 54 
rect 393 54 396 57 
rect 393 57 396 60 
rect 393 60 396 63 
rect 393 63 396 66 
rect 393 66 396 69 
rect 393 69 396 72 
rect 393 72 396 75 
rect 393 75 396 78 
rect 393 78 396 81 
rect 393 81 396 84 
rect 393 84 396 87 
rect 393 87 396 90 
rect 393 90 396 93 
rect 393 93 396 96 
rect 393 96 396 99 
rect 393 99 396 102 
rect 393 102 396 105 
rect 393 105 396 108 
rect 393 108 396 111 
rect 393 111 396 114 
rect 393 114 396 117 
rect 393 117 396 120 
rect 393 120 396 123 
rect 393 123 396 126 
rect 393 126 396 129 
rect 393 129 396 132 
rect 393 132 396 135 
rect 393 135 396 138 
rect 393 138 396 141 
rect 393 141 396 144 
rect 393 144 396 147 
rect 393 147 396 150 
rect 393 150 396 153 
rect 393 153 396 156 
rect 393 156 396 159 
rect 393 159 396 162 
rect 393 162 396 165 
rect 393 165 396 168 
rect 393 168 396 171 
rect 393 171 396 174 
rect 393 174 396 177 
rect 393 177 396 180 
rect 393 180 396 183 
rect 393 183 396 186 
rect 393 186 396 189 
rect 393 189 396 192 
rect 393 192 396 195 
rect 393 195 396 198 
rect 393 198 396 201 
rect 393 201 396 204 
rect 393 204 396 207 
rect 393 207 396 210 
rect 393 210 396 213 
rect 393 213 396 216 
rect 393 216 396 219 
rect 393 219 396 222 
rect 393 222 396 225 
rect 393 225 396 228 
rect 393 228 396 231 
rect 393 231 396 234 
rect 393 234 396 237 
rect 393 237 396 240 
rect 393 240 396 243 
rect 393 243 396 246 
rect 393 246 396 249 
rect 393 249 396 252 
rect 393 252 396 255 
rect 393 255 396 258 
rect 393 258 396 261 
rect 393 261 396 264 
rect 393 264 396 267 
rect 393 267 396 270 
rect 393 270 396 273 
rect 393 273 396 276 
rect 393 276 396 279 
rect 393 279 396 282 
rect 393 282 396 285 
rect 393 285 396 288 
rect 393 288 396 291 
rect 393 291 396 294 
rect 393 294 396 297 
rect 393 297 396 300 
rect 393 300 396 303 
rect 393 303 396 306 
rect 393 306 396 309 
rect 393 309 396 312 
rect 393 312 396 315 
rect 393 315 396 318 
rect 393 318 396 321 
rect 393 321 396 324 
rect 393 324 396 327 
rect 393 327 396 330 
rect 393 330 396 333 
rect 393 333 396 336 
rect 393 336 396 339 
rect 393 339 396 342 
rect 393 342 396 345 
rect 393 345 396 348 
rect 393 348 396 351 
rect 393 351 396 354 
rect 393 354 396 357 
rect 393 357 396 360 
rect 393 360 396 363 
rect 393 363 396 366 
rect 393 366 396 369 
rect 393 369 396 372 
rect 393 372 396 375 
rect 393 375 396 378 
rect 393 378 396 381 
rect 393 381 396 384 
rect 393 384 396 387 
rect 393 387 396 390 
rect 393 390 396 393 
rect 393 393 396 396 
rect 393 396 396 399 
rect 393 399 396 402 
rect 393 402 396 405 
rect 393 405 396 408 
rect 393 408 396 411 
rect 393 411 396 414 
rect 393 414 396 417 
rect 393 417 396 420 
rect 393 420 396 423 
rect 393 423 396 426 
rect 393 426 396 429 
rect 393 429 396 432 
rect 393 432 396 435 
rect 393 435 396 438 
rect 393 438 396 441 
rect 393 441 396 444 
rect 393 444 396 447 
rect 393 447 396 450 
rect 393 450 396 453 
rect 393 453 396 456 
rect 393 456 396 459 
rect 393 459 396 462 
rect 393 462 396 465 
rect 393 465 396 468 
rect 393 468 396 471 
rect 393 471 396 474 
rect 393 474 396 477 
rect 393 477 396 480 
rect 393 480 396 483 
rect 393 483 396 486 
rect 393 486 396 489 
rect 393 489 396 492 
rect 393 492 396 495 
rect 393 495 396 498 
rect 393 498 396 501 
rect 393 501 396 504 
rect 393 504 396 507 
rect 393 507 396 510 
rect 396 0 399 3 
rect 396 3 399 6 
rect 396 6 399 9 
rect 396 9 399 12 
rect 396 12 399 15 
rect 396 15 399 18 
rect 396 18 399 21 
rect 396 21 399 24 
rect 396 24 399 27 
rect 396 27 399 30 
rect 396 30 399 33 
rect 396 33 399 36 
rect 396 36 399 39 
rect 396 39 399 42 
rect 396 42 399 45 
rect 396 45 399 48 
rect 396 48 399 51 
rect 396 51 399 54 
rect 396 54 399 57 
rect 396 57 399 60 
rect 396 60 399 63 
rect 396 63 399 66 
rect 396 66 399 69 
rect 396 69 399 72 
rect 396 72 399 75 
rect 396 75 399 78 
rect 396 78 399 81 
rect 396 81 399 84 
rect 396 84 399 87 
rect 396 87 399 90 
rect 396 90 399 93 
rect 396 93 399 96 
rect 396 96 399 99 
rect 396 99 399 102 
rect 396 102 399 105 
rect 396 105 399 108 
rect 396 108 399 111 
rect 396 111 399 114 
rect 396 114 399 117 
rect 396 117 399 120 
rect 396 120 399 123 
rect 396 123 399 126 
rect 396 126 399 129 
rect 396 129 399 132 
rect 396 132 399 135 
rect 396 135 399 138 
rect 396 138 399 141 
rect 396 141 399 144 
rect 396 144 399 147 
rect 396 147 399 150 
rect 396 150 399 153 
rect 396 153 399 156 
rect 396 156 399 159 
rect 396 159 399 162 
rect 396 162 399 165 
rect 396 165 399 168 
rect 396 168 399 171 
rect 396 171 399 174 
rect 396 174 399 177 
rect 396 177 399 180 
rect 396 180 399 183 
rect 396 183 399 186 
rect 396 186 399 189 
rect 396 189 399 192 
rect 396 192 399 195 
rect 396 195 399 198 
rect 396 198 399 201 
rect 396 201 399 204 
rect 396 204 399 207 
rect 396 207 399 210 
rect 396 210 399 213 
rect 396 213 399 216 
rect 396 216 399 219 
rect 396 219 399 222 
rect 396 222 399 225 
rect 396 225 399 228 
rect 396 228 399 231 
rect 396 231 399 234 
rect 396 234 399 237 
rect 396 237 399 240 
rect 396 240 399 243 
rect 396 243 399 246 
rect 396 246 399 249 
rect 396 249 399 252 
rect 396 252 399 255 
rect 396 255 399 258 
rect 396 258 399 261 
rect 396 261 399 264 
rect 396 264 399 267 
rect 396 267 399 270 
rect 396 270 399 273 
rect 396 273 399 276 
rect 396 276 399 279 
rect 396 279 399 282 
rect 396 282 399 285 
rect 396 285 399 288 
rect 396 288 399 291 
rect 396 291 399 294 
rect 396 294 399 297 
rect 396 297 399 300 
rect 396 300 399 303 
rect 396 303 399 306 
rect 396 306 399 309 
rect 396 309 399 312 
rect 396 312 399 315 
rect 396 315 399 318 
rect 396 318 399 321 
rect 396 321 399 324 
rect 396 324 399 327 
rect 396 327 399 330 
rect 396 330 399 333 
rect 396 333 399 336 
rect 396 336 399 339 
rect 396 339 399 342 
rect 396 342 399 345 
rect 396 345 399 348 
rect 396 348 399 351 
rect 396 351 399 354 
rect 396 354 399 357 
rect 396 357 399 360 
rect 396 360 399 363 
rect 396 363 399 366 
rect 396 366 399 369 
rect 396 369 399 372 
rect 396 372 399 375 
rect 396 375 399 378 
rect 396 378 399 381 
rect 396 381 399 384 
rect 396 384 399 387 
rect 396 387 399 390 
rect 396 390 399 393 
rect 396 393 399 396 
rect 396 396 399 399 
rect 396 399 399 402 
rect 396 402 399 405 
rect 396 405 399 408 
rect 396 408 399 411 
rect 396 411 399 414 
rect 396 414 399 417 
rect 396 417 399 420 
rect 396 420 399 423 
rect 396 423 399 426 
rect 396 426 399 429 
rect 396 429 399 432 
rect 396 432 399 435 
rect 396 435 399 438 
rect 396 438 399 441 
rect 396 441 399 444 
rect 396 444 399 447 
rect 396 447 399 450 
rect 396 450 399 453 
rect 396 453 399 456 
rect 396 456 399 459 
rect 396 459 399 462 
rect 396 462 399 465 
rect 396 465 399 468 
rect 396 468 399 471 
rect 396 471 399 474 
rect 396 474 399 477 
rect 396 477 399 480 
rect 396 480 399 483 
rect 396 483 399 486 
rect 396 486 399 489 
rect 396 489 399 492 
rect 396 492 399 495 
rect 396 495 399 498 
rect 396 498 399 501 
rect 396 501 399 504 
rect 396 504 399 507 
rect 396 507 399 510 
rect 399 0 402 3 
rect 399 3 402 6 
rect 399 6 402 9 
rect 399 9 402 12 
rect 399 12 402 15 
rect 399 15 402 18 
rect 399 18 402 21 
rect 399 21 402 24 
rect 399 24 402 27 
rect 399 27 402 30 
rect 399 30 402 33 
rect 399 33 402 36 
rect 399 36 402 39 
rect 399 39 402 42 
rect 399 42 402 45 
rect 399 45 402 48 
rect 399 48 402 51 
rect 399 51 402 54 
rect 399 54 402 57 
rect 399 57 402 60 
rect 399 60 402 63 
rect 399 63 402 66 
rect 399 66 402 69 
rect 399 69 402 72 
rect 399 72 402 75 
rect 399 75 402 78 
rect 399 78 402 81 
rect 399 81 402 84 
rect 399 84 402 87 
rect 399 87 402 90 
rect 399 90 402 93 
rect 399 93 402 96 
rect 399 96 402 99 
rect 399 99 402 102 
rect 399 102 402 105 
rect 399 105 402 108 
rect 399 108 402 111 
rect 399 111 402 114 
rect 399 114 402 117 
rect 399 117 402 120 
rect 399 120 402 123 
rect 399 123 402 126 
rect 399 126 402 129 
rect 399 129 402 132 
rect 399 132 402 135 
rect 399 135 402 138 
rect 399 138 402 141 
rect 399 141 402 144 
rect 399 144 402 147 
rect 399 147 402 150 
rect 399 150 402 153 
rect 399 153 402 156 
rect 399 156 402 159 
rect 399 159 402 162 
rect 399 162 402 165 
rect 399 165 402 168 
rect 399 168 402 171 
rect 399 171 402 174 
rect 399 174 402 177 
rect 399 177 402 180 
rect 399 180 402 183 
rect 399 183 402 186 
rect 399 186 402 189 
rect 399 189 402 192 
rect 399 192 402 195 
rect 399 195 402 198 
rect 399 198 402 201 
rect 399 201 402 204 
rect 399 204 402 207 
rect 399 207 402 210 
rect 399 210 402 213 
rect 399 213 402 216 
rect 399 216 402 219 
rect 399 219 402 222 
rect 399 222 402 225 
rect 399 225 402 228 
rect 399 228 402 231 
rect 399 231 402 234 
rect 399 234 402 237 
rect 399 237 402 240 
rect 399 240 402 243 
rect 399 243 402 246 
rect 399 246 402 249 
rect 399 249 402 252 
rect 399 252 402 255 
rect 399 255 402 258 
rect 399 258 402 261 
rect 399 261 402 264 
rect 399 264 402 267 
rect 399 267 402 270 
rect 399 270 402 273 
rect 399 273 402 276 
rect 399 276 402 279 
rect 399 279 402 282 
rect 399 282 402 285 
rect 399 285 402 288 
rect 399 288 402 291 
rect 399 291 402 294 
rect 399 294 402 297 
rect 399 297 402 300 
rect 399 300 402 303 
rect 399 303 402 306 
rect 399 306 402 309 
rect 399 309 402 312 
rect 399 312 402 315 
rect 399 315 402 318 
rect 399 318 402 321 
rect 399 321 402 324 
rect 399 324 402 327 
rect 399 327 402 330 
rect 399 330 402 333 
rect 399 333 402 336 
rect 399 336 402 339 
rect 399 339 402 342 
rect 399 342 402 345 
rect 399 345 402 348 
rect 399 348 402 351 
rect 399 351 402 354 
rect 399 354 402 357 
rect 399 357 402 360 
rect 399 360 402 363 
rect 399 363 402 366 
rect 399 366 402 369 
rect 399 369 402 372 
rect 399 372 402 375 
rect 399 375 402 378 
rect 399 378 402 381 
rect 399 381 402 384 
rect 399 384 402 387 
rect 399 387 402 390 
rect 399 390 402 393 
rect 399 393 402 396 
rect 399 396 402 399 
rect 399 399 402 402 
rect 399 402 402 405 
rect 399 405 402 408 
rect 399 408 402 411 
rect 399 411 402 414 
rect 399 414 402 417 
rect 399 417 402 420 
rect 399 420 402 423 
rect 399 423 402 426 
rect 399 426 402 429 
rect 399 429 402 432 
rect 399 432 402 435 
rect 399 435 402 438 
rect 399 438 402 441 
rect 399 441 402 444 
rect 399 444 402 447 
rect 399 447 402 450 
rect 399 450 402 453 
rect 399 453 402 456 
rect 399 456 402 459 
rect 399 459 402 462 
rect 399 462 402 465 
rect 399 465 402 468 
rect 399 468 402 471 
rect 399 471 402 474 
rect 399 474 402 477 
rect 399 477 402 480 
rect 399 480 402 483 
rect 399 483 402 486 
rect 399 486 402 489 
rect 399 489 402 492 
rect 399 492 402 495 
rect 399 495 402 498 
rect 399 498 402 501 
rect 399 501 402 504 
rect 399 504 402 507 
rect 399 507 402 510 
rect 402 0 405 3 
rect 402 3 405 6 
rect 402 6 405 9 
rect 402 9 405 12 
rect 402 12 405 15 
rect 402 15 405 18 
rect 402 18 405 21 
rect 402 21 405 24 
rect 402 24 405 27 
rect 402 27 405 30 
rect 402 30 405 33 
rect 402 33 405 36 
rect 402 36 405 39 
rect 402 39 405 42 
rect 402 42 405 45 
rect 402 45 405 48 
rect 402 48 405 51 
rect 402 51 405 54 
rect 402 54 405 57 
rect 402 57 405 60 
rect 402 60 405 63 
rect 402 63 405 66 
rect 402 66 405 69 
rect 402 69 405 72 
rect 402 72 405 75 
rect 402 75 405 78 
rect 402 78 405 81 
rect 402 81 405 84 
rect 402 84 405 87 
rect 402 87 405 90 
rect 402 90 405 93 
rect 402 93 405 96 
rect 402 96 405 99 
rect 402 99 405 102 
rect 402 102 405 105 
rect 402 105 405 108 
rect 402 108 405 111 
rect 402 111 405 114 
rect 402 114 405 117 
rect 402 117 405 120 
rect 402 120 405 123 
rect 402 123 405 126 
rect 402 126 405 129 
rect 402 129 405 132 
rect 402 132 405 135 
rect 402 135 405 138 
rect 402 138 405 141 
rect 402 141 405 144 
rect 402 144 405 147 
rect 402 147 405 150 
rect 402 150 405 153 
rect 402 153 405 156 
rect 402 156 405 159 
rect 402 159 405 162 
rect 402 162 405 165 
rect 402 165 405 168 
rect 402 168 405 171 
rect 402 171 405 174 
rect 402 174 405 177 
rect 402 177 405 180 
rect 402 180 405 183 
rect 402 183 405 186 
rect 402 186 405 189 
rect 402 189 405 192 
rect 402 192 405 195 
rect 402 195 405 198 
rect 402 198 405 201 
rect 402 201 405 204 
rect 402 204 405 207 
rect 402 207 405 210 
rect 402 210 405 213 
rect 402 213 405 216 
rect 402 216 405 219 
rect 402 219 405 222 
rect 402 222 405 225 
rect 402 225 405 228 
rect 402 228 405 231 
rect 402 231 405 234 
rect 402 234 405 237 
rect 402 237 405 240 
rect 402 240 405 243 
rect 402 243 405 246 
rect 402 246 405 249 
rect 402 249 405 252 
rect 402 252 405 255 
rect 402 255 405 258 
rect 402 258 405 261 
rect 402 261 405 264 
rect 402 264 405 267 
rect 402 267 405 270 
rect 402 270 405 273 
rect 402 273 405 276 
rect 402 276 405 279 
rect 402 279 405 282 
rect 402 282 405 285 
rect 402 285 405 288 
rect 402 288 405 291 
rect 402 291 405 294 
rect 402 294 405 297 
rect 402 297 405 300 
rect 402 300 405 303 
rect 402 303 405 306 
rect 402 306 405 309 
rect 402 309 405 312 
rect 402 312 405 315 
rect 402 315 405 318 
rect 402 318 405 321 
rect 402 321 405 324 
rect 402 324 405 327 
rect 402 327 405 330 
rect 402 330 405 333 
rect 402 333 405 336 
rect 402 336 405 339 
rect 402 339 405 342 
rect 402 342 405 345 
rect 402 345 405 348 
rect 402 348 405 351 
rect 402 351 405 354 
rect 402 354 405 357 
rect 402 357 405 360 
rect 402 360 405 363 
rect 402 363 405 366 
rect 402 366 405 369 
rect 402 369 405 372 
rect 402 372 405 375 
rect 402 375 405 378 
rect 402 378 405 381 
rect 402 381 405 384 
rect 402 384 405 387 
rect 402 387 405 390 
rect 402 390 405 393 
rect 402 393 405 396 
rect 402 396 405 399 
rect 402 399 405 402 
rect 402 402 405 405 
rect 402 405 405 408 
rect 402 408 405 411 
rect 402 411 405 414 
rect 402 414 405 417 
rect 402 417 405 420 
rect 402 420 405 423 
rect 402 423 405 426 
rect 402 426 405 429 
rect 402 429 405 432 
rect 402 432 405 435 
rect 402 435 405 438 
rect 402 438 405 441 
rect 402 441 405 444 
rect 402 444 405 447 
rect 402 447 405 450 
rect 402 450 405 453 
rect 402 453 405 456 
rect 402 456 405 459 
rect 402 459 405 462 
rect 402 462 405 465 
rect 402 465 405 468 
rect 402 468 405 471 
rect 402 471 405 474 
rect 402 474 405 477 
rect 402 477 405 480 
rect 402 480 405 483 
rect 402 483 405 486 
rect 402 486 405 489 
rect 402 489 405 492 
rect 402 492 405 495 
rect 402 495 405 498 
rect 402 498 405 501 
rect 402 501 405 504 
rect 402 504 405 507 
rect 402 507 405 510 
rect 405 0 408 3 
rect 405 3 408 6 
rect 405 6 408 9 
rect 405 9 408 12 
rect 405 12 408 15 
rect 405 15 408 18 
rect 405 18 408 21 
rect 405 21 408 24 
rect 405 24 408 27 
rect 405 27 408 30 
rect 405 30 408 33 
rect 405 33 408 36 
rect 405 36 408 39 
rect 405 39 408 42 
rect 405 42 408 45 
rect 405 45 408 48 
rect 405 48 408 51 
rect 405 51 408 54 
rect 405 54 408 57 
rect 405 57 408 60 
rect 405 60 408 63 
rect 405 63 408 66 
rect 405 66 408 69 
rect 405 69 408 72 
rect 405 72 408 75 
rect 405 75 408 78 
rect 405 78 408 81 
rect 405 81 408 84 
rect 405 84 408 87 
rect 405 87 408 90 
rect 405 90 408 93 
rect 405 93 408 96 
rect 405 96 408 99 
rect 405 99 408 102 
rect 405 102 408 105 
rect 405 105 408 108 
rect 405 108 408 111 
rect 405 111 408 114 
rect 405 114 408 117 
rect 405 117 408 120 
rect 405 120 408 123 
rect 405 123 408 126 
rect 405 126 408 129 
rect 405 129 408 132 
rect 405 132 408 135 
rect 405 135 408 138 
rect 405 138 408 141 
rect 405 141 408 144 
rect 405 144 408 147 
rect 405 147 408 150 
rect 405 150 408 153 
rect 405 153 408 156 
rect 405 156 408 159 
rect 405 159 408 162 
rect 405 162 408 165 
rect 405 165 408 168 
rect 405 168 408 171 
rect 405 171 408 174 
rect 405 174 408 177 
rect 405 177 408 180 
rect 405 180 408 183 
rect 405 183 408 186 
rect 405 186 408 189 
rect 405 189 408 192 
rect 405 192 408 195 
rect 405 195 408 198 
rect 405 198 408 201 
rect 405 201 408 204 
rect 405 204 408 207 
rect 405 207 408 210 
rect 405 210 408 213 
rect 405 213 408 216 
rect 405 216 408 219 
rect 405 219 408 222 
rect 405 222 408 225 
rect 405 225 408 228 
rect 405 228 408 231 
rect 405 231 408 234 
rect 405 234 408 237 
rect 405 237 408 240 
rect 405 240 408 243 
rect 405 243 408 246 
rect 405 246 408 249 
rect 405 249 408 252 
rect 405 252 408 255 
rect 405 255 408 258 
rect 405 258 408 261 
rect 405 261 408 264 
rect 405 264 408 267 
rect 405 267 408 270 
rect 405 270 408 273 
rect 405 273 408 276 
rect 405 276 408 279 
rect 405 279 408 282 
rect 405 282 408 285 
rect 405 285 408 288 
rect 405 288 408 291 
rect 405 291 408 294 
rect 405 294 408 297 
rect 405 297 408 300 
rect 405 300 408 303 
rect 405 303 408 306 
rect 405 306 408 309 
rect 405 309 408 312 
rect 405 312 408 315 
rect 405 315 408 318 
rect 405 318 408 321 
rect 405 321 408 324 
rect 405 324 408 327 
rect 405 327 408 330 
rect 405 330 408 333 
rect 405 333 408 336 
rect 405 336 408 339 
rect 405 339 408 342 
rect 405 342 408 345 
rect 405 345 408 348 
rect 405 348 408 351 
rect 405 351 408 354 
rect 405 354 408 357 
rect 405 357 408 360 
rect 405 360 408 363 
rect 405 363 408 366 
rect 405 366 408 369 
rect 405 369 408 372 
rect 405 372 408 375 
rect 405 375 408 378 
rect 405 378 408 381 
rect 405 381 408 384 
rect 405 384 408 387 
rect 405 387 408 390 
rect 405 390 408 393 
rect 405 393 408 396 
rect 405 396 408 399 
rect 405 399 408 402 
rect 405 402 408 405 
rect 405 405 408 408 
rect 405 408 408 411 
rect 405 411 408 414 
rect 405 414 408 417 
rect 405 417 408 420 
rect 405 420 408 423 
rect 405 423 408 426 
rect 405 426 408 429 
rect 405 429 408 432 
rect 405 432 408 435 
rect 405 435 408 438 
rect 405 438 408 441 
rect 405 441 408 444 
rect 405 444 408 447 
rect 405 447 408 450 
rect 405 450 408 453 
rect 405 453 408 456 
rect 405 456 408 459 
rect 405 459 408 462 
rect 405 462 408 465 
rect 405 465 408 468 
rect 405 468 408 471 
rect 405 471 408 474 
rect 405 474 408 477 
rect 405 477 408 480 
rect 405 480 408 483 
rect 405 483 408 486 
rect 405 486 408 489 
rect 405 489 408 492 
rect 405 492 408 495 
rect 405 495 408 498 
rect 405 498 408 501 
rect 405 501 408 504 
rect 405 504 408 507 
rect 405 507 408 510 
rect 408 0 411 3 
rect 408 3 411 6 
rect 408 6 411 9 
rect 408 9 411 12 
rect 408 12 411 15 
rect 408 15 411 18 
rect 408 18 411 21 
rect 408 21 411 24 
rect 408 24 411 27 
rect 408 27 411 30 
rect 408 30 411 33 
rect 408 33 411 36 
rect 408 36 411 39 
rect 408 39 411 42 
rect 408 42 411 45 
rect 408 45 411 48 
rect 408 48 411 51 
rect 408 51 411 54 
rect 408 54 411 57 
rect 408 57 411 60 
rect 408 60 411 63 
rect 408 63 411 66 
rect 408 66 411 69 
rect 408 69 411 72 
rect 408 72 411 75 
rect 408 75 411 78 
rect 408 78 411 81 
rect 408 81 411 84 
rect 408 84 411 87 
rect 408 87 411 90 
rect 408 90 411 93 
rect 408 93 411 96 
rect 408 96 411 99 
rect 408 99 411 102 
rect 408 102 411 105 
rect 408 105 411 108 
rect 408 108 411 111 
rect 408 111 411 114 
rect 408 114 411 117 
rect 408 117 411 120 
rect 408 120 411 123 
rect 408 123 411 126 
rect 408 126 411 129 
rect 408 129 411 132 
rect 408 132 411 135 
rect 408 135 411 138 
rect 408 138 411 141 
rect 408 141 411 144 
rect 408 144 411 147 
rect 408 147 411 150 
rect 408 150 411 153 
rect 408 153 411 156 
rect 408 156 411 159 
rect 408 159 411 162 
rect 408 162 411 165 
rect 408 165 411 168 
rect 408 168 411 171 
rect 408 171 411 174 
rect 408 174 411 177 
rect 408 177 411 180 
rect 408 180 411 183 
rect 408 183 411 186 
rect 408 186 411 189 
rect 408 189 411 192 
rect 408 192 411 195 
rect 408 195 411 198 
rect 408 198 411 201 
rect 408 201 411 204 
rect 408 204 411 207 
rect 408 207 411 210 
rect 408 210 411 213 
rect 408 213 411 216 
rect 408 216 411 219 
rect 408 219 411 222 
rect 408 222 411 225 
rect 408 225 411 228 
rect 408 228 411 231 
rect 408 231 411 234 
rect 408 234 411 237 
rect 408 237 411 240 
rect 408 240 411 243 
rect 408 243 411 246 
rect 408 246 411 249 
rect 408 249 411 252 
rect 408 252 411 255 
rect 408 255 411 258 
rect 408 258 411 261 
rect 408 261 411 264 
rect 408 264 411 267 
rect 408 267 411 270 
rect 408 270 411 273 
rect 408 273 411 276 
rect 408 276 411 279 
rect 408 279 411 282 
rect 408 282 411 285 
rect 408 285 411 288 
rect 408 288 411 291 
rect 408 291 411 294 
rect 408 294 411 297 
rect 408 297 411 300 
rect 408 300 411 303 
rect 408 303 411 306 
rect 408 306 411 309 
rect 408 309 411 312 
rect 408 312 411 315 
rect 408 315 411 318 
rect 408 318 411 321 
rect 408 321 411 324 
rect 408 324 411 327 
rect 408 327 411 330 
rect 408 330 411 333 
rect 408 333 411 336 
rect 408 336 411 339 
rect 408 339 411 342 
rect 408 342 411 345 
rect 408 345 411 348 
rect 408 348 411 351 
rect 408 351 411 354 
rect 408 354 411 357 
rect 408 357 411 360 
rect 408 360 411 363 
rect 408 363 411 366 
rect 408 366 411 369 
rect 408 369 411 372 
rect 408 372 411 375 
rect 408 375 411 378 
rect 408 378 411 381 
rect 408 381 411 384 
rect 408 384 411 387 
rect 408 387 411 390 
rect 408 390 411 393 
rect 408 393 411 396 
rect 408 396 411 399 
rect 408 399 411 402 
rect 408 402 411 405 
rect 408 405 411 408 
rect 408 408 411 411 
rect 408 411 411 414 
rect 408 414 411 417 
rect 408 417 411 420 
rect 408 420 411 423 
rect 408 423 411 426 
rect 408 426 411 429 
rect 408 429 411 432 
rect 408 432 411 435 
rect 408 435 411 438 
rect 408 438 411 441 
rect 408 441 411 444 
rect 408 444 411 447 
rect 408 447 411 450 
rect 408 450 411 453 
rect 408 453 411 456 
rect 408 456 411 459 
rect 408 459 411 462 
rect 408 462 411 465 
rect 408 465 411 468 
rect 408 468 411 471 
rect 408 471 411 474 
rect 408 474 411 477 
rect 408 477 411 480 
rect 408 480 411 483 
rect 408 483 411 486 
rect 408 486 411 489 
rect 408 489 411 492 
rect 408 492 411 495 
rect 408 495 411 498 
rect 408 498 411 501 
rect 408 501 411 504 
rect 408 504 411 507 
rect 408 507 411 510 
rect 411 0 414 3 
rect 411 3 414 6 
rect 411 6 414 9 
rect 411 9 414 12 
rect 411 12 414 15 
rect 411 15 414 18 
rect 411 18 414 21 
rect 411 21 414 24 
rect 411 24 414 27 
rect 411 27 414 30 
rect 411 30 414 33 
rect 411 33 414 36 
rect 411 36 414 39 
rect 411 39 414 42 
rect 411 42 414 45 
rect 411 45 414 48 
rect 411 48 414 51 
rect 411 51 414 54 
rect 411 54 414 57 
rect 411 57 414 60 
rect 411 60 414 63 
rect 411 63 414 66 
rect 411 66 414 69 
rect 411 69 414 72 
rect 411 72 414 75 
rect 411 75 414 78 
rect 411 78 414 81 
rect 411 81 414 84 
rect 411 84 414 87 
rect 411 87 414 90 
rect 411 90 414 93 
rect 411 93 414 96 
rect 411 96 414 99 
rect 411 99 414 102 
rect 411 102 414 105 
rect 411 105 414 108 
rect 411 108 414 111 
rect 411 111 414 114 
rect 411 114 414 117 
rect 411 117 414 120 
rect 411 120 414 123 
rect 411 123 414 126 
rect 411 126 414 129 
rect 411 129 414 132 
rect 411 132 414 135 
rect 411 135 414 138 
rect 411 138 414 141 
rect 411 141 414 144 
rect 411 144 414 147 
rect 411 147 414 150 
rect 411 150 414 153 
rect 411 153 414 156 
rect 411 156 414 159 
rect 411 159 414 162 
rect 411 162 414 165 
rect 411 165 414 168 
rect 411 168 414 171 
rect 411 171 414 174 
rect 411 174 414 177 
rect 411 177 414 180 
rect 411 180 414 183 
rect 411 183 414 186 
rect 411 186 414 189 
rect 411 189 414 192 
rect 411 192 414 195 
rect 411 195 414 198 
rect 411 198 414 201 
rect 411 201 414 204 
rect 411 204 414 207 
rect 411 207 414 210 
rect 411 210 414 213 
rect 411 213 414 216 
rect 411 216 414 219 
rect 411 219 414 222 
rect 411 222 414 225 
rect 411 225 414 228 
rect 411 228 414 231 
rect 411 231 414 234 
rect 411 234 414 237 
rect 411 237 414 240 
rect 411 240 414 243 
rect 411 243 414 246 
rect 411 246 414 249 
rect 411 249 414 252 
rect 411 252 414 255 
rect 411 255 414 258 
rect 411 258 414 261 
rect 411 261 414 264 
rect 411 264 414 267 
rect 411 267 414 270 
rect 411 270 414 273 
rect 411 273 414 276 
rect 411 276 414 279 
rect 411 279 414 282 
rect 411 282 414 285 
rect 411 285 414 288 
rect 411 288 414 291 
rect 411 291 414 294 
rect 411 294 414 297 
rect 411 297 414 300 
rect 411 300 414 303 
rect 411 303 414 306 
rect 411 306 414 309 
rect 411 309 414 312 
rect 411 312 414 315 
rect 411 315 414 318 
rect 411 318 414 321 
rect 411 321 414 324 
rect 411 324 414 327 
rect 411 327 414 330 
rect 411 330 414 333 
rect 411 333 414 336 
rect 411 336 414 339 
rect 411 339 414 342 
rect 411 342 414 345 
rect 411 345 414 348 
rect 411 348 414 351 
rect 411 351 414 354 
rect 411 354 414 357 
rect 411 357 414 360 
rect 411 360 414 363 
rect 411 363 414 366 
rect 411 366 414 369 
rect 411 369 414 372 
rect 411 372 414 375 
rect 411 375 414 378 
rect 411 378 414 381 
rect 411 381 414 384 
rect 411 384 414 387 
rect 411 387 414 390 
rect 411 390 414 393 
rect 411 393 414 396 
rect 411 396 414 399 
rect 411 399 414 402 
rect 411 402 414 405 
rect 411 405 414 408 
rect 411 408 414 411 
rect 411 411 414 414 
rect 411 414 414 417 
rect 411 417 414 420 
rect 411 420 414 423 
rect 411 423 414 426 
rect 411 426 414 429 
rect 411 429 414 432 
rect 411 432 414 435 
rect 411 435 414 438 
rect 411 438 414 441 
rect 411 441 414 444 
rect 411 444 414 447 
rect 411 447 414 450 
rect 411 450 414 453 
rect 411 453 414 456 
rect 411 456 414 459 
rect 411 459 414 462 
rect 411 462 414 465 
rect 411 465 414 468 
rect 411 468 414 471 
rect 411 471 414 474 
rect 411 474 414 477 
rect 411 477 414 480 
rect 411 480 414 483 
rect 411 483 414 486 
rect 411 486 414 489 
rect 411 489 414 492 
rect 411 492 414 495 
rect 411 495 414 498 
rect 411 498 414 501 
rect 411 501 414 504 
rect 411 504 414 507 
rect 411 507 414 510 
rect 414 0 417 3 
rect 414 3 417 6 
rect 414 6 417 9 
rect 414 9 417 12 
rect 414 12 417 15 
rect 414 15 417 18 
rect 414 18 417 21 
rect 414 21 417 24 
rect 414 24 417 27 
rect 414 27 417 30 
rect 414 30 417 33 
rect 414 33 417 36 
rect 414 36 417 39 
rect 414 39 417 42 
rect 414 42 417 45 
rect 414 45 417 48 
rect 414 48 417 51 
rect 414 51 417 54 
rect 414 54 417 57 
rect 414 57 417 60 
rect 414 60 417 63 
rect 414 63 417 66 
rect 414 66 417 69 
rect 414 69 417 72 
rect 414 72 417 75 
rect 414 75 417 78 
rect 414 78 417 81 
rect 414 81 417 84 
rect 414 84 417 87 
rect 414 87 417 90 
rect 414 90 417 93 
rect 414 93 417 96 
rect 414 96 417 99 
rect 414 99 417 102 
rect 414 102 417 105 
rect 414 105 417 108 
rect 414 108 417 111 
rect 414 111 417 114 
rect 414 114 417 117 
rect 414 117 417 120 
rect 414 120 417 123 
rect 414 123 417 126 
rect 414 126 417 129 
rect 414 129 417 132 
rect 414 132 417 135 
rect 414 135 417 138 
rect 414 138 417 141 
rect 414 141 417 144 
rect 414 144 417 147 
rect 414 147 417 150 
rect 414 150 417 153 
rect 414 153 417 156 
rect 414 156 417 159 
rect 414 159 417 162 
rect 414 162 417 165 
rect 414 165 417 168 
rect 414 168 417 171 
rect 414 171 417 174 
rect 414 174 417 177 
rect 414 177 417 180 
rect 414 180 417 183 
rect 414 183 417 186 
rect 414 186 417 189 
rect 414 189 417 192 
rect 414 192 417 195 
rect 414 195 417 198 
rect 414 198 417 201 
rect 414 201 417 204 
rect 414 204 417 207 
rect 414 207 417 210 
rect 414 210 417 213 
rect 414 213 417 216 
rect 414 216 417 219 
rect 414 219 417 222 
rect 414 222 417 225 
rect 414 225 417 228 
rect 414 228 417 231 
rect 414 231 417 234 
rect 414 234 417 237 
rect 414 237 417 240 
rect 414 240 417 243 
rect 414 243 417 246 
rect 414 246 417 249 
rect 414 249 417 252 
rect 414 252 417 255 
rect 414 255 417 258 
rect 414 258 417 261 
rect 414 261 417 264 
rect 414 264 417 267 
rect 414 267 417 270 
rect 414 270 417 273 
rect 414 273 417 276 
rect 414 276 417 279 
rect 414 279 417 282 
rect 414 282 417 285 
rect 414 285 417 288 
rect 414 288 417 291 
rect 414 291 417 294 
rect 414 294 417 297 
rect 414 297 417 300 
rect 414 300 417 303 
rect 414 303 417 306 
rect 414 306 417 309 
rect 414 309 417 312 
rect 414 312 417 315 
rect 414 315 417 318 
rect 414 318 417 321 
rect 414 321 417 324 
rect 414 324 417 327 
rect 414 327 417 330 
rect 414 330 417 333 
rect 414 333 417 336 
rect 414 336 417 339 
rect 414 339 417 342 
rect 414 342 417 345 
rect 414 345 417 348 
rect 414 348 417 351 
rect 414 351 417 354 
rect 414 354 417 357 
rect 414 357 417 360 
rect 414 360 417 363 
rect 414 363 417 366 
rect 414 366 417 369 
rect 414 372 417 375 
rect 414 375 417 378 
rect 414 378 417 381 
rect 414 381 417 384 
rect 414 384 417 387 
rect 414 387 417 390 
rect 414 390 417 393 
rect 414 393 417 396 
rect 414 396 417 399 
rect 414 399 417 402 
rect 414 402 417 405 
rect 414 405 417 408 
rect 414 408 417 411 
rect 414 411 417 414 
rect 414 414 417 417 
rect 414 417 417 420 
rect 414 420 417 423 
rect 414 423 417 426 
rect 414 426 417 429 
rect 414 429 417 432 
rect 414 432 417 435 
rect 414 435 417 438 
rect 414 438 417 441 
rect 414 441 417 444 
rect 414 444 417 447 
rect 414 447 417 450 
rect 414 450 417 453 
rect 414 453 417 456 
rect 414 456 417 459 
rect 414 459 417 462 
rect 414 462 417 465 
rect 414 465 417 468 
rect 414 468 417 471 
rect 414 471 417 474 
rect 414 474 417 477 
rect 414 477 417 480 
rect 414 480 417 483 
rect 414 483 417 486 
rect 414 486 417 489 
rect 414 489 417 492 
rect 414 492 417 495 
rect 414 495 417 498 
rect 414 498 417 501 
rect 414 501 417 504 
rect 414 504 417 507 
rect 414 507 417 510 
rect 417 0 420 3 
rect 417 3 420 6 
rect 417 6 420 9 
rect 417 9 420 12 
rect 417 12 420 15 
rect 417 15 420 18 
rect 417 18 420 21 
rect 417 21 420 24 
rect 417 24 420 27 
rect 417 27 420 30 
rect 417 30 420 33 
rect 417 33 420 36 
rect 417 36 420 39 
rect 417 39 420 42 
rect 417 42 420 45 
rect 417 45 420 48 
rect 417 48 420 51 
rect 417 51 420 54 
rect 417 54 420 57 
rect 417 57 420 60 
rect 417 60 420 63 
rect 417 63 420 66 
rect 417 66 420 69 
rect 417 69 420 72 
rect 417 72 420 75 
rect 417 75 420 78 
rect 417 78 420 81 
rect 417 81 420 84 
rect 417 84 420 87 
rect 417 87 420 90 
rect 417 90 420 93 
rect 417 93 420 96 
rect 417 96 420 99 
rect 417 99 420 102 
rect 417 102 420 105 
rect 417 105 420 108 
rect 417 108 420 111 
rect 417 111 420 114 
rect 417 114 420 117 
rect 417 117 420 120 
rect 417 120 420 123 
rect 417 123 420 126 
rect 417 126 420 129 
rect 417 129 420 132 
rect 417 132 420 135 
rect 417 135 420 138 
rect 417 138 420 141 
rect 417 141 420 144 
rect 417 144 420 147 
rect 417 147 420 150 
rect 417 150 420 153 
rect 417 153 420 156 
rect 417 156 420 159 
rect 417 159 420 162 
rect 417 162 420 165 
rect 417 165 420 168 
rect 417 168 420 171 
rect 417 171 420 174 
rect 417 174 420 177 
rect 417 177 420 180 
rect 417 180 420 183 
rect 417 183 420 186 
rect 417 186 420 189 
rect 417 189 420 192 
rect 417 192 420 195 
rect 417 195 420 198 
rect 417 198 420 201 
rect 417 201 420 204 
rect 417 204 420 207 
rect 417 207 420 210 
rect 417 210 420 213 
rect 417 213 420 216 
rect 417 216 420 219 
rect 417 219 420 222 
rect 417 222 420 225 
rect 417 225 420 228 
rect 417 228 420 231 
rect 417 231 420 234 
rect 417 234 420 237 
rect 417 237 420 240 
rect 417 240 420 243 
rect 417 243 420 246 
rect 417 246 420 249 
rect 417 249 420 252 
rect 417 252 420 255 
rect 417 255 420 258 
rect 417 258 420 261 
rect 417 261 420 264 
rect 417 264 420 267 
rect 417 267 420 270 
rect 417 270 420 273 
rect 417 273 420 276 
rect 417 276 420 279 
rect 417 279 420 282 
rect 417 282 420 285 
rect 417 285 420 288 
rect 417 288 420 291 
rect 417 291 420 294 
rect 417 294 420 297 
rect 417 297 420 300 
rect 417 300 420 303 
rect 417 303 420 306 
rect 417 306 420 309 
rect 417 309 420 312 
rect 417 312 420 315 
rect 417 315 420 318 
rect 417 318 420 321 
rect 417 321 420 324 
rect 417 324 420 327 
rect 417 327 420 330 
rect 417 330 420 333 
rect 417 333 420 336 
rect 417 336 420 339 
rect 417 339 420 342 
rect 417 342 420 345 
rect 417 345 420 348 
rect 417 348 420 351 
rect 417 351 420 354 
rect 417 354 420 357 
rect 417 357 420 360 
rect 417 360 420 363 
rect 417 363 420 366 
rect 417 366 420 369 
rect 417 369 420 372 
rect 417 372 420 375 
rect 417 375 420 378 
rect 417 378 420 381 
rect 417 381 420 384 
rect 417 384 420 387 
rect 417 387 420 390 
rect 417 390 420 393 
rect 417 393 420 396 
rect 417 396 420 399 
rect 417 399 420 402 
rect 417 402 420 405 
rect 417 405 420 408 
rect 417 408 420 411 
rect 417 411 420 414 
rect 417 414 420 417 
rect 417 417 420 420 
rect 417 420 420 423 
rect 417 423 420 426 
rect 417 426 420 429 
rect 417 429 420 432 
rect 417 432 420 435 
rect 417 435 420 438 
rect 417 438 420 441 
rect 417 441 420 444 
rect 417 444 420 447 
rect 417 447 420 450 
rect 417 450 420 453 
rect 417 453 420 456 
rect 417 456 420 459 
rect 417 459 420 462 
rect 417 462 420 465 
rect 417 465 420 468 
rect 417 468 420 471 
rect 417 471 420 474 
rect 417 474 420 477 
rect 417 477 420 480 
rect 417 480 420 483 
rect 417 483 420 486 
rect 417 486 420 489 
rect 417 489 420 492 
rect 417 492 420 495 
rect 417 495 420 498 
rect 417 498 420 501 
rect 417 501 420 504 
rect 417 504 420 507 
rect 417 507 420 510 
rect 420 0 423 3 
rect 420 3 423 6 
rect 420 6 423 9 
rect 420 9 423 12 
rect 420 12 423 15 
rect 420 15 423 18 
rect 420 18 423 21 
rect 420 21 423 24 
rect 420 24 423 27 
rect 420 27 423 30 
rect 420 30 423 33 
rect 420 33 423 36 
rect 420 36 423 39 
rect 420 39 423 42 
rect 420 42 423 45 
rect 420 45 423 48 
rect 420 48 423 51 
rect 420 51 423 54 
rect 420 54 423 57 
rect 420 57 423 60 
rect 420 60 423 63 
rect 420 63 423 66 
rect 420 66 423 69 
rect 420 69 423 72 
rect 420 72 423 75 
rect 420 75 423 78 
rect 420 78 423 81 
rect 420 81 423 84 
rect 420 84 423 87 
rect 420 87 423 90 
rect 420 90 423 93 
rect 420 93 423 96 
rect 420 96 423 99 
rect 420 99 423 102 
rect 420 102 423 105 
rect 420 105 423 108 
rect 420 108 423 111 
rect 420 111 423 114 
rect 420 114 423 117 
rect 420 117 423 120 
rect 420 120 423 123 
rect 420 123 423 126 
rect 420 126 423 129 
rect 420 129 423 132 
rect 420 132 423 135 
rect 420 135 423 138 
rect 420 138 423 141 
rect 420 141 423 144 
rect 420 144 423 147 
rect 420 147 423 150 
rect 420 150 423 153 
rect 420 153 423 156 
rect 420 156 423 159 
rect 420 159 423 162 
rect 420 162 423 165 
rect 420 165 423 168 
rect 420 168 423 171 
rect 420 171 423 174 
rect 420 174 423 177 
rect 420 177 423 180 
rect 420 180 423 183 
rect 420 183 423 186 
rect 420 186 423 189 
rect 420 189 423 192 
rect 420 192 423 195 
rect 420 195 423 198 
rect 420 198 423 201 
rect 420 201 423 204 
rect 420 204 423 207 
rect 420 207 423 210 
rect 420 210 423 213 
rect 420 213 423 216 
rect 420 216 423 219 
rect 420 219 423 222 
rect 420 222 423 225 
rect 420 225 423 228 
rect 420 228 423 231 
rect 420 231 423 234 
rect 420 234 423 237 
rect 420 237 423 240 
rect 420 240 423 243 
rect 420 243 423 246 
rect 420 246 423 249 
rect 420 249 423 252 
rect 420 252 423 255 
rect 420 255 423 258 
rect 420 258 423 261 
rect 420 261 423 264 
rect 420 264 423 267 
rect 420 267 423 270 
rect 420 270 423 273 
rect 420 273 423 276 
rect 420 276 423 279 
rect 420 279 423 282 
rect 420 282 423 285 
rect 420 285 423 288 
rect 420 288 423 291 
rect 420 291 423 294 
rect 420 294 423 297 
rect 420 297 423 300 
rect 420 300 423 303 
rect 420 303 423 306 
rect 420 306 423 309 
rect 420 309 423 312 
rect 420 312 423 315 
rect 420 315 423 318 
rect 420 318 423 321 
rect 420 321 423 324 
rect 420 324 423 327 
rect 420 327 423 330 
rect 420 330 423 333 
rect 420 333 423 336 
rect 420 336 423 339 
rect 420 339 423 342 
rect 420 342 423 345 
rect 420 345 423 348 
rect 420 348 423 351 
rect 420 351 423 354 
rect 420 354 423 357 
rect 420 357 423 360 
rect 420 360 423 363 
rect 420 363 423 366 
rect 420 366 423 369 
rect 420 369 423 372 
rect 420 372 423 375 
rect 420 375 423 378 
rect 420 378 423 381 
rect 420 381 423 384 
rect 420 384 423 387 
rect 420 387 423 390 
rect 420 390 423 393 
rect 420 393 423 396 
rect 420 396 423 399 
rect 420 399 423 402 
rect 420 402 423 405 
rect 420 405 423 408 
rect 420 408 423 411 
rect 420 411 423 414 
rect 420 414 423 417 
rect 420 417 423 420 
rect 420 420 423 423 
rect 420 423 423 426 
rect 420 426 423 429 
rect 420 429 423 432 
rect 420 432 423 435 
rect 420 435 423 438 
rect 420 438 423 441 
rect 420 441 423 444 
rect 420 444 423 447 
rect 420 447 423 450 
rect 420 450 423 453 
rect 420 453 423 456 
rect 420 456 423 459 
rect 420 459 423 462 
rect 420 462 423 465 
rect 420 465 423 468 
rect 420 468 423 471 
rect 420 471 423 474 
rect 420 474 423 477 
rect 420 477 423 480 
rect 420 480 423 483 
rect 420 483 423 486 
rect 420 486 423 489 
rect 420 489 423 492 
rect 420 492 423 495 
rect 420 495 423 498 
rect 420 498 423 501 
rect 420 501 423 504 
rect 420 504 423 507 
rect 420 507 423 510 
rect 423 0 426 3 
rect 423 3 426 6 
rect 423 6 426 9 
rect 423 9 426 12 
rect 423 12 426 15 
rect 423 15 426 18 
rect 423 18 426 21 
rect 423 21 426 24 
rect 423 24 426 27 
rect 423 27 426 30 
rect 423 30 426 33 
rect 423 33 426 36 
rect 423 36 426 39 
rect 423 39 426 42 
rect 423 42 426 45 
rect 423 45 426 48 
rect 423 48 426 51 
rect 423 51 426 54 
rect 423 54 426 57 
rect 423 57 426 60 
rect 423 60 426 63 
rect 423 63 426 66 
rect 423 66 426 69 
rect 423 69 426 72 
rect 423 72 426 75 
rect 423 75 426 78 
rect 423 78 426 81 
rect 423 81 426 84 
rect 423 84 426 87 
rect 423 87 426 90 
rect 423 90 426 93 
rect 423 93 426 96 
rect 423 96 426 99 
rect 423 99 426 102 
rect 423 102 426 105 
rect 423 105 426 108 
rect 423 108 426 111 
rect 423 111 426 114 
rect 423 114 426 117 
rect 423 117 426 120 
rect 423 120 426 123 
rect 423 123 426 126 
rect 423 126 426 129 
rect 423 129 426 132 
rect 423 132 426 135 
rect 423 135 426 138 
rect 423 138 426 141 
rect 423 141 426 144 
rect 423 144 426 147 
rect 423 147 426 150 
rect 423 150 426 153 
rect 423 153 426 156 
rect 423 156 426 159 
rect 423 159 426 162 
rect 423 162 426 165 
rect 423 165 426 168 
rect 423 168 426 171 
rect 423 171 426 174 
rect 423 174 426 177 
rect 423 177 426 180 
rect 423 180 426 183 
rect 423 183 426 186 
rect 423 186 426 189 
rect 423 189 426 192 
rect 423 192 426 195 
rect 423 195 426 198 
rect 423 198 426 201 
rect 423 201 426 204 
rect 423 204 426 207 
rect 423 207 426 210 
rect 423 210 426 213 
rect 423 213 426 216 
rect 423 216 426 219 
rect 423 219 426 222 
rect 423 222 426 225 
rect 423 225 426 228 
rect 423 228 426 231 
rect 423 231 426 234 
rect 423 234 426 237 
rect 423 237 426 240 
rect 423 240 426 243 
rect 423 243 426 246 
rect 423 246 426 249 
rect 423 249 426 252 
rect 423 252 426 255 
rect 423 255 426 258 
rect 423 258 426 261 
rect 423 261 426 264 
rect 423 264 426 267 
rect 423 267 426 270 
rect 423 270 426 273 
rect 423 273 426 276 
rect 423 276 426 279 
rect 423 279 426 282 
rect 423 282 426 285 
rect 423 285 426 288 
rect 423 288 426 291 
rect 423 291 426 294 
rect 423 294 426 297 
rect 423 297 426 300 
rect 423 300 426 303 
rect 423 303 426 306 
rect 423 306 426 309 
rect 423 309 426 312 
rect 423 312 426 315 
rect 423 315 426 318 
rect 423 318 426 321 
rect 423 321 426 324 
rect 423 324 426 327 
rect 423 327 426 330 
rect 423 330 426 333 
rect 423 333 426 336 
rect 423 336 426 339 
rect 423 339 426 342 
rect 423 342 426 345 
rect 423 345 426 348 
rect 423 348 426 351 
rect 423 351 426 354 
rect 423 354 426 357 
rect 423 357 426 360 
rect 423 360 426 363 
rect 423 363 426 366 
rect 423 366 426 369 
rect 423 369 426 372 
rect 423 372 426 375 
rect 423 375 426 378 
rect 423 378 426 381 
rect 423 381 426 384 
rect 423 384 426 387 
rect 423 387 426 390 
rect 423 390 426 393 
rect 423 393 426 396 
rect 423 396 426 399 
rect 423 399 426 402 
rect 423 402 426 405 
rect 423 405 426 408 
rect 423 408 426 411 
rect 423 411 426 414 
rect 423 414 426 417 
rect 423 417 426 420 
rect 423 420 426 423 
rect 423 423 426 426 
rect 423 426 426 429 
rect 423 429 426 432 
rect 423 432 426 435 
rect 423 435 426 438 
rect 423 438 426 441 
rect 423 441 426 444 
rect 423 444 426 447 
rect 423 447 426 450 
rect 423 450 426 453 
rect 423 453 426 456 
rect 423 456 426 459 
rect 423 459 426 462 
rect 423 462 426 465 
rect 423 465 426 468 
rect 423 468 426 471 
rect 423 471 426 474 
rect 423 474 426 477 
rect 423 477 426 480 
rect 423 480 426 483 
rect 423 483 426 486 
rect 423 486 426 489 
rect 423 489 426 492 
rect 423 492 426 495 
rect 423 495 426 498 
rect 423 498 426 501 
rect 423 501 426 504 
rect 423 504 426 507 
rect 423 507 426 510 
rect 426 0 429 3 
rect 426 3 429 6 
rect 426 6 429 9 
rect 426 9 429 12 
rect 426 12 429 15 
rect 426 15 429 18 
rect 426 18 429 21 
rect 426 21 429 24 
rect 426 24 429 27 
rect 426 27 429 30 
rect 426 30 429 33 
rect 426 33 429 36 
rect 426 36 429 39 
rect 426 39 429 42 
rect 426 42 429 45 
rect 426 45 429 48 
rect 426 48 429 51 
rect 426 51 429 54 
rect 426 54 429 57 
rect 426 57 429 60 
rect 426 60 429 63 
rect 426 63 429 66 
rect 426 66 429 69 
rect 426 69 429 72 
rect 426 72 429 75 
rect 426 75 429 78 
rect 426 78 429 81 
rect 426 81 429 84 
rect 426 84 429 87 
rect 426 87 429 90 
rect 426 90 429 93 
rect 426 93 429 96 
rect 426 96 429 99 
rect 426 99 429 102 
rect 426 102 429 105 
rect 426 105 429 108 
rect 426 108 429 111 
rect 426 111 429 114 
rect 426 114 429 117 
rect 426 117 429 120 
rect 426 120 429 123 
rect 426 123 429 126 
rect 426 126 429 129 
rect 426 129 429 132 
rect 426 132 429 135 
rect 426 135 429 138 
rect 426 138 429 141 
rect 426 141 429 144 
rect 426 144 429 147 
rect 426 147 429 150 
rect 426 150 429 153 
rect 426 153 429 156 
rect 426 156 429 159 
rect 426 159 429 162 
rect 426 162 429 165 
rect 426 165 429 168 
rect 426 168 429 171 
rect 426 171 429 174 
rect 426 174 429 177 
rect 426 177 429 180 
rect 426 180 429 183 
rect 426 183 429 186 
rect 426 186 429 189 
rect 426 189 429 192 
rect 426 192 429 195 
rect 426 195 429 198 
rect 426 198 429 201 
rect 426 201 429 204 
rect 426 204 429 207 
rect 426 207 429 210 
rect 426 210 429 213 
rect 426 213 429 216 
rect 426 216 429 219 
rect 426 219 429 222 
rect 426 222 429 225 
rect 426 225 429 228 
rect 426 228 429 231 
rect 426 231 429 234 
rect 426 234 429 237 
rect 426 237 429 240 
rect 426 240 429 243 
rect 426 243 429 246 
rect 426 246 429 249 
rect 426 249 429 252 
rect 426 252 429 255 
rect 426 255 429 258 
rect 426 258 429 261 
rect 426 261 429 264 
rect 426 264 429 267 
rect 426 267 429 270 
rect 426 270 429 273 
rect 426 273 429 276 
rect 426 276 429 279 
rect 426 279 429 282 
rect 426 282 429 285 
rect 426 285 429 288 
rect 426 288 429 291 
rect 426 291 429 294 
rect 426 294 429 297 
rect 426 297 429 300 
rect 426 300 429 303 
rect 426 303 429 306 
rect 426 306 429 309 
rect 426 309 429 312 
rect 426 312 429 315 
rect 426 315 429 318 
rect 426 318 429 321 
rect 426 321 429 324 
rect 426 324 429 327 
rect 426 327 429 330 
rect 426 330 429 333 
rect 426 333 429 336 
rect 426 336 429 339 
rect 426 339 429 342 
rect 426 342 429 345 
rect 426 345 429 348 
rect 426 348 429 351 
rect 426 351 429 354 
rect 426 354 429 357 
rect 426 357 429 360 
rect 426 360 429 363 
rect 426 363 429 366 
rect 426 366 429 369 
rect 426 369 429 372 
rect 426 372 429 375 
rect 426 375 429 378 
rect 426 378 429 381 
rect 426 381 429 384 
rect 426 384 429 387 
rect 426 387 429 390 
rect 426 390 429 393 
rect 426 393 429 396 
rect 426 396 429 399 
rect 426 399 429 402 
rect 426 402 429 405 
rect 426 405 429 408 
rect 426 408 429 411 
rect 426 411 429 414 
rect 426 414 429 417 
rect 426 417 429 420 
rect 426 420 429 423 
rect 426 423 429 426 
rect 426 426 429 429 
rect 426 429 429 432 
rect 426 432 429 435 
rect 426 435 429 438 
rect 426 438 429 441 
rect 426 441 429 444 
rect 426 444 429 447 
rect 426 447 429 450 
rect 426 450 429 453 
rect 426 453 429 456 
rect 426 456 429 459 
rect 426 459 429 462 
rect 426 462 429 465 
rect 426 465 429 468 
rect 426 468 429 471 
rect 426 471 429 474 
rect 426 474 429 477 
rect 426 477 429 480 
rect 426 480 429 483 
rect 426 483 429 486 
rect 426 486 429 489 
rect 426 489 429 492 
rect 426 492 429 495 
rect 426 495 429 498 
rect 426 498 429 501 
rect 426 501 429 504 
rect 426 504 429 507 
rect 426 507 429 510 
rect 429 0 432 3 
rect 429 3 432 6 
rect 429 6 432 9 
rect 429 9 432 12 
rect 429 12 432 15 
rect 429 15 432 18 
rect 429 18 432 21 
rect 429 21 432 24 
rect 429 24 432 27 
rect 429 27 432 30 
rect 429 30 432 33 
rect 429 33 432 36 
rect 429 36 432 39 
rect 429 39 432 42 
rect 429 45 432 48 
rect 429 48 432 51 
rect 429 51 432 54 
rect 429 54 432 57 
rect 429 57 432 60 
rect 429 60 432 63 
rect 429 63 432 66 
rect 429 66 432 69 
rect 429 69 432 72 
rect 429 72 432 75 
rect 429 75 432 78 
rect 429 78 432 81 
rect 429 81 432 84 
rect 429 84 432 87 
rect 429 87 432 90 
rect 429 90 432 93 
rect 429 93 432 96 
rect 429 96 432 99 
rect 429 99 432 102 
rect 429 102 432 105 
rect 429 105 432 108 
rect 429 108 432 111 
rect 429 111 432 114 
rect 429 114 432 117 
rect 429 117 432 120 
rect 429 120 432 123 
rect 429 123 432 126 
rect 429 126 432 129 
rect 429 132 432 135 
rect 429 135 432 138 
rect 429 138 432 141 
rect 429 141 432 144 
rect 429 144 432 147 
rect 429 147 432 150 
rect 429 150 432 153 
rect 429 153 432 156 
rect 429 156 432 159 
rect 429 159 432 162 
rect 429 162 432 165 
rect 429 165 432 168 
rect 429 168 432 171 
rect 429 171 432 174 
rect 429 174 432 177 
rect 429 177 432 180 
rect 429 180 432 183 
rect 429 183 432 186 
rect 429 186 432 189 
rect 429 189 432 192 
rect 429 192 432 195 
rect 429 195 432 198 
rect 429 198 432 201 
rect 429 201 432 204 
rect 429 204 432 207 
rect 429 207 432 210 
rect 429 210 432 213 
rect 429 213 432 216 
rect 429 216 432 219 
rect 429 219 432 222 
rect 429 222 432 225 
rect 429 225 432 228 
rect 429 228 432 231 
rect 429 231 432 234 
rect 429 234 432 237 
rect 429 237 432 240 
rect 429 240 432 243 
rect 429 243 432 246 
rect 429 246 432 249 
rect 429 249 432 252 
rect 429 252 432 255 
rect 429 255 432 258 
rect 429 258 432 261 
rect 429 261 432 264 
rect 429 264 432 267 
rect 429 267 432 270 
rect 429 270 432 273 
rect 429 273 432 276 
rect 429 276 432 279 
rect 429 279 432 282 
rect 429 282 432 285 
rect 429 285 432 288 
rect 429 288 432 291 
rect 429 291 432 294 
rect 429 294 432 297 
rect 429 297 432 300 
rect 429 300 432 303 
rect 429 303 432 306 
rect 429 306 432 309 
rect 429 309 432 312 
rect 429 312 432 315 
rect 429 315 432 318 
rect 429 318 432 321 
rect 429 324 432 327 
rect 429 327 432 330 
rect 429 330 432 333 
rect 429 333 432 336 
rect 429 336 432 339 
rect 429 339 432 342 
rect 429 342 432 345 
rect 429 345 432 348 
rect 429 348 432 351 
rect 429 351 432 354 
rect 429 354 432 357 
rect 429 357 432 360 
rect 429 360 432 363 
rect 429 363 432 366 
rect 429 366 432 369 
rect 429 369 432 372 
rect 429 372 432 375 
rect 429 375 432 378 
rect 429 378 432 381 
rect 429 381 432 384 
rect 429 384 432 387 
rect 429 387 432 390 
rect 429 390 432 393 
rect 429 393 432 396 
rect 429 396 432 399 
rect 429 399 432 402 
rect 429 402 432 405 
rect 429 405 432 408 
rect 429 408 432 411 
rect 429 411 432 414 
rect 429 414 432 417 
rect 429 417 432 420 
rect 429 420 432 423 
rect 429 423 432 426 
rect 429 429 432 432 
rect 429 432 432 435 
rect 429 435 432 438 
rect 429 438 432 441 
rect 429 441 432 444 
rect 429 444 432 447 
rect 429 447 432 450 
rect 429 450 432 453 
rect 429 453 432 456 
rect 429 456 432 459 
rect 429 459 432 462 
rect 429 462 432 465 
rect 429 465 432 468 
rect 429 468 432 471 
rect 429 471 432 474 
rect 429 474 432 477 
rect 429 477 432 480 
rect 429 480 432 483 
rect 429 483 432 486 
rect 429 486 432 489 
rect 429 489 432 492 
rect 429 492 432 495 
rect 429 495 432 498 
rect 429 498 432 501 
rect 429 501 432 504 
rect 429 504 432 507 
rect 429 507 432 510 
rect 432 0 435 3 
rect 432 3 435 6 
rect 432 6 435 9 
rect 432 9 435 12 
rect 432 12 435 15 
rect 432 15 435 18 
rect 432 18 435 21 
rect 432 21 435 24 
rect 432 24 435 27 
rect 432 27 435 30 
rect 432 30 435 33 
rect 432 33 435 36 
rect 432 36 435 39 
rect 432 39 435 42 
rect 432 42 435 45 
rect 432 45 435 48 
rect 432 48 435 51 
rect 432 51 435 54 
rect 432 54 435 57 
rect 432 57 435 60 
rect 432 60 435 63 
rect 432 63 435 66 
rect 432 66 435 69 
rect 432 69 435 72 
rect 432 72 435 75 
rect 432 75 435 78 
rect 432 78 435 81 
rect 432 81 435 84 
rect 432 84 435 87 
rect 432 87 435 90 
rect 432 90 435 93 
rect 432 93 435 96 
rect 432 96 435 99 
rect 432 99 435 102 
rect 432 102 435 105 
rect 432 105 435 108 
rect 432 108 435 111 
rect 432 111 435 114 
rect 432 114 435 117 
rect 432 117 435 120 
rect 432 120 435 123 
rect 432 123 435 126 
rect 432 126 435 129 
rect 432 129 435 132 
rect 432 132 435 135 
rect 432 135 435 138 
rect 432 138 435 141 
rect 432 141 435 144 
rect 432 144 435 147 
rect 432 147 435 150 
rect 432 150 435 153 
rect 432 153 435 156 
rect 432 156 435 159 
rect 432 159 435 162 
rect 432 162 435 165 
rect 432 165 435 168 
rect 432 168 435 171 
rect 432 171 435 174 
rect 432 174 435 177 
rect 432 177 435 180 
rect 432 180 435 183 
rect 432 183 435 186 
rect 432 186 435 189 
rect 432 189 435 192 
rect 432 192 435 195 
rect 432 195 435 198 
rect 432 198 435 201 
rect 432 201 435 204 
rect 432 204 435 207 
rect 432 207 435 210 
rect 432 210 435 213 
rect 432 213 435 216 
rect 432 216 435 219 
rect 432 219 435 222 
rect 432 222 435 225 
rect 432 225 435 228 
rect 432 228 435 231 
rect 432 231 435 234 
rect 432 234 435 237 
rect 432 237 435 240 
rect 432 240 435 243 
rect 432 243 435 246 
rect 432 246 435 249 
rect 432 249 435 252 
rect 432 252 435 255 
rect 432 255 435 258 
rect 432 258 435 261 
rect 432 261 435 264 
rect 432 264 435 267 
rect 432 267 435 270 
rect 432 270 435 273 
rect 432 273 435 276 
rect 432 276 435 279 
rect 432 279 435 282 
rect 432 282 435 285 
rect 432 285 435 288 
rect 432 288 435 291 
rect 432 291 435 294 
rect 432 294 435 297 
rect 432 297 435 300 
rect 432 300 435 303 
rect 432 303 435 306 
rect 432 306 435 309 
rect 432 309 435 312 
rect 432 312 435 315 
rect 432 315 435 318 
rect 432 318 435 321 
rect 432 321 435 324 
rect 432 324 435 327 
rect 432 327 435 330 
rect 432 330 435 333 
rect 432 333 435 336 
rect 432 336 435 339 
rect 432 339 435 342 
rect 432 342 435 345 
rect 432 345 435 348 
rect 432 348 435 351 
rect 432 351 435 354 
rect 432 354 435 357 
rect 432 357 435 360 
rect 432 360 435 363 
rect 432 363 435 366 
rect 432 366 435 369 
rect 432 369 435 372 
rect 432 372 435 375 
rect 432 375 435 378 
rect 432 378 435 381 
rect 432 381 435 384 
rect 432 384 435 387 
rect 432 387 435 390 
rect 432 390 435 393 
rect 432 393 435 396 
rect 432 396 435 399 
rect 432 399 435 402 
rect 432 402 435 405 
rect 432 405 435 408 
rect 432 408 435 411 
rect 432 411 435 414 
rect 432 414 435 417 
rect 432 417 435 420 
rect 432 420 435 423 
rect 432 423 435 426 
rect 432 426 435 429 
rect 432 429 435 432 
rect 432 432 435 435 
rect 432 435 435 438 
rect 432 438 435 441 
rect 432 441 435 444 
rect 432 444 435 447 
rect 432 447 435 450 
rect 432 450 435 453 
rect 432 453 435 456 
rect 432 456 435 459 
rect 432 459 435 462 
rect 432 462 435 465 
rect 432 465 435 468 
rect 432 468 435 471 
rect 432 471 435 474 
rect 432 474 435 477 
rect 432 477 435 480 
rect 432 480 435 483 
rect 432 483 435 486 
rect 432 486 435 489 
rect 432 489 435 492 
rect 432 492 435 495 
rect 432 495 435 498 
rect 432 498 435 501 
rect 432 501 435 504 
rect 432 504 435 507 
rect 432 507 435 510 
rect 435 0 438 3 
rect 435 3 438 6 
rect 435 6 438 9 
rect 435 9 438 12 
rect 435 12 438 15 
rect 435 15 438 18 
rect 435 18 438 21 
rect 435 21 438 24 
rect 435 24 438 27 
rect 435 27 438 30 
rect 435 30 438 33 
rect 435 33 438 36 
rect 435 36 438 39 
rect 435 39 438 42 
rect 435 42 438 45 
rect 435 45 438 48 
rect 435 48 438 51 
rect 435 51 438 54 
rect 435 54 438 57 
rect 435 57 438 60 
rect 435 60 438 63 
rect 435 63 438 66 
rect 435 66 438 69 
rect 435 69 438 72 
rect 435 72 438 75 
rect 435 75 438 78 
rect 435 78 438 81 
rect 435 81 438 84 
rect 435 84 438 87 
rect 435 87 438 90 
rect 435 90 438 93 
rect 435 93 438 96 
rect 435 96 438 99 
rect 435 99 438 102 
rect 435 102 438 105 
rect 435 105 438 108 
rect 435 108 438 111 
rect 435 111 438 114 
rect 435 114 438 117 
rect 435 117 438 120 
rect 435 120 438 123 
rect 435 123 438 126 
rect 435 126 438 129 
rect 435 129 438 132 
rect 435 132 438 135 
rect 435 135 438 138 
rect 435 138 438 141 
rect 435 141 438 144 
rect 435 144 438 147 
rect 435 147 438 150 
rect 435 150 438 153 
rect 435 153 438 156 
rect 435 156 438 159 
rect 435 159 438 162 
rect 435 162 438 165 
rect 435 165 438 168 
rect 435 168 438 171 
rect 435 171 438 174 
rect 435 174 438 177 
rect 435 177 438 180 
rect 435 180 438 183 
rect 435 183 438 186 
rect 435 186 438 189 
rect 435 189 438 192 
rect 435 192 438 195 
rect 435 195 438 198 
rect 435 198 438 201 
rect 435 201 438 204 
rect 435 204 438 207 
rect 435 207 438 210 
rect 435 210 438 213 
rect 435 213 438 216 
rect 435 216 438 219 
rect 435 219 438 222 
rect 435 222 438 225 
rect 435 225 438 228 
rect 435 228 438 231 
rect 435 231 438 234 
rect 435 234 438 237 
rect 435 237 438 240 
rect 435 240 438 243 
rect 435 243 438 246 
rect 435 246 438 249 
rect 435 249 438 252 
rect 435 252 438 255 
rect 435 255 438 258 
rect 435 258 438 261 
rect 435 261 438 264 
rect 435 264 438 267 
rect 435 267 438 270 
rect 435 270 438 273 
rect 435 273 438 276 
rect 435 276 438 279 
rect 435 279 438 282 
rect 435 282 438 285 
rect 435 285 438 288 
rect 435 288 438 291 
rect 435 291 438 294 
rect 435 294 438 297 
rect 435 297 438 300 
rect 435 300 438 303 
rect 435 303 438 306 
rect 435 306 438 309 
rect 435 309 438 312 
rect 435 312 438 315 
rect 435 315 438 318 
rect 435 318 438 321 
rect 435 321 438 324 
rect 435 324 438 327 
rect 435 327 438 330 
rect 435 330 438 333 
rect 435 333 438 336 
rect 435 336 438 339 
rect 435 339 438 342 
rect 435 342 438 345 
rect 435 345 438 348 
rect 435 348 438 351 
rect 435 351 438 354 
rect 435 354 438 357 
rect 435 357 438 360 
rect 435 360 438 363 
rect 435 363 438 366 
rect 435 366 438 369 
rect 435 369 438 372 
rect 435 372 438 375 
rect 435 375 438 378 
rect 435 378 438 381 
rect 435 381 438 384 
rect 435 384 438 387 
rect 435 387 438 390 
rect 435 390 438 393 
rect 435 393 438 396 
rect 435 396 438 399 
rect 435 399 438 402 
rect 435 402 438 405 
rect 435 405 438 408 
rect 435 408 438 411 
rect 435 411 438 414 
rect 435 414 438 417 
rect 435 417 438 420 
rect 435 420 438 423 
rect 435 423 438 426 
rect 435 426 438 429 
rect 435 429 438 432 
rect 435 432 438 435 
rect 435 435 438 438 
rect 435 438 438 441 
rect 435 441 438 444 
rect 435 444 438 447 
rect 435 447 438 450 
rect 435 450 438 453 
rect 435 453 438 456 
rect 435 456 438 459 
rect 435 459 438 462 
rect 435 462 438 465 
rect 435 465 438 468 
rect 435 468 438 471 
rect 435 471 438 474 
rect 435 474 438 477 
rect 435 477 438 480 
rect 435 480 438 483 
rect 435 483 438 486 
rect 435 486 438 489 
rect 435 489 438 492 
rect 435 492 438 495 
rect 435 495 438 498 
rect 435 498 438 501 
rect 435 501 438 504 
rect 435 504 438 507 
rect 435 507 438 510 
rect 438 0 441 3 
rect 438 3 441 6 
rect 438 6 441 9 
rect 438 9 441 12 
rect 438 12 441 15 
rect 438 15 441 18 
rect 438 18 441 21 
rect 438 21 441 24 
rect 438 24 441 27 
rect 438 27 441 30 
rect 438 30 441 33 
rect 438 33 441 36 
rect 438 36 441 39 
rect 438 39 441 42 
rect 438 42 441 45 
rect 438 45 441 48 
rect 438 48 441 51 
rect 438 51 441 54 
rect 438 54 441 57 
rect 438 57 441 60 
rect 438 60 441 63 
rect 438 63 441 66 
rect 438 66 441 69 
rect 438 69 441 72 
rect 438 72 441 75 
rect 438 75 441 78 
rect 438 78 441 81 
rect 438 81 441 84 
rect 438 84 441 87 
rect 438 87 441 90 
rect 438 90 441 93 
rect 438 93 441 96 
rect 438 96 441 99 
rect 438 99 441 102 
rect 438 102 441 105 
rect 438 105 441 108 
rect 438 108 441 111 
rect 438 111 441 114 
rect 438 114 441 117 
rect 438 117 441 120 
rect 438 120 441 123 
rect 438 123 441 126 
rect 438 126 441 129 
rect 438 129 441 132 
rect 438 132 441 135 
rect 438 135 441 138 
rect 438 138 441 141 
rect 438 141 441 144 
rect 438 144 441 147 
rect 438 147 441 150 
rect 438 150 441 153 
rect 438 153 441 156 
rect 438 156 441 159 
rect 438 159 441 162 
rect 438 162 441 165 
rect 438 165 441 168 
rect 438 168 441 171 
rect 438 171 441 174 
rect 438 174 441 177 
rect 438 177 441 180 
rect 438 180 441 183 
rect 438 183 441 186 
rect 438 186 441 189 
rect 438 189 441 192 
rect 438 192 441 195 
rect 438 195 441 198 
rect 438 198 441 201 
rect 438 201 441 204 
rect 438 204 441 207 
rect 438 207 441 210 
rect 438 210 441 213 
rect 438 213 441 216 
rect 438 216 441 219 
rect 438 219 441 222 
rect 438 222 441 225 
rect 438 225 441 228 
rect 438 228 441 231 
rect 438 231 441 234 
rect 438 234 441 237 
rect 438 237 441 240 
rect 438 240 441 243 
rect 438 243 441 246 
rect 438 246 441 249 
rect 438 249 441 252 
rect 438 252 441 255 
rect 438 255 441 258 
rect 438 258 441 261 
rect 438 261 441 264 
rect 438 264 441 267 
rect 438 267 441 270 
rect 438 270 441 273 
rect 438 273 441 276 
rect 438 276 441 279 
rect 438 279 441 282 
rect 438 282 441 285 
rect 438 285 441 288 
rect 438 288 441 291 
rect 438 291 441 294 
rect 438 294 441 297 
rect 438 297 441 300 
rect 438 300 441 303 
rect 438 303 441 306 
rect 438 306 441 309 
rect 438 309 441 312 
rect 438 312 441 315 
rect 438 315 441 318 
rect 438 318 441 321 
rect 438 321 441 324 
rect 438 324 441 327 
rect 438 327 441 330 
rect 438 330 441 333 
rect 438 333 441 336 
rect 438 336 441 339 
rect 438 339 441 342 
rect 438 342 441 345 
rect 438 345 441 348 
rect 438 348 441 351 
rect 438 351 441 354 
rect 438 354 441 357 
rect 438 357 441 360 
rect 438 360 441 363 
rect 438 363 441 366 
rect 438 366 441 369 
rect 438 369 441 372 
rect 438 372 441 375 
rect 438 375 441 378 
rect 438 378 441 381 
rect 438 381 441 384 
rect 438 384 441 387 
rect 438 387 441 390 
rect 438 390 441 393 
rect 438 393 441 396 
rect 438 396 441 399 
rect 438 399 441 402 
rect 438 402 441 405 
rect 438 405 441 408 
rect 438 408 441 411 
rect 438 411 441 414 
rect 438 414 441 417 
rect 438 417 441 420 
rect 438 420 441 423 
rect 438 423 441 426 
rect 438 426 441 429 
rect 438 429 441 432 
rect 438 432 441 435 
rect 438 435 441 438 
rect 438 438 441 441 
rect 438 441 441 444 
rect 438 444 441 447 
rect 438 447 441 450 
rect 438 450 441 453 
rect 438 453 441 456 
rect 438 456 441 459 
rect 438 459 441 462 
rect 438 462 441 465 
rect 438 465 441 468 
rect 438 468 441 471 
rect 438 471 441 474 
rect 438 474 441 477 
rect 438 477 441 480 
rect 438 480 441 483 
rect 438 483 441 486 
rect 438 486 441 489 
rect 438 489 441 492 
rect 438 492 441 495 
rect 438 495 441 498 
rect 438 498 441 501 
rect 438 501 441 504 
rect 438 504 441 507 
rect 438 507 441 510 
rect 441 0 444 3 
rect 441 3 444 6 
rect 441 6 444 9 
rect 441 9 444 12 
rect 441 12 444 15 
rect 441 15 444 18 
rect 441 18 444 21 
rect 441 21 444 24 
rect 441 24 444 27 
rect 441 27 444 30 
rect 441 30 444 33 
rect 441 33 444 36 
rect 441 36 444 39 
rect 441 39 444 42 
rect 441 42 444 45 
rect 441 45 444 48 
rect 441 48 444 51 
rect 441 51 444 54 
rect 441 54 444 57 
rect 441 57 444 60 
rect 441 60 444 63 
rect 441 63 444 66 
rect 441 66 444 69 
rect 441 69 444 72 
rect 441 72 444 75 
rect 441 75 444 78 
rect 441 78 444 81 
rect 441 81 444 84 
rect 441 84 444 87 
rect 441 87 444 90 
rect 441 90 444 93 
rect 441 93 444 96 
rect 441 96 444 99 
rect 441 99 444 102 
rect 441 102 444 105 
rect 441 105 444 108 
rect 441 108 444 111 
rect 441 111 444 114 
rect 441 114 444 117 
rect 441 117 444 120 
rect 441 120 444 123 
rect 441 123 444 126 
rect 441 126 444 129 
rect 441 129 444 132 
rect 441 132 444 135 
rect 441 135 444 138 
rect 441 138 444 141 
rect 441 141 444 144 
rect 441 144 444 147 
rect 441 147 444 150 
rect 441 150 444 153 
rect 441 153 444 156 
rect 441 156 444 159 
rect 441 159 444 162 
rect 441 162 444 165 
rect 441 165 444 168 
rect 441 168 444 171 
rect 441 171 444 174 
rect 441 174 444 177 
rect 441 177 444 180 
rect 441 180 444 183 
rect 441 183 444 186 
rect 441 186 444 189 
rect 441 189 444 192 
rect 441 192 444 195 
rect 441 195 444 198 
rect 441 198 444 201 
rect 441 201 444 204 
rect 441 204 444 207 
rect 441 207 444 210 
rect 441 210 444 213 
rect 441 213 444 216 
rect 441 216 444 219 
rect 441 219 444 222 
rect 441 222 444 225 
rect 441 225 444 228 
rect 441 228 444 231 
rect 441 231 444 234 
rect 441 234 444 237 
rect 441 237 444 240 
rect 441 240 444 243 
rect 441 243 444 246 
rect 441 246 444 249 
rect 441 249 444 252 
rect 441 252 444 255 
rect 441 255 444 258 
rect 441 258 444 261 
rect 441 261 444 264 
rect 441 264 444 267 
rect 441 267 444 270 
rect 441 270 444 273 
rect 441 273 444 276 
rect 441 276 444 279 
rect 441 279 444 282 
rect 441 282 444 285 
rect 441 285 444 288 
rect 441 288 444 291 
rect 441 291 444 294 
rect 441 294 444 297 
rect 441 297 444 300 
rect 441 300 444 303 
rect 441 303 444 306 
rect 441 306 444 309 
rect 441 309 444 312 
rect 441 312 444 315 
rect 441 315 444 318 
rect 441 318 444 321 
rect 441 321 444 324 
rect 441 324 444 327 
rect 441 327 444 330 
rect 441 330 444 333 
rect 441 333 444 336 
rect 441 336 444 339 
rect 441 339 444 342 
rect 441 342 444 345 
rect 441 345 444 348 
rect 441 348 444 351 
rect 441 351 444 354 
rect 441 354 444 357 
rect 441 357 444 360 
rect 441 360 444 363 
rect 441 363 444 366 
rect 441 366 444 369 
rect 441 369 444 372 
rect 441 372 444 375 
rect 441 375 444 378 
rect 441 378 444 381 
rect 441 381 444 384 
rect 441 384 444 387 
rect 441 387 444 390 
rect 441 390 444 393 
rect 441 393 444 396 
rect 441 396 444 399 
rect 441 399 444 402 
rect 441 402 444 405 
rect 441 405 444 408 
rect 441 408 444 411 
rect 441 411 444 414 
rect 441 414 444 417 
rect 441 417 444 420 
rect 441 420 444 423 
rect 441 423 444 426 
rect 441 426 444 429 
rect 441 429 444 432 
rect 441 432 444 435 
rect 441 435 444 438 
rect 441 438 444 441 
rect 441 441 444 444 
rect 441 444 444 447 
rect 441 447 444 450 
rect 441 450 444 453 
rect 441 453 444 456 
rect 441 456 444 459 
rect 441 459 444 462 
rect 441 462 444 465 
rect 441 465 444 468 
rect 441 468 444 471 
rect 441 471 444 474 
rect 441 474 444 477 
rect 441 477 444 480 
rect 441 480 444 483 
rect 441 483 444 486 
rect 441 486 444 489 
rect 441 489 444 492 
rect 441 492 444 495 
rect 441 495 444 498 
rect 441 498 444 501 
rect 441 501 444 504 
rect 441 504 444 507 
rect 441 507 444 510 
rect 444 0 447 3 
rect 444 3 447 6 
rect 444 6 447 9 
rect 444 9 447 12 
rect 444 12 447 15 
rect 444 15 447 18 
rect 444 18 447 21 
rect 444 21 447 24 
rect 444 24 447 27 
rect 444 27 447 30 
rect 444 30 447 33 
rect 444 33 447 36 
rect 444 36 447 39 
rect 444 39 447 42 
rect 444 42 447 45 
rect 444 45 447 48 
rect 444 48 447 51 
rect 444 51 447 54 
rect 444 54 447 57 
rect 444 57 447 60 
rect 444 60 447 63 
rect 444 63 447 66 
rect 444 66 447 69 
rect 444 69 447 72 
rect 444 72 447 75 
rect 444 75 447 78 
rect 444 78 447 81 
rect 444 81 447 84 
rect 444 84 447 87 
rect 444 87 447 90 
rect 444 90 447 93 
rect 444 93 447 96 
rect 444 96 447 99 
rect 444 99 447 102 
rect 444 102 447 105 
rect 444 105 447 108 
rect 444 108 447 111 
rect 444 111 447 114 
rect 444 114 447 117 
rect 444 117 447 120 
rect 444 120 447 123 
rect 444 123 447 126 
rect 444 126 447 129 
rect 444 129 447 132 
rect 444 132 447 135 
rect 444 135 447 138 
rect 444 138 447 141 
rect 444 141 447 144 
rect 444 144 447 147 
rect 444 147 447 150 
rect 444 150 447 153 
rect 444 153 447 156 
rect 444 156 447 159 
rect 444 159 447 162 
rect 444 162 447 165 
rect 444 165 447 168 
rect 444 168 447 171 
rect 444 171 447 174 
rect 444 174 447 177 
rect 444 177 447 180 
rect 444 180 447 183 
rect 444 183 447 186 
rect 444 186 447 189 
rect 444 189 447 192 
rect 444 192 447 195 
rect 444 195 447 198 
rect 444 198 447 201 
rect 444 201 447 204 
rect 444 204 447 207 
rect 444 207 447 210 
rect 444 210 447 213 
rect 444 213 447 216 
rect 444 216 447 219 
rect 444 219 447 222 
rect 444 222 447 225 
rect 444 225 447 228 
rect 444 228 447 231 
rect 444 231 447 234 
rect 444 234 447 237 
rect 444 237 447 240 
rect 444 240 447 243 
rect 444 243 447 246 
rect 444 246 447 249 
rect 444 249 447 252 
rect 444 252 447 255 
rect 444 255 447 258 
rect 444 258 447 261 
rect 444 261 447 264 
rect 444 264 447 267 
rect 444 267 447 270 
rect 444 270 447 273 
rect 444 273 447 276 
rect 444 276 447 279 
rect 444 279 447 282 
rect 444 282 447 285 
rect 444 285 447 288 
rect 444 288 447 291 
rect 444 291 447 294 
rect 444 294 447 297 
rect 444 297 447 300 
rect 444 300 447 303 
rect 444 303 447 306 
rect 444 306 447 309 
rect 444 309 447 312 
rect 444 312 447 315 
rect 444 315 447 318 
rect 444 318 447 321 
rect 444 321 447 324 
rect 444 324 447 327 
rect 444 327 447 330 
rect 444 330 447 333 
rect 444 333 447 336 
rect 444 336 447 339 
rect 444 339 447 342 
rect 444 342 447 345 
rect 444 345 447 348 
rect 444 348 447 351 
rect 444 351 447 354 
rect 444 354 447 357 
rect 444 357 447 360 
rect 444 360 447 363 
rect 444 363 447 366 
rect 444 366 447 369 
rect 444 369 447 372 
rect 444 372 447 375 
rect 444 375 447 378 
rect 444 378 447 381 
rect 444 381 447 384 
rect 444 384 447 387 
rect 444 387 447 390 
rect 444 390 447 393 
rect 444 393 447 396 
rect 444 396 447 399 
rect 444 399 447 402 
rect 444 402 447 405 
rect 444 405 447 408 
rect 444 408 447 411 
rect 444 411 447 414 
rect 444 414 447 417 
rect 444 417 447 420 
rect 444 420 447 423 
rect 444 423 447 426 
rect 444 426 447 429 
rect 444 429 447 432 
rect 444 432 447 435 
rect 444 435 447 438 
rect 444 438 447 441 
rect 444 441 447 444 
rect 444 444 447 447 
rect 444 447 447 450 
rect 444 450 447 453 
rect 444 453 447 456 
rect 444 456 447 459 
rect 444 459 447 462 
rect 444 462 447 465 
rect 444 465 447 468 
rect 444 468 447 471 
rect 444 471 447 474 
rect 444 474 447 477 
rect 444 477 447 480 
rect 444 480 447 483 
rect 444 483 447 486 
rect 444 486 447 489 
rect 444 489 447 492 
rect 444 492 447 495 
rect 444 495 447 498 
rect 444 498 447 501 
rect 444 501 447 504 
rect 444 504 447 507 
rect 444 507 447 510 
rect 447 0 450 3 
rect 447 3 450 6 
rect 447 6 450 9 
rect 447 9 450 12 
rect 447 12 450 15 
rect 447 15 450 18 
rect 447 18 450 21 
rect 447 21 450 24 
rect 447 24 450 27 
rect 447 27 450 30 
rect 447 30 450 33 
rect 447 33 450 36 
rect 447 36 450 39 
rect 447 39 450 42 
rect 447 42 450 45 
rect 447 45 450 48 
rect 447 48 450 51 
rect 447 51 450 54 
rect 447 54 450 57 
rect 447 57 450 60 
rect 447 60 450 63 
rect 447 63 450 66 
rect 447 66 450 69 
rect 447 69 450 72 
rect 447 72 450 75 
rect 447 75 450 78 
rect 447 78 450 81 
rect 447 81 450 84 
rect 447 84 450 87 
rect 447 87 450 90 
rect 447 90 450 93 
rect 447 93 450 96 
rect 447 96 450 99 
rect 447 99 450 102 
rect 447 102 450 105 
rect 447 105 450 108 
rect 447 108 450 111 
rect 447 111 450 114 
rect 447 114 450 117 
rect 447 117 450 120 
rect 447 120 450 123 
rect 447 123 450 126 
rect 447 126 450 129 
rect 447 129 450 132 
rect 447 132 450 135 
rect 447 135 450 138 
rect 447 138 450 141 
rect 447 141 450 144 
rect 447 144 450 147 
rect 447 147 450 150 
rect 447 150 450 153 
rect 447 153 450 156 
rect 447 156 450 159 
rect 447 159 450 162 
rect 447 162 450 165 
rect 447 165 450 168 
rect 447 168 450 171 
rect 447 171 450 174 
rect 447 174 450 177 
rect 447 177 450 180 
rect 447 180 450 183 
rect 447 183 450 186 
rect 447 186 450 189 
rect 447 189 450 192 
rect 447 192 450 195 
rect 447 195 450 198 
rect 447 198 450 201 
rect 447 201 450 204 
rect 447 204 450 207 
rect 447 207 450 210 
rect 447 210 450 213 
rect 447 213 450 216 
rect 447 216 450 219 
rect 447 219 450 222 
rect 447 222 450 225 
rect 447 225 450 228 
rect 447 228 450 231 
rect 447 231 450 234 
rect 447 234 450 237 
rect 447 237 450 240 
rect 447 240 450 243 
rect 447 243 450 246 
rect 447 246 450 249 
rect 447 249 450 252 
rect 447 252 450 255 
rect 447 255 450 258 
rect 447 258 450 261 
rect 447 261 450 264 
rect 447 264 450 267 
rect 447 267 450 270 
rect 447 270 450 273 
rect 447 273 450 276 
rect 447 276 450 279 
rect 447 279 450 282 
rect 447 282 450 285 
rect 447 285 450 288 
rect 447 288 450 291 
rect 447 291 450 294 
rect 447 294 450 297 
rect 447 297 450 300 
rect 447 300 450 303 
rect 447 303 450 306 
rect 447 306 450 309 
rect 447 309 450 312 
rect 447 312 450 315 
rect 447 315 450 318 
rect 447 318 450 321 
rect 447 321 450 324 
rect 447 324 450 327 
rect 447 327 450 330 
rect 447 330 450 333 
rect 447 333 450 336 
rect 447 336 450 339 
rect 447 339 450 342 
rect 447 342 450 345 
rect 447 345 450 348 
rect 447 348 450 351 
rect 447 351 450 354 
rect 447 354 450 357 
rect 447 357 450 360 
rect 447 360 450 363 
rect 447 363 450 366 
rect 447 366 450 369 
rect 447 369 450 372 
rect 447 372 450 375 
rect 447 375 450 378 
rect 447 378 450 381 
rect 447 381 450 384 
rect 447 384 450 387 
rect 447 387 450 390 
rect 447 390 450 393 
rect 447 393 450 396 
rect 447 396 450 399 
rect 447 399 450 402 
rect 447 402 450 405 
rect 447 405 450 408 
rect 447 408 450 411 
rect 447 411 450 414 
rect 447 414 450 417 
rect 447 417 450 420 
rect 447 420 450 423 
rect 447 423 450 426 
rect 447 426 450 429 
rect 447 429 450 432 
rect 447 432 450 435 
rect 447 435 450 438 
rect 447 438 450 441 
rect 447 441 450 444 
rect 447 444 450 447 
rect 447 447 450 450 
rect 447 450 450 453 
rect 447 453 450 456 
rect 447 456 450 459 
rect 447 459 450 462 
rect 447 462 450 465 
rect 447 465 450 468 
rect 447 468 450 471 
rect 447 471 450 474 
rect 447 474 450 477 
rect 447 477 450 480 
rect 447 480 450 483 
rect 447 483 450 486 
rect 447 486 450 489 
rect 447 489 450 492 
rect 447 492 450 495 
rect 447 495 450 498 
rect 447 498 450 501 
rect 447 501 450 504 
rect 447 504 450 507 
rect 447 507 450 510 
rect 450 0 453 3 
rect 450 3 453 6 
rect 450 6 453 9 
rect 450 9 453 12 
rect 450 12 453 15 
rect 450 15 453 18 
rect 450 18 453 21 
rect 450 21 453 24 
rect 450 24 453 27 
rect 450 27 453 30 
rect 450 30 453 33 
rect 450 33 453 36 
rect 450 36 453 39 
rect 450 39 453 42 
rect 450 42 453 45 
rect 450 45 453 48 
rect 450 48 453 51 
rect 450 51 453 54 
rect 450 54 453 57 
rect 450 57 453 60 
rect 450 60 453 63 
rect 450 63 453 66 
rect 450 66 453 69 
rect 450 69 453 72 
rect 450 72 453 75 
rect 450 75 453 78 
rect 450 78 453 81 
rect 450 81 453 84 
rect 450 84 453 87 
rect 450 87 453 90 
rect 450 90 453 93 
rect 450 93 453 96 
rect 450 96 453 99 
rect 450 99 453 102 
rect 450 102 453 105 
rect 450 105 453 108 
rect 450 108 453 111 
rect 450 111 453 114 
rect 450 114 453 117 
rect 450 117 453 120 
rect 450 120 453 123 
rect 450 123 453 126 
rect 450 126 453 129 
rect 450 129 453 132 
rect 450 132 453 135 
rect 450 135 453 138 
rect 450 138 453 141 
rect 450 141 453 144 
rect 450 144 453 147 
rect 450 147 453 150 
rect 450 150 453 153 
rect 450 153 453 156 
rect 450 156 453 159 
rect 450 159 453 162 
rect 450 162 453 165 
rect 450 165 453 168 
rect 450 168 453 171 
rect 450 171 453 174 
rect 450 174 453 177 
rect 450 177 453 180 
rect 450 180 453 183 
rect 450 183 453 186 
rect 450 186 453 189 
rect 450 189 453 192 
rect 450 192 453 195 
rect 450 195 453 198 
rect 450 198 453 201 
rect 450 201 453 204 
rect 450 204 453 207 
rect 450 207 453 210 
rect 450 210 453 213 
rect 450 213 453 216 
rect 450 216 453 219 
rect 450 219 453 222 
rect 450 222 453 225 
rect 450 225 453 228 
rect 450 228 453 231 
rect 450 231 453 234 
rect 450 234 453 237 
rect 450 237 453 240 
rect 450 240 453 243 
rect 450 243 453 246 
rect 450 246 453 249 
rect 450 249 453 252 
rect 450 252 453 255 
rect 450 255 453 258 
rect 450 258 453 261 
rect 450 261 453 264 
rect 450 264 453 267 
rect 450 267 453 270 
rect 450 270 453 273 
rect 450 273 453 276 
rect 450 276 453 279 
rect 450 279 453 282 
rect 450 282 453 285 
rect 450 285 453 288 
rect 450 288 453 291 
rect 450 291 453 294 
rect 450 294 453 297 
rect 450 297 453 300 
rect 450 300 453 303 
rect 450 303 453 306 
rect 450 306 453 309 
rect 450 309 453 312 
rect 450 312 453 315 
rect 450 315 453 318 
rect 450 318 453 321 
rect 450 321 453 324 
rect 450 324 453 327 
rect 450 327 453 330 
rect 450 330 453 333 
rect 450 333 453 336 
rect 450 336 453 339 
rect 450 339 453 342 
rect 450 342 453 345 
rect 450 345 453 348 
rect 450 348 453 351 
rect 450 351 453 354 
rect 450 354 453 357 
rect 450 357 453 360 
rect 450 360 453 363 
rect 450 363 453 366 
rect 450 366 453 369 
rect 450 369 453 372 
rect 450 372 453 375 
rect 450 375 453 378 
rect 450 378 453 381 
rect 450 381 453 384 
rect 450 384 453 387 
rect 450 387 453 390 
rect 450 390 453 393 
rect 450 393 453 396 
rect 450 396 453 399 
rect 450 399 453 402 
rect 450 402 453 405 
rect 450 405 453 408 
rect 450 408 453 411 
rect 450 411 453 414 
rect 450 414 453 417 
rect 450 417 453 420 
rect 450 420 453 423 
rect 450 423 453 426 
rect 450 426 453 429 
rect 450 429 453 432 
rect 450 432 453 435 
rect 450 435 453 438 
rect 450 438 453 441 
rect 450 441 453 444 
rect 450 444 453 447 
rect 450 447 453 450 
rect 450 450 453 453 
rect 450 453 453 456 
rect 450 456 453 459 
rect 450 459 453 462 
rect 450 462 453 465 
rect 450 465 453 468 
rect 450 468 453 471 
rect 450 471 453 474 
rect 450 474 453 477 
rect 450 477 453 480 
rect 450 480 453 483 
rect 450 483 453 486 
rect 450 486 453 489 
rect 450 489 453 492 
rect 450 492 453 495 
rect 450 495 453 498 
rect 450 498 453 501 
rect 450 501 453 504 
rect 450 504 453 507 
rect 450 507 453 510 
rect 453 0 456 3 
rect 453 3 456 6 
rect 453 6 456 9 
rect 453 9 456 12 
rect 453 12 456 15 
rect 453 15 456 18 
rect 453 18 456 21 
rect 453 21 456 24 
rect 453 24 456 27 
rect 453 27 456 30 
rect 453 30 456 33 
rect 453 33 456 36 
rect 453 36 456 39 
rect 453 39 456 42 
rect 453 42 456 45 
rect 453 45 456 48 
rect 453 48 456 51 
rect 453 51 456 54 
rect 453 54 456 57 
rect 453 57 456 60 
rect 453 60 456 63 
rect 453 63 456 66 
rect 453 66 456 69 
rect 453 69 456 72 
rect 453 72 456 75 
rect 453 75 456 78 
rect 453 78 456 81 
rect 453 81 456 84 
rect 453 84 456 87 
rect 453 87 456 90 
rect 453 90 456 93 
rect 453 93 456 96 
rect 453 96 456 99 
rect 453 99 456 102 
rect 453 102 456 105 
rect 453 105 456 108 
rect 453 108 456 111 
rect 453 111 456 114 
rect 453 114 456 117 
rect 453 117 456 120 
rect 453 120 456 123 
rect 453 123 456 126 
rect 453 126 456 129 
rect 453 129 456 132 
rect 453 132 456 135 
rect 453 135 456 138 
rect 453 138 456 141 
rect 453 141 456 144 
rect 453 144 456 147 
rect 453 147 456 150 
rect 453 150 456 153 
rect 453 153 456 156 
rect 453 156 456 159 
rect 453 159 456 162 
rect 453 162 456 165 
rect 453 165 456 168 
rect 453 168 456 171 
rect 453 171 456 174 
rect 453 174 456 177 
rect 453 177 456 180 
rect 453 180 456 183 
rect 453 183 456 186 
rect 453 186 456 189 
rect 453 189 456 192 
rect 453 192 456 195 
rect 453 195 456 198 
rect 453 198 456 201 
rect 453 201 456 204 
rect 453 204 456 207 
rect 453 207 456 210 
rect 453 210 456 213 
rect 453 213 456 216 
rect 453 216 456 219 
rect 453 219 456 222 
rect 453 222 456 225 
rect 453 225 456 228 
rect 453 228 456 231 
rect 453 231 456 234 
rect 453 234 456 237 
rect 453 237 456 240 
rect 453 240 456 243 
rect 453 243 456 246 
rect 453 246 456 249 
rect 453 249 456 252 
rect 453 252 456 255 
rect 453 255 456 258 
rect 453 258 456 261 
rect 453 261 456 264 
rect 453 264 456 267 
rect 453 267 456 270 
rect 453 270 456 273 
rect 453 273 456 276 
rect 453 276 456 279 
rect 453 279 456 282 
rect 453 282 456 285 
rect 453 285 456 288 
rect 453 288 456 291 
rect 453 291 456 294 
rect 453 294 456 297 
rect 453 297 456 300 
rect 453 300 456 303 
rect 453 303 456 306 
rect 453 306 456 309 
rect 453 309 456 312 
rect 453 312 456 315 
rect 453 315 456 318 
rect 453 318 456 321 
rect 453 321 456 324 
rect 453 324 456 327 
rect 453 327 456 330 
rect 453 330 456 333 
rect 453 333 456 336 
rect 453 336 456 339 
rect 453 339 456 342 
rect 453 342 456 345 
rect 453 345 456 348 
rect 453 348 456 351 
rect 453 351 456 354 
rect 453 354 456 357 
rect 453 357 456 360 
rect 453 360 456 363 
rect 453 363 456 366 
rect 453 366 456 369 
rect 453 369 456 372 
rect 453 372 456 375 
rect 453 375 456 378 
rect 453 378 456 381 
rect 453 381 456 384 
rect 453 384 456 387 
rect 453 387 456 390 
rect 453 390 456 393 
rect 453 393 456 396 
rect 453 396 456 399 
rect 453 399 456 402 
rect 453 402 456 405 
rect 453 405 456 408 
rect 453 408 456 411 
rect 453 411 456 414 
rect 453 414 456 417 
rect 453 417 456 420 
rect 453 420 456 423 
rect 453 423 456 426 
rect 453 426 456 429 
rect 453 429 456 432 
rect 453 432 456 435 
rect 453 435 456 438 
rect 453 438 456 441 
rect 453 441 456 444 
rect 453 444 456 447 
rect 453 447 456 450 
rect 453 450 456 453 
rect 453 453 456 456 
rect 453 456 456 459 
rect 453 459 456 462 
rect 453 462 456 465 
rect 453 465 456 468 
rect 453 468 456 471 
rect 453 471 456 474 
rect 453 474 456 477 
rect 453 477 456 480 
rect 453 480 456 483 
rect 453 483 456 486 
rect 453 486 456 489 
rect 453 489 456 492 
rect 453 492 456 495 
rect 453 495 456 498 
rect 453 498 456 501 
rect 453 501 456 504 
rect 453 504 456 507 
rect 453 507 456 510 
rect 456 0 459 3 
rect 456 3 459 6 
rect 456 6 459 9 
rect 456 9 459 12 
rect 456 12 459 15 
rect 456 15 459 18 
rect 456 18 459 21 
rect 456 21 459 24 
rect 456 24 459 27 
rect 456 27 459 30 
rect 456 30 459 33 
rect 456 33 459 36 
rect 456 36 459 39 
rect 456 39 459 42 
rect 456 42 459 45 
rect 456 45 459 48 
rect 456 48 459 51 
rect 456 51 459 54 
rect 456 54 459 57 
rect 456 57 459 60 
rect 456 60 459 63 
rect 456 63 459 66 
rect 456 66 459 69 
rect 456 69 459 72 
rect 456 72 459 75 
rect 456 75 459 78 
rect 456 78 459 81 
rect 456 81 459 84 
rect 456 84 459 87 
rect 456 87 459 90 
rect 456 90 459 93 
rect 456 93 459 96 
rect 456 96 459 99 
rect 456 99 459 102 
rect 456 102 459 105 
rect 456 105 459 108 
rect 456 108 459 111 
rect 456 111 459 114 
rect 456 114 459 117 
rect 456 117 459 120 
rect 456 120 459 123 
rect 456 123 459 126 
rect 456 126 459 129 
rect 456 129 459 132 
rect 456 132 459 135 
rect 456 135 459 138 
rect 456 138 459 141 
rect 456 141 459 144 
rect 456 144 459 147 
rect 456 147 459 150 
rect 456 150 459 153 
rect 456 153 459 156 
rect 456 156 459 159 
rect 456 159 459 162 
rect 456 162 459 165 
rect 456 165 459 168 
rect 456 168 459 171 
rect 456 171 459 174 
rect 456 174 459 177 
rect 456 177 459 180 
rect 456 180 459 183 
rect 456 183 459 186 
rect 456 186 459 189 
rect 456 189 459 192 
rect 456 192 459 195 
rect 456 195 459 198 
rect 456 198 459 201 
rect 456 201 459 204 
rect 456 204 459 207 
rect 456 207 459 210 
rect 456 210 459 213 
rect 456 213 459 216 
rect 456 216 459 219 
rect 456 219 459 222 
rect 456 222 459 225 
rect 456 225 459 228 
rect 456 228 459 231 
rect 456 231 459 234 
rect 456 234 459 237 
rect 456 237 459 240 
rect 456 240 459 243 
rect 456 243 459 246 
rect 456 246 459 249 
rect 456 249 459 252 
rect 456 252 459 255 
rect 456 255 459 258 
rect 456 258 459 261 
rect 456 261 459 264 
rect 456 264 459 267 
rect 456 267 459 270 
rect 456 270 459 273 
rect 456 273 459 276 
rect 456 276 459 279 
rect 456 279 459 282 
rect 456 282 459 285 
rect 456 285 459 288 
rect 456 288 459 291 
rect 456 291 459 294 
rect 456 294 459 297 
rect 456 297 459 300 
rect 456 300 459 303 
rect 456 303 459 306 
rect 456 306 459 309 
rect 456 309 459 312 
rect 456 312 459 315 
rect 456 315 459 318 
rect 456 318 459 321 
rect 456 321 459 324 
rect 456 324 459 327 
rect 456 327 459 330 
rect 456 330 459 333 
rect 456 333 459 336 
rect 456 336 459 339 
rect 456 339 459 342 
rect 456 342 459 345 
rect 456 345 459 348 
rect 456 348 459 351 
rect 456 351 459 354 
rect 456 354 459 357 
rect 456 357 459 360 
rect 456 360 459 363 
rect 456 363 459 366 
rect 456 366 459 369 
rect 456 369 459 372 
rect 456 372 459 375 
rect 456 375 459 378 
rect 456 378 459 381 
rect 456 381 459 384 
rect 456 384 459 387 
rect 456 387 459 390 
rect 456 390 459 393 
rect 456 393 459 396 
rect 456 396 459 399 
rect 456 399 459 402 
rect 456 402 459 405 
rect 456 405 459 408 
rect 456 408 459 411 
rect 456 411 459 414 
rect 456 414 459 417 
rect 456 417 459 420 
rect 456 420 459 423 
rect 456 423 459 426 
rect 456 426 459 429 
rect 456 429 459 432 
rect 456 432 459 435 
rect 456 435 459 438 
rect 456 438 459 441 
rect 456 441 459 444 
rect 456 444 459 447 
rect 456 447 459 450 
rect 456 450 459 453 
rect 456 453 459 456 
rect 456 456 459 459 
rect 456 459 459 462 
rect 456 462 459 465 
rect 456 465 459 468 
rect 456 468 459 471 
rect 456 471 459 474 
rect 456 474 459 477 
rect 456 477 459 480 
rect 456 480 459 483 
rect 456 483 459 486 
rect 456 486 459 489 
rect 456 489 459 492 
rect 456 492 459 495 
rect 456 495 459 498 
rect 456 498 459 501 
rect 456 501 459 504 
rect 456 504 459 507 
rect 456 507 459 510 
rect 459 0 462 3 
rect 459 3 462 6 
rect 459 6 462 9 
rect 459 9 462 12 
rect 459 12 462 15 
rect 459 15 462 18 
rect 459 18 462 21 
rect 459 21 462 24 
rect 459 24 462 27 
rect 459 27 462 30 
rect 459 30 462 33 
rect 459 33 462 36 
rect 459 36 462 39 
rect 459 39 462 42 
rect 459 42 462 45 
rect 459 45 462 48 
rect 459 48 462 51 
rect 459 51 462 54 
rect 459 54 462 57 
rect 459 57 462 60 
rect 459 60 462 63 
rect 459 63 462 66 
rect 459 66 462 69 
rect 459 69 462 72 
rect 459 72 462 75 
rect 459 75 462 78 
rect 459 78 462 81 
rect 459 81 462 84 
rect 459 84 462 87 
rect 459 87 462 90 
rect 459 90 462 93 
rect 459 93 462 96 
rect 459 96 462 99 
rect 459 99 462 102 
rect 459 102 462 105 
rect 459 105 462 108 
rect 459 108 462 111 
rect 459 111 462 114 
rect 459 114 462 117 
rect 459 117 462 120 
rect 459 120 462 123 
rect 459 123 462 126 
rect 459 126 462 129 
rect 459 129 462 132 
rect 459 132 462 135 
rect 459 135 462 138 
rect 459 138 462 141 
rect 459 141 462 144 
rect 459 144 462 147 
rect 459 147 462 150 
rect 459 150 462 153 
rect 459 153 462 156 
rect 459 156 462 159 
rect 459 159 462 162 
rect 459 162 462 165 
rect 459 165 462 168 
rect 459 168 462 171 
rect 459 171 462 174 
rect 459 174 462 177 
rect 459 177 462 180 
rect 459 180 462 183 
rect 459 183 462 186 
rect 459 186 462 189 
rect 459 189 462 192 
rect 459 192 462 195 
rect 459 195 462 198 
rect 459 198 462 201 
rect 459 201 462 204 
rect 459 204 462 207 
rect 459 207 462 210 
rect 459 210 462 213 
rect 459 213 462 216 
rect 459 216 462 219 
rect 459 219 462 222 
rect 459 222 462 225 
rect 459 225 462 228 
rect 459 228 462 231 
rect 459 231 462 234 
rect 459 234 462 237 
rect 459 237 462 240 
rect 459 240 462 243 
rect 459 243 462 246 
rect 459 246 462 249 
rect 459 249 462 252 
rect 459 252 462 255 
rect 459 255 462 258 
rect 459 258 462 261 
rect 459 261 462 264 
rect 459 264 462 267 
rect 459 267 462 270 
rect 459 270 462 273 
rect 459 273 462 276 
rect 459 276 462 279 
rect 459 279 462 282 
rect 459 282 462 285 
rect 459 285 462 288 
rect 459 288 462 291 
rect 459 291 462 294 
rect 459 294 462 297 
rect 459 297 462 300 
rect 459 300 462 303 
rect 459 303 462 306 
rect 459 306 462 309 
rect 459 309 462 312 
rect 459 312 462 315 
rect 459 315 462 318 
rect 459 318 462 321 
rect 459 321 462 324 
rect 459 324 462 327 
rect 459 327 462 330 
rect 459 330 462 333 
rect 459 333 462 336 
rect 459 336 462 339 
rect 459 339 462 342 
rect 459 342 462 345 
rect 459 345 462 348 
rect 459 348 462 351 
rect 459 351 462 354 
rect 459 354 462 357 
rect 459 357 462 360 
rect 459 360 462 363 
rect 459 363 462 366 
rect 459 366 462 369 
rect 459 369 462 372 
rect 459 372 462 375 
rect 459 375 462 378 
rect 459 378 462 381 
rect 459 381 462 384 
rect 459 384 462 387 
rect 459 387 462 390 
rect 459 390 462 393 
rect 459 393 462 396 
rect 459 396 462 399 
rect 459 399 462 402 
rect 459 402 462 405 
rect 459 405 462 408 
rect 459 408 462 411 
rect 459 411 462 414 
rect 459 414 462 417 
rect 459 417 462 420 
rect 459 420 462 423 
rect 459 423 462 426 
rect 459 426 462 429 
rect 459 429 462 432 
rect 459 432 462 435 
rect 459 435 462 438 
rect 459 438 462 441 
rect 459 441 462 444 
rect 459 444 462 447 
rect 459 447 462 450 
rect 459 450 462 453 
rect 459 453 462 456 
rect 459 456 462 459 
rect 459 459 462 462 
rect 459 462 462 465 
rect 459 465 462 468 
rect 459 468 462 471 
rect 459 471 462 474 
rect 459 474 462 477 
rect 459 477 462 480 
rect 459 480 462 483 
rect 459 483 462 486 
rect 459 486 462 489 
rect 459 489 462 492 
rect 459 492 462 495 
rect 459 495 462 498 
rect 459 498 462 501 
rect 459 501 462 504 
rect 459 504 462 507 
rect 459 507 462 510 
rect 462 0 465 3 
rect 462 3 465 6 
rect 462 6 465 9 
rect 462 9 465 12 
rect 462 12 465 15 
rect 462 15 465 18 
rect 462 18 465 21 
rect 462 21 465 24 
rect 462 24 465 27 
rect 462 27 465 30 
rect 462 30 465 33 
rect 462 33 465 36 
rect 462 36 465 39 
rect 462 39 465 42 
rect 462 42 465 45 
rect 462 45 465 48 
rect 462 48 465 51 
rect 462 51 465 54 
rect 462 54 465 57 
rect 462 57 465 60 
rect 462 60 465 63 
rect 462 63 465 66 
rect 462 66 465 69 
rect 462 69 465 72 
rect 462 72 465 75 
rect 462 75 465 78 
rect 462 78 465 81 
rect 462 81 465 84 
rect 462 84 465 87 
rect 462 87 465 90 
rect 462 90 465 93 
rect 462 93 465 96 
rect 462 96 465 99 
rect 462 99 465 102 
rect 462 102 465 105 
rect 462 105 465 108 
rect 462 108 465 111 
rect 462 111 465 114 
rect 462 114 465 117 
rect 462 117 465 120 
rect 462 120 465 123 
rect 462 123 465 126 
rect 462 126 465 129 
rect 462 129 465 132 
rect 462 132 465 135 
rect 462 135 465 138 
rect 462 138 465 141 
rect 462 141 465 144 
rect 462 144 465 147 
rect 462 147 465 150 
rect 462 150 465 153 
rect 462 153 465 156 
rect 462 156 465 159 
rect 462 159 465 162 
rect 462 162 465 165 
rect 462 165 465 168 
rect 462 168 465 171 
rect 462 171 465 174 
rect 462 174 465 177 
rect 462 177 465 180 
rect 462 180 465 183 
rect 462 183 465 186 
rect 462 186 465 189 
rect 462 189 465 192 
rect 462 192 465 195 
rect 462 195 465 198 
rect 462 198 465 201 
rect 462 201 465 204 
rect 462 204 465 207 
rect 462 207 465 210 
rect 462 210 465 213 
rect 462 213 465 216 
rect 462 216 465 219 
rect 462 219 465 222 
rect 462 222 465 225 
rect 462 225 465 228 
rect 462 228 465 231 
rect 462 231 465 234 
rect 462 234 465 237 
rect 462 237 465 240 
rect 462 240 465 243 
rect 462 243 465 246 
rect 462 246 465 249 
rect 462 249 465 252 
rect 462 252 465 255 
rect 462 255 465 258 
rect 462 258 465 261 
rect 462 261 465 264 
rect 462 264 465 267 
rect 462 267 465 270 
rect 462 270 465 273 
rect 462 273 465 276 
rect 462 276 465 279 
rect 462 279 465 282 
rect 462 285 465 288 
rect 462 288 465 291 
rect 462 291 465 294 
rect 462 294 465 297 
rect 462 297 465 300 
rect 462 300 465 303 
rect 462 303 465 306 
rect 462 306 465 309 
rect 462 309 465 312 
rect 462 312 465 315 
rect 462 315 465 318 
rect 462 318 465 321 
rect 462 321 465 324 
rect 462 324 465 327 
rect 462 327 465 330 
rect 462 333 465 336 
rect 462 336 465 339 
rect 462 339 465 342 
rect 462 342 465 345 
rect 462 345 465 348 
rect 462 348 465 351 
rect 462 351 465 354 
rect 462 354 465 357 
rect 462 357 465 360 
rect 462 360 465 363 
rect 462 363 465 366 
rect 462 366 465 369 
rect 462 372 465 375 
rect 462 375 465 378 
rect 462 381 465 384 
rect 462 384 465 387 
rect 462 387 465 390 
rect 462 390 465 393 
rect 462 393 465 396 
rect 462 396 465 399 
rect 462 399 465 402 
rect 462 402 465 405 
rect 462 405 465 408 
rect 462 408 465 411 
rect 462 411 465 414 
rect 462 414 465 417 
rect 462 417 465 420 
rect 462 420 465 423 
rect 462 423 465 426 
rect 462 429 465 432 
rect 462 432 465 435 
rect 462 435 465 438 
rect 462 438 465 441 
rect 462 441 465 444 
rect 462 444 465 447 
rect 462 447 465 450 
rect 462 450 465 453 
rect 462 453 465 456 
rect 462 456 465 459 
rect 462 459 465 462 
rect 462 462 465 465 
rect 462 465 465 468 
rect 462 468 465 471 
rect 462 471 465 474 
rect 462 474 465 477 
rect 462 477 465 480 
rect 462 480 465 483 
rect 462 483 465 486 
rect 462 486 465 489 
rect 462 489 465 492 
rect 462 492 465 495 
rect 462 495 465 498 
rect 462 498 465 501 
rect 462 501 465 504 
rect 462 504 465 507 
rect 462 507 465 510 
rect 465 0 468 3 
rect 465 3 468 6 
rect 465 6 468 9 
rect 465 9 468 12 
rect 465 12 468 15 
rect 465 15 468 18 
rect 465 18 468 21 
rect 465 21 468 24 
rect 465 24 468 27 
rect 465 27 468 30 
rect 465 30 468 33 
rect 465 33 468 36 
rect 465 36 468 39 
rect 465 39 468 42 
rect 465 42 468 45 
rect 465 45 468 48 
rect 465 48 468 51 
rect 465 51 468 54 
rect 465 54 468 57 
rect 465 57 468 60 
rect 465 60 468 63 
rect 465 63 468 66 
rect 465 66 468 69 
rect 465 69 468 72 
rect 465 72 468 75 
rect 465 75 468 78 
rect 465 78 468 81 
rect 465 81 468 84 
rect 465 84 468 87 
rect 465 87 468 90 
rect 465 90 468 93 
rect 465 93 468 96 
rect 465 96 468 99 
rect 465 99 468 102 
rect 465 102 468 105 
rect 465 105 468 108 
rect 465 108 468 111 
rect 465 111 468 114 
rect 465 114 468 117 
rect 465 117 468 120 
rect 465 120 468 123 
rect 465 123 468 126 
rect 465 126 468 129 
rect 465 129 468 132 
rect 465 132 468 135 
rect 465 135 468 138 
rect 465 138 468 141 
rect 465 141 468 144 
rect 465 144 468 147 
rect 465 147 468 150 
rect 465 150 468 153 
rect 465 153 468 156 
rect 465 156 468 159 
rect 465 159 468 162 
rect 465 162 468 165 
rect 465 165 468 168 
rect 465 168 468 171 
rect 465 171 468 174 
rect 465 174 468 177 
rect 465 177 468 180 
rect 465 180 468 183 
rect 465 183 468 186 
rect 465 186 468 189 
rect 465 189 468 192 
rect 465 192 468 195 
rect 465 195 468 198 
rect 465 198 468 201 
rect 465 201 468 204 
rect 465 204 468 207 
rect 465 207 468 210 
rect 465 210 468 213 
rect 465 213 468 216 
rect 465 216 468 219 
rect 465 219 468 222 
rect 465 222 468 225 
rect 465 225 468 228 
rect 465 228 468 231 
rect 465 231 468 234 
rect 465 234 468 237 
rect 465 237 468 240 
rect 465 240 468 243 
rect 465 243 468 246 
rect 465 246 468 249 
rect 465 249 468 252 
rect 465 252 468 255 
rect 465 255 468 258 
rect 465 258 468 261 
rect 465 261 468 264 
rect 465 264 468 267 
rect 465 267 468 270 
rect 465 270 468 273 
rect 465 273 468 276 
rect 465 276 468 279 
rect 465 279 468 282 
rect 465 282 468 285 
rect 465 285 468 288 
rect 465 288 468 291 
rect 465 291 468 294 
rect 465 294 468 297 
rect 465 297 468 300 
rect 465 300 468 303 
rect 465 303 468 306 
rect 465 306 468 309 
rect 465 309 468 312 
rect 465 312 468 315 
rect 465 315 468 318 
rect 465 318 468 321 
rect 465 321 468 324 
rect 465 324 468 327 
rect 465 327 468 330 
rect 465 330 468 333 
rect 465 333 468 336 
rect 465 336 468 339 
rect 465 339 468 342 
rect 465 342 468 345 
rect 465 345 468 348 
rect 465 348 468 351 
rect 465 351 468 354 
rect 465 354 468 357 
rect 465 357 468 360 
rect 465 360 468 363 
rect 465 363 468 366 
rect 465 366 468 369 
rect 465 369 468 372 
rect 465 372 468 375 
rect 465 375 468 378 
rect 465 378 468 381 
rect 465 381 468 384 
rect 465 384 468 387 
rect 465 387 468 390 
rect 465 390 468 393 
rect 465 393 468 396 
rect 465 396 468 399 
rect 465 399 468 402 
rect 465 402 468 405 
rect 465 405 468 408 
rect 465 408 468 411 
rect 465 411 468 414 
rect 465 414 468 417 
rect 465 417 468 420 
rect 465 420 468 423 
rect 465 423 468 426 
rect 465 426 468 429 
rect 465 429 468 432 
rect 465 432 468 435 
rect 465 435 468 438 
rect 465 438 468 441 
rect 465 441 468 444 
rect 465 444 468 447 
rect 465 447 468 450 
rect 465 450 468 453 
rect 465 453 468 456 
rect 465 456 468 459 
rect 465 459 468 462 
rect 465 462 468 465 
rect 465 465 468 468 
rect 465 468 468 471 
rect 465 471 468 474 
rect 465 474 468 477 
rect 465 477 468 480 
rect 465 480 468 483 
rect 465 483 468 486 
rect 465 486 468 489 
rect 465 489 468 492 
rect 465 492 468 495 
rect 465 495 468 498 
rect 465 498 468 501 
rect 465 501 468 504 
rect 465 504 468 507 
rect 465 507 468 510 
rect 468 0 471 3 
rect 468 3 471 6 
rect 468 6 471 9 
rect 468 9 471 12 
rect 468 12 471 15 
rect 468 15 471 18 
rect 468 18 471 21 
rect 468 21 471 24 
rect 468 24 471 27 
rect 468 27 471 30 
rect 468 30 471 33 
rect 468 33 471 36 
rect 468 36 471 39 
rect 468 39 471 42 
rect 468 42 471 45 
rect 468 45 471 48 
rect 468 48 471 51 
rect 468 51 471 54 
rect 468 54 471 57 
rect 468 57 471 60 
rect 468 60 471 63 
rect 468 63 471 66 
rect 468 66 471 69 
rect 468 69 471 72 
rect 468 72 471 75 
rect 468 75 471 78 
rect 468 78 471 81 
rect 468 81 471 84 
rect 468 84 471 87 
rect 468 87 471 90 
rect 468 90 471 93 
rect 468 93 471 96 
rect 468 96 471 99 
rect 468 99 471 102 
rect 468 102 471 105 
rect 468 105 471 108 
rect 468 108 471 111 
rect 468 111 471 114 
rect 468 114 471 117 
rect 468 117 471 120 
rect 468 120 471 123 
rect 468 123 471 126 
rect 468 126 471 129 
rect 468 129 471 132 
rect 468 132 471 135 
rect 468 135 471 138 
rect 468 138 471 141 
rect 468 141 471 144 
rect 468 144 471 147 
rect 468 147 471 150 
rect 468 150 471 153 
rect 468 153 471 156 
rect 468 156 471 159 
rect 468 159 471 162 
rect 468 162 471 165 
rect 468 165 471 168 
rect 468 168 471 171 
rect 468 171 471 174 
rect 468 174 471 177 
rect 468 177 471 180 
rect 468 180 471 183 
rect 468 183 471 186 
rect 468 186 471 189 
rect 468 189 471 192 
rect 468 192 471 195 
rect 468 195 471 198 
rect 468 198 471 201 
rect 468 201 471 204 
rect 468 204 471 207 
rect 468 207 471 210 
rect 468 210 471 213 
rect 468 213 471 216 
rect 468 216 471 219 
rect 468 219 471 222 
rect 468 222 471 225 
rect 468 225 471 228 
rect 468 228 471 231 
rect 468 231 471 234 
rect 468 234 471 237 
rect 468 237 471 240 
rect 468 240 471 243 
rect 468 243 471 246 
rect 468 246 471 249 
rect 468 249 471 252 
rect 468 252 471 255 
rect 468 255 471 258 
rect 468 258 471 261 
rect 468 261 471 264 
rect 468 264 471 267 
rect 468 267 471 270 
rect 468 270 471 273 
rect 468 273 471 276 
rect 468 276 471 279 
rect 468 279 471 282 
rect 468 282 471 285 
rect 468 285 471 288 
rect 468 288 471 291 
rect 468 291 471 294 
rect 468 294 471 297 
rect 468 297 471 300 
rect 468 300 471 303 
rect 468 303 471 306 
rect 468 306 471 309 
rect 468 309 471 312 
rect 468 312 471 315 
rect 468 315 471 318 
rect 468 318 471 321 
rect 468 321 471 324 
rect 468 324 471 327 
rect 468 327 471 330 
rect 468 330 471 333 
rect 468 333 471 336 
rect 468 336 471 339 
rect 468 339 471 342 
rect 468 342 471 345 
rect 468 345 471 348 
rect 468 348 471 351 
rect 468 351 471 354 
rect 468 354 471 357 
rect 468 357 471 360 
rect 468 360 471 363 
rect 468 363 471 366 
rect 468 366 471 369 
rect 468 369 471 372 
rect 468 372 471 375 
rect 468 375 471 378 
rect 468 378 471 381 
rect 468 381 471 384 
rect 468 384 471 387 
rect 468 387 471 390 
rect 468 390 471 393 
rect 468 393 471 396 
rect 468 396 471 399 
rect 468 399 471 402 
rect 468 402 471 405 
rect 468 405 471 408 
rect 468 408 471 411 
rect 468 411 471 414 
rect 468 414 471 417 
rect 468 417 471 420 
rect 468 420 471 423 
rect 468 423 471 426 
rect 468 426 471 429 
rect 468 429 471 432 
rect 468 432 471 435 
rect 468 435 471 438 
rect 468 438 471 441 
rect 468 441 471 444 
rect 468 444 471 447 
rect 468 447 471 450 
rect 468 450 471 453 
rect 468 453 471 456 
rect 468 456 471 459 
rect 468 459 471 462 
rect 468 462 471 465 
rect 468 465 471 468 
rect 468 468 471 471 
rect 468 471 471 474 
rect 468 474 471 477 
rect 468 477 471 480 
rect 468 480 471 483 
rect 468 483 471 486 
rect 468 486 471 489 
rect 468 489 471 492 
rect 468 492 471 495 
rect 468 495 471 498 
rect 468 498 471 501 
rect 468 501 471 504 
rect 468 504 471 507 
rect 468 507 471 510 
rect 471 0 474 3 
rect 471 3 474 6 
rect 471 6 474 9 
rect 471 9 474 12 
rect 471 12 474 15 
rect 471 15 474 18 
rect 471 18 474 21 
rect 471 21 474 24 
rect 471 24 474 27 
rect 471 27 474 30 
rect 471 30 474 33 
rect 471 33 474 36 
rect 471 36 474 39 
rect 471 39 474 42 
rect 471 42 474 45 
rect 471 45 474 48 
rect 471 48 474 51 
rect 471 51 474 54 
rect 471 54 474 57 
rect 471 57 474 60 
rect 471 60 474 63 
rect 471 63 474 66 
rect 471 66 474 69 
rect 471 69 474 72 
rect 471 72 474 75 
rect 471 75 474 78 
rect 471 78 474 81 
rect 471 81 474 84 
rect 471 84 474 87 
rect 471 87 474 90 
rect 471 90 474 93 
rect 471 93 474 96 
rect 471 96 474 99 
rect 471 99 474 102 
rect 471 102 474 105 
rect 471 105 474 108 
rect 471 108 474 111 
rect 471 111 474 114 
rect 471 114 474 117 
rect 471 117 474 120 
rect 471 120 474 123 
rect 471 123 474 126 
rect 471 126 474 129 
rect 471 129 474 132 
rect 471 132 474 135 
rect 471 135 474 138 
rect 471 138 474 141 
rect 471 141 474 144 
rect 471 144 474 147 
rect 471 147 474 150 
rect 471 150 474 153 
rect 471 153 474 156 
rect 471 156 474 159 
rect 471 159 474 162 
rect 471 162 474 165 
rect 471 165 474 168 
rect 471 168 474 171 
rect 471 171 474 174 
rect 471 174 474 177 
rect 471 177 474 180 
rect 471 180 474 183 
rect 471 183 474 186 
rect 471 186 474 189 
rect 471 189 474 192 
rect 471 192 474 195 
rect 471 195 474 198 
rect 471 198 474 201 
rect 471 201 474 204 
rect 471 204 474 207 
rect 471 207 474 210 
rect 471 210 474 213 
rect 471 213 474 216 
rect 471 216 474 219 
rect 471 219 474 222 
rect 471 222 474 225 
rect 471 225 474 228 
rect 471 228 474 231 
rect 471 231 474 234 
rect 471 234 474 237 
rect 471 237 474 240 
rect 471 240 474 243 
rect 471 243 474 246 
rect 471 246 474 249 
rect 471 249 474 252 
rect 471 252 474 255 
rect 471 255 474 258 
rect 471 258 474 261 
rect 471 261 474 264 
rect 471 264 474 267 
rect 471 267 474 270 
rect 471 270 474 273 
rect 471 273 474 276 
rect 471 276 474 279 
rect 471 279 474 282 
rect 471 282 474 285 
rect 471 285 474 288 
rect 471 288 474 291 
rect 471 291 474 294 
rect 471 294 474 297 
rect 471 297 474 300 
rect 471 300 474 303 
rect 471 303 474 306 
rect 471 306 474 309 
rect 471 309 474 312 
rect 471 312 474 315 
rect 471 315 474 318 
rect 471 318 474 321 
rect 471 321 474 324 
rect 471 324 474 327 
rect 471 327 474 330 
rect 471 330 474 333 
rect 471 333 474 336 
rect 471 336 474 339 
rect 471 339 474 342 
rect 471 342 474 345 
rect 471 345 474 348 
rect 471 348 474 351 
rect 471 351 474 354 
rect 471 354 474 357 
rect 471 357 474 360 
rect 471 360 474 363 
rect 471 363 474 366 
rect 471 366 474 369 
rect 471 369 474 372 
rect 471 372 474 375 
rect 471 375 474 378 
rect 471 378 474 381 
rect 471 381 474 384 
rect 471 384 474 387 
rect 471 387 474 390 
rect 471 390 474 393 
rect 471 393 474 396 
rect 471 396 474 399 
rect 471 399 474 402 
rect 471 402 474 405 
rect 471 405 474 408 
rect 471 408 474 411 
rect 471 411 474 414 
rect 471 414 474 417 
rect 471 417 474 420 
rect 471 420 474 423 
rect 471 423 474 426 
rect 471 426 474 429 
rect 471 429 474 432 
rect 471 432 474 435 
rect 471 435 474 438 
rect 471 438 474 441 
rect 471 441 474 444 
rect 471 444 474 447 
rect 471 447 474 450 
rect 471 450 474 453 
rect 471 453 474 456 
rect 471 456 474 459 
rect 471 459 474 462 
rect 471 462 474 465 
rect 471 465 474 468 
rect 471 468 474 471 
rect 471 471 474 474 
rect 471 474 474 477 
rect 471 477 474 480 
rect 471 480 474 483 
rect 471 483 474 486 
rect 471 486 474 489 
rect 471 489 474 492 
rect 471 492 474 495 
rect 471 495 474 498 
rect 471 498 474 501 
rect 471 501 474 504 
rect 471 504 474 507 
rect 471 507 474 510 
rect 474 0 477 3 
rect 474 3 477 6 
rect 474 6 477 9 
rect 474 9 477 12 
rect 474 12 477 15 
rect 474 15 477 18 
rect 474 18 477 21 
rect 474 21 477 24 
rect 474 24 477 27 
rect 474 27 477 30 
rect 474 30 477 33 
rect 474 33 477 36 
rect 474 36 477 39 
rect 474 39 477 42 
rect 474 42 477 45 
rect 474 45 477 48 
rect 474 48 477 51 
rect 474 51 477 54 
rect 474 54 477 57 
rect 474 57 477 60 
rect 474 60 477 63 
rect 474 63 477 66 
rect 474 66 477 69 
rect 474 69 477 72 
rect 474 72 477 75 
rect 474 75 477 78 
rect 474 78 477 81 
rect 474 81 477 84 
rect 474 84 477 87 
rect 474 87 477 90 
rect 474 90 477 93 
rect 474 93 477 96 
rect 474 96 477 99 
rect 474 99 477 102 
rect 474 102 477 105 
rect 474 105 477 108 
rect 474 108 477 111 
rect 474 111 477 114 
rect 474 114 477 117 
rect 474 117 477 120 
rect 474 120 477 123 
rect 474 123 477 126 
rect 474 126 477 129 
rect 474 129 477 132 
rect 474 132 477 135 
rect 474 135 477 138 
rect 474 138 477 141 
rect 474 141 477 144 
rect 474 144 477 147 
rect 474 147 477 150 
rect 474 150 477 153 
rect 474 153 477 156 
rect 474 156 477 159 
rect 474 159 477 162 
rect 474 162 477 165 
rect 474 165 477 168 
rect 474 168 477 171 
rect 474 171 477 174 
rect 474 174 477 177 
rect 474 177 477 180 
rect 474 180 477 183 
rect 474 183 477 186 
rect 474 186 477 189 
rect 474 189 477 192 
rect 474 192 477 195 
rect 474 195 477 198 
rect 474 198 477 201 
rect 474 201 477 204 
rect 474 204 477 207 
rect 474 207 477 210 
rect 474 210 477 213 
rect 474 213 477 216 
rect 474 216 477 219 
rect 474 219 477 222 
rect 474 222 477 225 
rect 474 225 477 228 
rect 474 228 477 231 
rect 474 231 477 234 
rect 474 234 477 237 
rect 474 237 477 240 
rect 474 240 477 243 
rect 474 243 477 246 
rect 474 246 477 249 
rect 474 249 477 252 
rect 474 252 477 255 
rect 474 255 477 258 
rect 474 258 477 261 
rect 474 261 477 264 
rect 474 264 477 267 
rect 474 267 477 270 
rect 474 270 477 273 
rect 474 273 477 276 
rect 474 276 477 279 
rect 474 279 477 282 
rect 474 282 477 285 
rect 474 285 477 288 
rect 474 288 477 291 
rect 474 291 477 294 
rect 474 294 477 297 
rect 474 297 477 300 
rect 474 300 477 303 
rect 474 303 477 306 
rect 474 306 477 309 
rect 474 309 477 312 
rect 474 312 477 315 
rect 474 315 477 318 
rect 474 318 477 321 
rect 474 321 477 324 
rect 474 324 477 327 
rect 474 327 477 330 
rect 474 330 477 333 
rect 474 333 477 336 
rect 474 336 477 339 
rect 474 339 477 342 
rect 474 342 477 345 
rect 474 345 477 348 
rect 474 348 477 351 
rect 474 351 477 354 
rect 474 354 477 357 
rect 474 357 477 360 
rect 474 360 477 363 
rect 474 363 477 366 
rect 474 366 477 369 
rect 474 369 477 372 
rect 474 372 477 375 
rect 474 375 477 378 
rect 474 378 477 381 
rect 474 381 477 384 
rect 474 384 477 387 
rect 474 387 477 390 
rect 474 390 477 393 
rect 474 393 477 396 
rect 474 396 477 399 
rect 474 399 477 402 
rect 474 402 477 405 
rect 474 405 477 408 
rect 474 408 477 411 
rect 474 411 477 414 
rect 474 414 477 417 
rect 474 417 477 420 
rect 474 420 477 423 
rect 474 423 477 426 
rect 474 426 477 429 
rect 474 429 477 432 
rect 474 432 477 435 
rect 474 435 477 438 
rect 474 438 477 441 
rect 474 441 477 444 
rect 474 444 477 447 
rect 474 447 477 450 
rect 474 450 477 453 
rect 474 453 477 456 
rect 474 456 477 459 
rect 474 459 477 462 
rect 474 462 477 465 
rect 474 465 477 468 
rect 474 468 477 471 
rect 474 471 477 474 
rect 474 474 477 477 
rect 474 477 477 480 
rect 474 480 477 483 
rect 474 483 477 486 
rect 474 486 477 489 
rect 474 489 477 492 
rect 474 492 477 495 
rect 474 495 477 498 
rect 474 498 477 501 
rect 474 501 477 504 
rect 474 504 477 507 
rect 474 507 477 510 
rect 477 0 480 3 
rect 477 3 480 6 
rect 477 6 480 9 
rect 477 9 480 12 
rect 477 12 480 15 
rect 477 15 480 18 
rect 477 18 480 21 
rect 477 21 480 24 
rect 477 24 480 27 
rect 477 27 480 30 
rect 477 30 480 33 
rect 477 33 480 36 
rect 477 36 480 39 
rect 477 39 480 42 
rect 477 42 480 45 
rect 477 45 480 48 
rect 477 48 480 51 
rect 477 51 480 54 
rect 477 54 480 57 
rect 477 57 480 60 
rect 477 60 480 63 
rect 477 63 480 66 
rect 477 66 480 69 
rect 477 69 480 72 
rect 477 72 480 75 
rect 477 75 480 78 
rect 477 78 480 81 
rect 477 81 480 84 
rect 477 84 480 87 
rect 477 87 480 90 
rect 477 90 480 93 
rect 477 93 480 96 
rect 477 96 480 99 
rect 477 99 480 102 
rect 477 102 480 105 
rect 477 105 480 108 
rect 477 108 480 111 
rect 477 111 480 114 
rect 477 114 480 117 
rect 477 117 480 120 
rect 477 120 480 123 
rect 477 123 480 126 
rect 477 126 480 129 
rect 477 129 480 132 
rect 477 132 480 135 
rect 477 135 480 138 
rect 477 138 480 141 
rect 477 141 480 144 
rect 477 144 480 147 
rect 477 147 480 150 
rect 477 150 480 153 
rect 477 153 480 156 
rect 477 156 480 159 
rect 477 159 480 162 
rect 477 162 480 165 
rect 477 165 480 168 
rect 477 168 480 171 
rect 477 171 480 174 
rect 477 174 480 177 
rect 477 177 480 180 
rect 477 180 480 183 
rect 477 183 480 186 
rect 477 186 480 189 
rect 477 189 480 192 
rect 477 192 480 195 
rect 477 195 480 198 
rect 477 198 480 201 
rect 477 201 480 204 
rect 477 204 480 207 
rect 477 207 480 210 
rect 477 210 480 213 
rect 477 213 480 216 
rect 477 216 480 219 
rect 477 219 480 222 
rect 477 222 480 225 
rect 477 228 480 231 
rect 477 231 480 234 
rect 477 234 480 237 
rect 477 237 480 240 
rect 477 240 480 243 
rect 477 243 480 246 
rect 477 246 480 249 
rect 477 249 480 252 
rect 477 252 480 255 
rect 477 255 480 258 
rect 477 258 480 261 
rect 477 261 480 264 
rect 477 264 480 267 
rect 477 267 480 270 
rect 477 270 480 273 
rect 477 273 480 276 
rect 477 276 480 279 
rect 477 279 480 282 
rect 477 282 480 285 
rect 477 285 480 288 
rect 477 288 480 291 
rect 477 291 480 294 
rect 477 294 480 297 
rect 477 297 480 300 
rect 477 300 480 303 
rect 477 303 480 306 
rect 477 306 480 309 
rect 477 309 480 312 
rect 477 312 480 315 
rect 477 315 480 318 
rect 477 318 480 321 
rect 477 321 480 324 
rect 477 324 480 327 
rect 477 327 480 330 
rect 477 333 480 336 
rect 477 336 480 339 
rect 477 339 480 342 
rect 477 342 480 345 
rect 477 345 480 348 
rect 477 348 480 351 
rect 477 351 480 354 
rect 477 354 480 357 
rect 477 357 480 360 
rect 477 360 480 363 
rect 477 363 480 366 
rect 477 366 480 369 
rect 477 372 480 375 
rect 477 375 480 378 
rect 477 378 480 381 
rect 477 381 480 384 
rect 477 384 480 387 
rect 477 387 480 390 
rect 477 390 480 393 
rect 477 393 480 396 
rect 477 396 480 399 
rect 477 399 480 402 
rect 477 402 480 405 
rect 477 405 480 408 
rect 477 408 480 411 
rect 477 411 480 414 
rect 477 414 480 417 
rect 477 417 480 420 
rect 477 420 480 423 
rect 477 423 480 426 
rect 477 426 480 429 
rect 477 429 480 432 
rect 477 432 480 435 
rect 477 435 480 438 
rect 477 438 480 441 
rect 477 441 480 444 
rect 477 444 480 447 
rect 477 447 480 450 
rect 477 450 480 453 
rect 477 453 480 456 
rect 477 456 480 459 
rect 477 459 480 462 
rect 477 462 480 465 
rect 477 465 480 468 
rect 477 468 480 471 
rect 477 471 480 474 
rect 477 474 480 477 
rect 477 477 480 480 
rect 477 480 480 483 
rect 477 483 480 486 
rect 477 486 480 489 
rect 477 489 480 492 
rect 477 492 480 495 
rect 477 495 480 498 
rect 477 498 480 501 
rect 477 501 480 504 
rect 477 504 480 507 
rect 477 507 480 510 
rect 480 0 483 3 
rect 480 3 483 6 
rect 480 6 483 9 
rect 480 9 483 12 
rect 480 12 483 15 
rect 480 15 483 18 
rect 480 18 483 21 
rect 480 21 483 24 
rect 480 24 483 27 
rect 480 27 483 30 
rect 480 30 483 33 
rect 480 33 483 36 
rect 480 36 483 39 
rect 480 39 483 42 
rect 480 42 483 45 
rect 480 45 483 48 
rect 480 48 483 51 
rect 480 51 483 54 
rect 480 54 483 57 
rect 480 57 483 60 
rect 480 60 483 63 
rect 480 63 483 66 
rect 480 66 483 69 
rect 480 69 483 72 
rect 480 72 483 75 
rect 480 75 483 78 
rect 480 78 483 81 
rect 480 81 483 84 
rect 480 84 483 87 
rect 480 87 483 90 
rect 480 90 483 93 
rect 480 93 483 96 
rect 480 96 483 99 
rect 480 99 483 102 
rect 480 102 483 105 
rect 480 105 483 108 
rect 480 108 483 111 
rect 480 111 483 114 
rect 480 114 483 117 
rect 480 117 483 120 
rect 480 120 483 123 
rect 480 123 483 126 
rect 480 126 483 129 
rect 480 129 483 132 
rect 480 132 483 135 
rect 480 135 483 138 
rect 480 138 483 141 
rect 480 141 483 144 
rect 480 144 483 147 
rect 480 147 483 150 
rect 480 150 483 153 
rect 480 153 483 156 
rect 480 156 483 159 
rect 480 159 483 162 
rect 480 162 483 165 
rect 480 165 483 168 
rect 480 168 483 171 
rect 480 171 483 174 
rect 480 174 483 177 
rect 480 177 483 180 
rect 480 180 483 183 
rect 480 183 483 186 
rect 480 186 483 189 
rect 480 189 483 192 
rect 480 192 483 195 
rect 480 195 483 198 
rect 480 198 483 201 
rect 480 201 483 204 
rect 480 204 483 207 
rect 480 207 483 210 
rect 480 210 483 213 
rect 480 213 483 216 
rect 480 216 483 219 
rect 480 219 483 222 
rect 480 222 483 225 
rect 480 225 483 228 
rect 480 228 483 231 
rect 480 231 483 234 
rect 480 234 483 237 
rect 480 237 483 240 
rect 480 240 483 243 
rect 480 243 483 246 
rect 480 246 483 249 
rect 480 249 483 252 
rect 480 252 483 255 
rect 480 255 483 258 
rect 480 258 483 261 
rect 480 261 483 264 
rect 480 264 483 267 
rect 480 267 483 270 
rect 480 270 483 273 
rect 480 273 483 276 
rect 480 276 483 279 
rect 480 279 483 282 
rect 480 282 483 285 
rect 480 285 483 288 
rect 480 288 483 291 
rect 480 291 483 294 
rect 480 294 483 297 
rect 480 297 483 300 
rect 480 300 483 303 
rect 480 303 483 306 
rect 480 306 483 309 
rect 480 309 483 312 
rect 480 312 483 315 
rect 480 315 483 318 
rect 480 318 483 321 
rect 480 321 483 324 
rect 480 324 483 327 
rect 480 327 483 330 
rect 480 330 483 333 
rect 480 333 483 336 
rect 480 336 483 339 
rect 480 339 483 342 
rect 480 342 483 345 
rect 480 345 483 348 
rect 480 348 483 351 
rect 480 351 483 354 
rect 480 354 483 357 
rect 480 357 483 360 
rect 480 360 483 363 
rect 480 363 483 366 
rect 480 366 483 369 
rect 480 369 483 372 
rect 480 372 483 375 
rect 480 375 483 378 
rect 480 378 483 381 
rect 480 381 483 384 
rect 480 384 483 387 
rect 480 387 483 390 
rect 480 390 483 393 
rect 480 393 483 396 
rect 480 396 483 399 
rect 480 399 483 402 
rect 480 402 483 405 
rect 480 405 483 408 
rect 480 408 483 411 
rect 480 411 483 414 
rect 480 414 483 417 
rect 480 417 483 420 
rect 480 420 483 423 
rect 480 423 483 426 
rect 480 426 483 429 
rect 480 429 483 432 
rect 480 432 483 435 
rect 480 435 483 438 
rect 480 438 483 441 
rect 480 441 483 444 
rect 480 444 483 447 
rect 480 447 483 450 
rect 480 450 483 453 
rect 480 453 483 456 
rect 480 456 483 459 
rect 480 459 483 462 
rect 480 462 483 465 
rect 480 465 483 468 
rect 480 468 483 471 
rect 480 471 483 474 
rect 480 474 483 477 
rect 480 477 483 480 
rect 480 480 483 483 
rect 480 483 483 486 
rect 480 486 483 489 
rect 480 489 483 492 
rect 480 492 483 495 
rect 480 495 483 498 
rect 480 498 483 501 
rect 480 501 483 504 
rect 480 504 483 507 
rect 480 507 483 510 
rect 483 0 486 3 
rect 483 3 486 6 
rect 483 6 486 9 
rect 483 9 486 12 
rect 483 12 486 15 
rect 483 15 486 18 
rect 483 18 486 21 
rect 483 21 486 24 
rect 483 24 486 27 
rect 483 27 486 30 
rect 483 30 486 33 
rect 483 33 486 36 
rect 483 36 486 39 
rect 483 39 486 42 
rect 483 42 486 45 
rect 483 45 486 48 
rect 483 48 486 51 
rect 483 51 486 54 
rect 483 54 486 57 
rect 483 57 486 60 
rect 483 60 486 63 
rect 483 63 486 66 
rect 483 66 486 69 
rect 483 69 486 72 
rect 483 72 486 75 
rect 483 75 486 78 
rect 483 78 486 81 
rect 483 81 486 84 
rect 483 84 486 87 
rect 483 87 486 90 
rect 483 90 486 93 
rect 483 93 486 96 
rect 483 96 486 99 
rect 483 99 486 102 
rect 483 102 486 105 
rect 483 105 486 108 
rect 483 108 486 111 
rect 483 111 486 114 
rect 483 114 486 117 
rect 483 117 486 120 
rect 483 120 486 123 
rect 483 123 486 126 
rect 483 126 486 129 
rect 483 129 486 132 
rect 483 132 486 135 
rect 483 135 486 138 
rect 483 138 486 141 
rect 483 141 486 144 
rect 483 144 486 147 
rect 483 147 486 150 
rect 483 150 486 153 
rect 483 153 486 156 
rect 483 156 486 159 
rect 483 159 486 162 
rect 483 162 486 165 
rect 483 165 486 168 
rect 483 168 486 171 
rect 483 171 486 174 
rect 483 174 486 177 
rect 483 177 486 180 
rect 483 180 486 183 
rect 483 183 486 186 
rect 483 186 486 189 
rect 483 189 486 192 
rect 483 192 486 195 
rect 483 195 486 198 
rect 483 198 486 201 
rect 483 201 486 204 
rect 483 204 486 207 
rect 483 207 486 210 
rect 483 210 486 213 
rect 483 213 486 216 
rect 483 216 486 219 
rect 483 219 486 222 
rect 483 222 486 225 
rect 483 225 486 228 
rect 483 228 486 231 
rect 483 231 486 234 
rect 483 234 486 237 
rect 483 237 486 240 
rect 483 240 486 243 
rect 483 243 486 246 
rect 483 246 486 249 
rect 483 249 486 252 
rect 483 252 486 255 
rect 483 255 486 258 
rect 483 258 486 261 
rect 483 261 486 264 
rect 483 264 486 267 
rect 483 267 486 270 
rect 483 270 486 273 
rect 483 273 486 276 
rect 483 276 486 279 
rect 483 279 486 282 
rect 483 282 486 285 
rect 483 285 486 288 
rect 483 288 486 291 
rect 483 291 486 294 
rect 483 294 486 297 
rect 483 297 486 300 
rect 483 300 486 303 
rect 483 303 486 306 
rect 483 306 486 309 
rect 483 309 486 312 
rect 483 312 486 315 
rect 483 315 486 318 
rect 483 318 486 321 
rect 483 321 486 324 
rect 483 324 486 327 
rect 483 327 486 330 
rect 483 330 486 333 
rect 483 333 486 336 
rect 483 336 486 339 
rect 483 339 486 342 
rect 483 342 486 345 
rect 483 345 486 348 
rect 483 348 486 351 
rect 483 351 486 354 
rect 483 354 486 357 
rect 483 357 486 360 
rect 483 360 486 363 
rect 483 363 486 366 
rect 483 366 486 369 
rect 483 369 486 372 
rect 483 372 486 375 
rect 483 375 486 378 
rect 483 378 486 381 
rect 483 381 486 384 
rect 483 384 486 387 
rect 483 387 486 390 
rect 483 390 486 393 
rect 483 393 486 396 
rect 483 396 486 399 
rect 483 399 486 402 
rect 483 402 486 405 
rect 483 405 486 408 
rect 483 408 486 411 
rect 483 411 486 414 
rect 483 414 486 417 
rect 483 417 486 420 
rect 483 420 486 423 
rect 483 423 486 426 
rect 483 426 486 429 
rect 483 429 486 432 
rect 483 432 486 435 
rect 483 435 486 438 
rect 483 438 486 441 
rect 483 441 486 444 
rect 483 444 486 447 
rect 483 447 486 450 
rect 483 450 486 453 
rect 483 453 486 456 
rect 483 456 486 459 
rect 483 459 486 462 
rect 483 462 486 465 
rect 483 465 486 468 
rect 483 468 486 471 
rect 483 471 486 474 
rect 483 474 486 477 
rect 483 477 486 480 
rect 483 480 486 483 
rect 483 483 486 486 
rect 483 486 486 489 
rect 483 489 486 492 
rect 483 492 486 495 
rect 483 495 486 498 
rect 483 498 486 501 
rect 483 501 486 504 
rect 483 504 486 507 
rect 483 507 486 510 
rect 486 0 489 3 
rect 486 3 489 6 
rect 486 6 489 9 
rect 486 9 489 12 
rect 486 12 489 15 
rect 486 15 489 18 
rect 486 18 489 21 
rect 486 21 489 24 
rect 486 24 489 27 
rect 486 27 489 30 
rect 486 30 489 33 
rect 486 33 489 36 
rect 486 36 489 39 
rect 486 39 489 42 
rect 486 42 489 45 
rect 486 45 489 48 
rect 486 48 489 51 
rect 486 51 489 54 
rect 486 54 489 57 
rect 486 57 489 60 
rect 486 60 489 63 
rect 486 63 489 66 
rect 486 66 489 69 
rect 486 69 489 72 
rect 486 72 489 75 
rect 486 75 489 78 
rect 486 78 489 81 
rect 486 81 489 84 
rect 486 84 489 87 
rect 486 87 489 90 
rect 486 90 489 93 
rect 486 93 489 96 
rect 486 96 489 99 
rect 486 99 489 102 
rect 486 102 489 105 
rect 486 105 489 108 
rect 486 108 489 111 
rect 486 111 489 114 
rect 486 114 489 117 
rect 486 117 489 120 
rect 486 120 489 123 
rect 486 123 489 126 
rect 486 126 489 129 
rect 486 129 489 132 
rect 486 132 489 135 
rect 486 135 489 138 
rect 486 138 489 141 
rect 486 141 489 144 
rect 486 144 489 147 
rect 486 147 489 150 
rect 486 150 489 153 
rect 486 153 489 156 
rect 486 156 489 159 
rect 486 159 489 162 
rect 486 162 489 165 
rect 486 165 489 168 
rect 486 168 489 171 
rect 486 171 489 174 
rect 486 174 489 177 
rect 486 177 489 180 
rect 486 180 489 183 
rect 486 183 489 186 
rect 486 186 489 189 
rect 486 189 489 192 
rect 486 192 489 195 
rect 486 195 489 198 
rect 486 198 489 201 
rect 486 201 489 204 
rect 486 204 489 207 
rect 486 207 489 210 
rect 486 210 489 213 
rect 486 213 489 216 
rect 486 216 489 219 
rect 486 219 489 222 
rect 486 222 489 225 
rect 486 225 489 228 
rect 486 228 489 231 
rect 486 231 489 234 
rect 486 234 489 237 
rect 486 237 489 240 
rect 486 240 489 243 
rect 486 243 489 246 
rect 486 246 489 249 
rect 486 249 489 252 
rect 486 252 489 255 
rect 486 255 489 258 
rect 486 258 489 261 
rect 486 261 489 264 
rect 486 264 489 267 
rect 486 267 489 270 
rect 486 270 489 273 
rect 486 273 489 276 
rect 486 276 489 279 
rect 486 279 489 282 
rect 486 282 489 285 
rect 486 285 489 288 
rect 486 288 489 291 
rect 486 291 489 294 
rect 486 294 489 297 
rect 486 297 489 300 
rect 486 300 489 303 
rect 486 303 489 306 
rect 486 306 489 309 
rect 486 309 489 312 
rect 486 312 489 315 
rect 486 315 489 318 
rect 486 318 489 321 
rect 486 321 489 324 
rect 486 324 489 327 
rect 486 327 489 330 
rect 486 330 489 333 
rect 486 333 489 336 
rect 486 336 489 339 
rect 486 339 489 342 
rect 486 342 489 345 
rect 486 345 489 348 
rect 486 348 489 351 
rect 486 351 489 354 
rect 486 354 489 357 
rect 486 357 489 360 
rect 486 360 489 363 
rect 486 363 489 366 
rect 486 366 489 369 
rect 486 369 489 372 
rect 486 372 489 375 
rect 486 375 489 378 
rect 486 378 489 381 
rect 486 381 489 384 
rect 486 384 489 387 
rect 486 387 489 390 
rect 486 390 489 393 
rect 486 393 489 396 
rect 486 396 489 399 
rect 486 399 489 402 
rect 486 402 489 405 
rect 486 405 489 408 
rect 486 408 489 411 
rect 486 411 489 414 
rect 486 414 489 417 
rect 486 417 489 420 
rect 486 420 489 423 
rect 486 423 489 426 
rect 486 426 489 429 
rect 486 429 489 432 
rect 486 432 489 435 
rect 486 435 489 438 
rect 486 438 489 441 
rect 486 441 489 444 
rect 486 444 489 447 
rect 486 447 489 450 
rect 486 450 489 453 
rect 486 453 489 456 
rect 486 456 489 459 
rect 486 459 489 462 
rect 486 462 489 465 
rect 486 465 489 468 
rect 486 468 489 471 
rect 486 471 489 474 
rect 486 474 489 477 
rect 486 477 489 480 
rect 486 480 489 483 
rect 486 483 489 486 
rect 486 486 489 489 
rect 486 489 489 492 
rect 486 492 489 495 
rect 486 495 489 498 
rect 486 498 489 501 
rect 486 501 489 504 
rect 486 504 489 507 
rect 486 507 489 510 
rect 489 0 492 3 
rect 489 3 492 6 
rect 489 6 492 9 
rect 489 9 492 12 
rect 489 12 492 15 
rect 489 15 492 18 
rect 489 18 492 21 
rect 489 21 492 24 
rect 489 24 492 27 
rect 489 27 492 30 
rect 489 30 492 33 
rect 489 33 492 36 
rect 489 36 492 39 
rect 489 39 492 42 
rect 489 42 492 45 
rect 489 45 492 48 
rect 489 48 492 51 
rect 489 51 492 54 
rect 489 54 492 57 
rect 489 57 492 60 
rect 489 60 492 63 
rect 489 63 492 66 
rect 489 66 492 69 
rect 489 69 492 72 
rect 489 72 492 75 
rect 489 75 492 78 
rect 489 78 492 81 
rect 489 81 492 84 
rect 489 84 492 87 
rect 489 87 492 90 
rect 489 90 492 93 
rect 489 93 492 96 
rect 489 96 492 99 
rect 489 99 492 102 
rect 489 102 492 105 
rect 489 105 492 108 
rect 489 108 492 111 
rect 489 111 492 114 
rect 489 114 492 117 
rect 489 117 492 120 
rect 489 120 492 123 
rect 489 123 492 126 
rect 489 126 492 129 
rect 489 129 492 132 
rect 489 132 492 135 
rect 489 135 492 138 
rect 489 138 492 141 
rect 489 141 492 144 
rect 489 144 492 147 
rect 489 147 492 150 
rect 489 150 492 153 
rect 489 153 492 156 
rect 489 156 492 159 
rect 489 159 492 162 
rect 489 162 492 165 
rect 489 165 492 168 
rect 489 168 492 171 
rect 489 171 492 174 
rect 489 174 492 177 
rect 489 177 492 180 
rect 489 180 492 183 
rect 489 183 492 186 
rect 489 186 492 189 
rect 489 189 492 192 
rect 489 192 492 195 
rect 489 195 492 198 
rect 489 198 492 201 
rect 489 201 492 204 
rect 489 204 492 207 
rect 489 207 492 210 
rect 489 210 492 213 
rect 489 213 492 216 
rect 489 216 492 219 
rect 489 219 492 222 
rect 489 222 492 225 
rect 489 225 492 228 
rect 489 228 492 231 
rect 489 231 492 234 
rect 489 234 492 237 
rect 489 237 492 240 
rect 489 240 492 243 
rect 489 243 492 246 
rect 489 246 492 249 
rect 489 249 492 252 
rect 489 252 492 255 
rect 489 255 492 258 
rect 489 258 492 261 
rect 489 261 492 264 
rect 489 264 492 267 
rect 489 267 492 270 
rect 489 270 492 273 
rect 489 273 492 276 
rect 489 276 492 279 
rect 489 279 492 282 
rect 489 282 492 285 
rect 489 285 492 288 
rect 489 288 492 291 
rect 489 291 492 294 
rect 489 294 492 297 
rect 489 297 492 300 
rect 489 300 492 303 
rect 489 303 492 306 
rect 489 306 492 309 
rect 489 309 492 312 
rect 489 312 492 315 
rect 489 315 492 318 
rect 489 318 492 321 
rect 489 321 492 324 
rect 489 324 492 327 
rect 489 327 492 330 
rect 489 330 492 333 
rect 489 333 492 336 
rect 489 336 492 339 
rect 489 339 492 342 
rect 489 342 492 345 
rect 489 345 492 348 
rect 489 348 492 351 
rect 489 351 492 354 
rect 489 354 492 357 
rect 489 357 492 360 
rect 489 360 492 363 
rect 489 363 492 366 
rect 489 366 492 369 
rect 489 369 492 372 
rect 489 372 492 375 
rect 489 375 492 378 
rect 489 378 492 381 
rect 489 381 492 384 
rect 489 384 492 387 
rect 489 387 492 390 
rect 489 390 492 393 
rect 489 393 492 396 
rect 489 396 492 399 
rect 489 399 492 402 
rect 489 402 492 405 
rect 489 405 492 408 
rect 489 408 492 411 
rect 489 411 492 414 
rect 489 414 492 417 
rect 489 417 492 420 
rect 489 420 492 423 
rect 489 423 492 426 
rect 489 426 492 429 
rect 489 429 492 432 
rect 489 432 492 435 
rect 489 435 492 438 
rect 489 438 492 441 
rect 489 441 492 444 
rect 489 444 492 447 
rect 489 447 492 450 
rect 489 450 492 453 
rect 489 453 492 456 
rect 489 456 492 459 
rect 489 459 492 462 
rect 489 462 492 465 
rect 489 465 492 468 
rect 489 468 492 471 
rect 489 471 492 474 
rect 489 474 492 477 
rect 489 477 492 480 
rect 489 480 492 483 
rect 489 483 492 486 
rect 489 486 492 489 
rect 489 489 492 492 
rect 489 492 492 495 
rect 489 495 492 498 
rect 489 498 492 501 
rect 489 501 492 504 
rect 489 504 492 507 
rect 489 507 492 510 
rect 492 0 495 3 
rect 492 3 495 6 
rect 492 6 495 9 
rect 492 9 495 12 
rect 492 12 495 15 
rect 492 15 495 18 
rect 492 18 495 21 
rect 492 21 495 24 
rect 492 24 495 27 
rect 492 27 495 30 
rect 492 30 495 33 
rect 492 33 495 36 
rect 492 36 495 39 
rect 492 39 495 42 
rect 492 42 495 45 
rect 492 45 495 48 
rect 492 48 495 51 
rect 492 51 495 54 
rect 492 54 495 57 
rect 492 57 495 60 
rect 492 60 495 63 
rect 492 63 495 66 
rect 492 66 495 69 
rect 492 69 495 72 
rect 492 72 495 75 
rect 492 75 495 78 
rect 492 78 495 81 
rect 492 81 495 84 
rect 492 84 495 87 
rect 492 87 495 90 
rect 492 90 495 93 
rect 492 93 495 96 
rect 492 96 495 99 
rect 492 99 495 102 
rect 492 102 495 105 
rect 492 105 495 108 
rect 492 108 495 111 
rect 492 111 495 114 
rect 492 114 495 117 
rect 492 117 495 120 
rect 492 120 495 123 
rect 492 123 495 126 
rect 492 126 495 129 
rect 492 129 495 132 
rect 492 132 495 135 
rect 492 135 495 138 
rect 492 138 495 141 
rect 492 141 495 144 
rect 492 144 495 147 
rect 492 147 495 150 
rect 492 150 495 153 
rect 492 153 495 156 
rect 492 156 495 159 
rect 492 159 495 162 
rect 492 162 495 165 
rect 492 165 495 168 
rect 492 168 495 171 
rect 492 171 495 174 
rect 492 174 495 177 
rect 492 177 495 180 
rect 492 180 495 183 
rect 492 183 495 186 
rect 492 186 495 189 
rect 492 189 495 192 
rect 492 192 495 195 
rect 492 195 495 198 
rect 492 198 495 201 
rect 492 201 495 204 
rect 492 204 495 207 
rect 492 207 495 210 
rect 492 210 495 213 
rect 492 213 495 216 
rect 492 216 495 219 
rect 492 219 495 222 
rect 492 222 495 225 
rect 492 225 495 228 
rect 492 228 495 231 
rect 492 231 495 234 
rect 492 234 495 237 
rect 492 237 495 240 
rect 492 240 495 243 
rect 492 243 495 246 
rect 492 246 495 249 
rect 492 249 495 252 
rect 492 252 495 255 
rect 492 255 495 258 
rect 492 258 495 261 
rect 492 261 495 264 
rect 492 264 495 267 
rect 492 267 495 270 
rect 492 270 495 273 
rect 492 273 495 276 
rect 492 276 495 279 
rect 492 279 495 282 
rect 492 282 495 285 
rect 492 285 495 288 
rect 492 288 495 291 
rect 492 291 495 294 
rect 492 294 495 297 
rect 492 297 495 300 
rect 492 300 495 303 
rect 492 303 495 306 
rect 492 306 495 309 
rect 492 309 495 312 
rect 492 312 495 315 
rect 492 315 495 318 
rect 492 318 495 321 
rect 492 321 495 324 
rect 492 324 495 327 
rect 492 327 495 330 
rect 492 330 495 333 
rect 492 333 495 336 
rect 492 336 495 339 
rect 492 339 495 342 
rect 492 342 495 345 
rect 492 345 495 348 
rect 492 348 495 351 
rect 492 351 495 354 
rect 492 354 495 357 
rect 492 357 495 360 
rect 492 360 495 363 
rect 492 363 495 366 
rect 492 366 495 369 
rect 492 369 495 372 
rect 492 372 495 375 
rect 492 375 495 378 
rect 492 378 495 381 
rect 492 381 495 384 
rect 492 384 495 387 
rect 492 387 495 390 
rect 492 390 495 393 
rect 492 393 495 396 
rect 492 396 495 399 
rect 492 399 495 402 
rect 492 402 495 405 
rect 492 405 495 408 
rect 492 408 495 411 
rect 492 411 495 414 
rect 492 414 495 417 
rect 492 417 495 420 
rect 492 420 495 423 
rect 492 423 495 426 
rect 492 426 495 429 
rect 492 429 495 432 
rect 492 432 495 435 
rect 492 435 495 438 
rect 492 438 495 441 
rect 492 441 495 444 
rect 492 444 495 447 
rect 492 447 495 450 
rect 492 450 495 453 
rect 492 453 495 456 
rect 492 456 495 459 
rect 492 459 495 462 
rect 492 462 495 465 
rect 492 465 495 468 
rect 492 468 495 471 
rect 492 471 495 474 
rect 492 474 495 477 
rect 492 477 495 480 
rect 492 480 495 483 
rect 492 483 495 486 
rect 492 486 495 489 
rect 492 489 495 492 
rect 492 492 495 495 
rect 492 495 495 498 
rect 492 498 495 501 
rect 492 501 495 504 
rect 492 504 495 507 
rect 492 507 495 510 
rect 495 0 498 3 
rect 495 3 498 6 
rect 495 6 498 9 
rect 495 9 498 12 
rect 495 12 498 15 
rect 495 15 498 18 
rect 495 18 498 21 
rect 495 21 498 24 
rect 495 24 498 27 
rect 495 27 498 30 
rect 495 30 498 33 
rect 495 33 498 36 
rect 495 36 498 39 
rect 495 39 498 42 
rect 495 42 498 45 
rect 495 45 498 48 
rect 495 48 498 51 
rect 495 51 498 54 
rect 495 54 498 57 
rect 495 57 498 60 
rect 495 60 498 63 
rect 495 63 498 66 
rect 495 66 498 69 
rect 495 69 498 72 
rect 495 72 498 75 
rect 495 75 498 78 
rect 495 78 498 81 
rect 495 81 498 84 
rect 495 84 498 87 
rect 495 87 498 90 
rect 495 90 498 93 
rect 495 93 498 96 
rect 495 96 498 99 
rect 495 99 498 102 
rect 495 102 498 105 
rect 495 105 498 108 
rect 495 108 498 111 
rect 495 111 498 114 
rect 495 114 498 117 
rect 495 117 498 120 
rect 495 120 498 123 
rect 495 123 498 126 
rect 495 126 498 129 
rect 495 129 498 132 
rect 495 132 498 135 
rect 495 135 498 138 
rect 495 138 498 141 
rect 495 141 498 144 
rect 495 144 498 147 
rect 495 147 498 150 
rect 495 150 498 153 
rect 495 153 498 156 
rect 495 156 498 159 
rect 495 159 498 162 
rect 495 162 498 165 
rect 495 165 498 168 
rect 495 168 498 171 
rect 495 171 498 174 
rect 495 174 498 177 
rect 495 177 498 180 
rect 495 180 498 183 
rect 495 183 498 186 
rect 495 186 498 189 
rect 495 189 498 192 
rect 495 192 498 195 
rect 495 195 498 198 
rect 495 198 498 201 
rect 495 201 498 204 
rect 495 204 498 207 
rect 495 207 498 210 
rect 495 210 498 213 
rect 495 213 498 216 
rect 495 216 498 219 
rect 495 219 498 222 
rect 495 222 498 225 
rect 495 225 498 228 
rect 495 228 498 231 
rect 495 231 498 234 
rect 495 234 498 237 
rect 495 237 498 240 
rect 495 240 498 243 
rect 495 243 498 246 
rect 495 246 498 249 
rect 495 249 498 252 
rect 495 252 498 255 
rect 495 255 498 258 
rect 495 258 498 261 
rect 495 261 498 264 
rect 495 264 498 267 
rect 495 267 498 270 
rect 495 270 498 273 
rect 495 273 498 276 
rect 495 276 498 279 
rect 495 279 498 282 
rect 495 282 498 285 
rect 495 285 498 288 
rect 495 288 498 291 
rect 495 291 498 294 
rect 495 294 498 297 
rect 495 297 498 300 
rect 495 300 498 303 
rect 495 303 498 306 
rect 495 306 498 309 
rect 495 309 498 312 
rect 495 312 498 315 
rect 495 315 498 318 
rect 495 318 498 321 
rect 495 321 498 324 
rect 495 324 498 327 
rect 495 327 498 330 
rect 495 330 498 333 
rect 495 333 498 336 
rect 495 336 498 339 
rect 495 339 498 342 
rect 495 342 498 345 
rect 495 345 498 348 
rect 495 348 498 351 
rect 495 351 498 354 
rect 495 354 498 357 
rect 495 357 498 360 
rect 495 360 498 363 
rect 495 363 498 366 
rect 495 366 498 369 
rect 495 369 498 372 
rect 495 372 498 375 
rect 495 375 498 378 
rect 495 378 498 381 
rect 495 381 498 384 
rect 495 384 498 387 
rect 495 387 498 390 
rect 495 390 498 393 
rect 495 393 498 396 
rect 495 396 498 399 
rect 495 399 498 402 
rect 495 402 498 405 
rect 495 405 498 408 
rect 495 408 498 411 
rect 495 411 498 414 
rect 495 414 498 417 
rect 495 417 498 420 
rect 495 420 498 423 
rect 495 423 498 426 
rect 495 426 498 429 
rect 495 429 498 432 
rect 495 432 498 435 
rect 495 435 498 438 
rect 495 438 498 441 
rect 495 441 498 444 
rect 495 444 498 447 
rect 495 447 498 450 
rect 495 450 498 453 
rect 495 453 498 456 
rect 495 456 498 459 
rect 495 459 498 462 
rect 495 462 498 465 
rect 495 465 498 468 
rect 495 468 498 471 
rect 495 471 498 474 
rect 495 474 498 477 
rect 495 477 498 480 
rect 495 480 498 483 
rect 495 483 498 486 
rect 495 486 498 489 
rect 495 489 498 492 
rect 495 492 498 495 
rect 495 495 498 498 
rect 495 498 498 501 
rect 495 501 498 504 
rect 495 504 498 507 
rect 495 507 498 510 
rect 498 0 501 3 
rect 498 3 501 6 
rect 498 6 501 9 
rect 498 9 501 12 
rect 498 12 501 15 
rect 498 15 501 18 
rect 498 18 501 21 
rect 498 21 501 24 
rect 498 24 501 27 
rect 498 27 501 30 
rect 498 30 501 33 
rect 498 33 501 36 
rect 498 36 501 39 
rect 498 39 501 42 
rect 498 42 501 45 
rect 498 45 501 48 
rect 498 48 501 51 
rect 498 51 501 54 
rect 498 54 501 57 
rect 498 57 501 60 
rect 498 60 501 63 
rect 498 63 501 66 
rect 498 66 501 69 
rect 498 69 501 72 
rect 498 72 501 75 
rect 498 75 501 78 
rect 498 78 501 81 
rect 498 81 501 84 
rect 498 84 501 87 
rect 498 87 501 90 
rect 498 90 501 93 
rect 498 93 501 96 
rect 498 96 501 99 
rect 498 99 501 102 
rect 498 102 501 105 
rect 498 105 501 108 
rect 498 108 501 111 
rect 498 111 501 114 
rect 498 114 501 117 
rect 498 117 501 120 
rect 498 120 501 123 
rect 498 123 501 126 
rect 498 126 501 129 
rect 498 129 501 132 
rect 498 132 501 135 
rect 498 135 501 138 
rect 498 138 501 141 
rect 498 141 501 144 
rect 498 144 501 147 
rect 498 147 501 150 
rect 498 150 501 153 
rect 498 153 501 156 
rect 498 156 501 159 
rect 498 159 501 162 
rect 498 162 501 165 
rect 498 165 501 168 
rect 498 168 501 171 
rect 498 171 501 174 
rect 498 174 501 177 
rect 498 177 501 180 
rect 498 180 501 183 
rect 498 183 501 186 
rect 498 186 501 189 
rect 498 189 501 192 
rect 498 192 501 195 
rect 498 195 501 198 
rect 498 198 501 201 
rect 498 201 501 204 
rect 498 204 501 207 
rect 498 207 501 210 
rect 498 210 501 213 
rect 498 213 501 216 
rect 498 216 501 219 
rect 498 219 501 222 
rect 498 222 501 225 
rect 498 225 501 228 
rect 498 228 501 231 
rect 498 231 501 234 
rect 498 234 501 237 
rect 498 237 501 240 
rect 498 240 501 243 
rect 498 243 501 246 
rect 498 246 501 249 
rect 498 249 501 252 
rect 498 252 501 255 
rect 498 255 501 258 
rect 498 258 501 261 
rect 498 261 501 264 
rect 498 264 501 267 
rect 498 267 501 270 
rect 498 270 501 273 
rect 498 273 501 276 
rect 498 276 501 279 
rect 498 279 501 282 
rect 498 282 501 285 
rect 498 285 501 288 
rect 498 288 501 291 
rect 498 291 501 294 
rect 498 294 501 297 
rect 498 297 501 300 
rect 498 300 501 303 
rect 498 303 501 306 
rect 498 306 501 309 
rect 498 309 501 312 
rect 498 312 501 315 
rect 498 315 501 318 
rect 498 318 501 321 
rect 498 321 501 324 
rect 498 324 501 327 
rect 498 327 501 330 
rect 498 330 501 333 
rect 498 333 501 336 
rect 498 336 501 339 
rect 498 339 501 342 
rect 498 342 501 345 
rect 498 345 501 348 
rect 498 348 501 351 
rect 498 351 501 354 
rect 498 354 501 357 
rect 498 357 501 360 
rect 498 360 501 363 
rect 498 363 501 366 
rect 498 366 501 369 
rect 498 369 501 372 
rect 498 372 501 375 
rect 498 375 501 378 
rect 498 378 501 381 
rect 498 381 501 384 
rect 498 384 501 387 
rect 498 387 501 390 
rect 498 390 501 393 
rect 498 393 501 396 
rect 498 396 501 399 
rect 498 399 501 402 
rect 498 402 501 405 
rect 498 405 501 408 
rect 498 408 501 411 
rect 498 411 501 414 
rect 498 414 501 417 
rect 498 417 501 420 
rect 498 420 501 423 
rect 498 423 501 426 
rect 498 426 501 429 
rect 498 429 501 432 
rect 498 432 501 435 
rect 498 435 501 438 
rect 498 438 501 441 
rect 498 441 501 444 
rect 498 444 501 447 
rect 498 447 501 450 
rect 498 450 501 453 
rect 498 453 501 456 
rect 498 456 501 459 
rect 498 459 501 462 
rect 498 462 501 465 
rect 498 465 501 468 
rect 498 468 501 471 
rect 498 471 501 474 
rect 498 474 501 477 
rect 498 477 501 480 
rect 498 480 501 483 
rect 498 483 501 486 
rect 498 486 501 489 
rect 498 489 501 492 
rect 498 492 501 495 
rect 498 495 501 498 
rect 498 498 501 501 
rect 498 501 501 504 
rect 498 504 501 507 
rect 498 507 501 510 
rect 501 0 504 3 
rect 501 3 504 6 
rect 501 6 504 9 
rect 501 9 504 12 
rect 501 12 504 15 
rect 501 15 504 18 
rect 501 18 504 21 
rect 501 21 504 24 
rect 501 24 504 27 
rect 501 27 504 30 
rect 501 30 504 33 
rect 501 33 504 36 
rect 501 36 504 39 
rect 501 39 504 42 
rect 501 42 504 45 
rect 501 45 504 48 
rect 501 48 504 51 
rect 501 51 504 54 
rect 501 54 504 57 
rect 501 57 504 60 
rect 501 60 504 63 
rect 501 63 504 66 
rect 501 66 504 69 
rect 501 69 504 72 
rect 501 72 504 75 
rect 501 75 504 78 
rect 501 78 504 81 
rect 501 81 504 84 
rect 501 84 504 87 
rect 501 87 504 90 
rect 501 90 504 93 
rect 501 93 504 96 
rect 501 96 504 99 
rect 501 99 504 102 
rect 501 102 504 105 
rect 501 105 504 108 
rect 501 108 504 111 
rect 501 111 504 114 
rect 501 114 504 117 
rect 501 117 504 120 
rect 501 120 504 123 
rect 501 123 504 126 
rect 501 126 504 129 
rect 501 129 504 132 
rect 501 132 504 135 
rect 501 135 504 138 
rect 501 138 504 141 
rect 501 141 504 144 
rect 501 144 504 147 
rect 501 147 504 150 
rect 501 150 504 153 
rect 501 153 504 156 
rect 501 156 504 159 
rect 501 159 504 162 
rect 501 162 504 165 
rect 501 165 504 168 
rect 501 168 504 171 
rect 501 171 504 174 
rect 501 174 504 177 
rect 501 177 504 180 
rect 501 180 504 183 
rect 501 183 504 186 
rect 501 186 504 189 
rect 501 189 504 192 
rect 501 192 504 195 
rect 501 195 504 198 
rect 501 198 504 201 
rect 501 201 504 204 
rect 501 204 504 207 
rect 501 207 504 210 
rect 501 210 504 213 
rect 501 213 504 216 
rect 501 216 504 219 
rect 501 219 504 222 
rect 501 222 504 225 
rect 501 225 504 228 
rect 501 228 504 231 
rect 501 231 504 234 
rect 501 234 504 237 
rect 501 237 504 240 
rect 501 240 504 243 
rect 501 243 504 246 
rect 501 246 504 249 
rect 501 249 504 252 
rect 501 252 504 255 
rect 501 255 504 258 
rect 501 258 504 261 
rect 501 261 504 264 
rect 501 264 504 267 
rect 501 267 504 270 
rect 501 270 504 273 
rect 501 273 504 276 
rect 501 276 504 279 
rect 501 279 504 282 
rect 501 282 504 285 
rect 501 285 504 288 
rect 501 288 504 291 
rect 501 291 504 294 
rect 501 294 504 297 
rect 501 297 504 300 
rect 501 300 504 303 
rect 501 303 504 306 
rect 501 306 504 309 
rect 501 309 504 312 
rect 501 312 504 315 
rect 501 315 504 318 
rect 501 318 504 321 
rect 501 321 504 324 
rect 501 324 504 327 
rect 501 327 504 330 
rect 501 330 504 333 
rect 501 333 504 336 
rect 501 336 504 339 
rect 501 339 504 342 
rect 501 342 504 345 
rect 501 345 504 348 
rect 501 348 504 351 
rect 501 351 504 354 
rect 501 354 504 357 
rect 501 357 504 360 
rect 501 360 504 363 
rect 501 363 504 366 
rect 501 366 504 369 
rect 501 369 504 372 
rect 501 372 504 375 
rect 501 375 504 378 
rect 501 378 504 381 
rect 501 381 504 384 
rect 501 384 504 387 
rect 501 387 504 390 
rect 501 390 504 393 
rect 501 393 504 396 
rect 501 396 504 399 
rect 501 399 504 402 
rect 501 402 504 405 
rect 501 405 504 408 
rect 501 408 504 411 
rect 501 411 504 414 
rect 501 414 504 417 
rect 501 417 504 420 
rect 501 420 504 423 
rect 501 423 504 426 
rect 501 426 504 429 
rect 501 429 504 432 
rect 501 432 504 435 
rect 501 435 504 438 
rect 501 438 504 441 
rect 501 441 504 444 
rect 501 444 504 447 
rect 501 447 504 450 
rect 501 450 504 453 
rect 501 453 504 456 
rect 501 456 504 459 
rect 501 459 504 462 
rect 501 462 504 465 
rect 501 465 504 468 
rect 501 468 504 471 
rect 501 471 504 474 
rect 501 474 504 477 
rect 501 477 504 480 
rect 501 480 504 483 
rect 501 483 504 486 
rect 501 486 504 489 
rect 501 489 504 492 
rect 501 492 504 495 
rect 501 495 504 498 
rect 501 498 504 501 
rect 501 501 504 504 
rect 501 504 504 507 
rect 501 507 504 510 
rect 504 0 507 3 
rect 504 3 507 6 
rect 504 6 507 9 
rect 504 9 507 12 
rect 504 12 507 15 
rect 504 15 507 18 
rect 504 18 507 21 
rect 504 21 507 24 
rect 504 24 507 27 
rect 504 27 507 30 
rect 504 30 507 33 
rect 504 33 507 36 
rect 504 36 507 39 
rect 504 39 507 42 
rect 504 42 507 45 
rect 504 45 507 48 
rect 504 48 507 51 
rect 504 51 507 54 
rect 504 54 507 57 
rect 504 57 507 60 
rect 504 60 507 63 
rect 504 63 507 66 
rect 504 66 507 69 
rect 504 69 507 72 
rect 504 72 507 75 
rect 504 75 507 78 
rect 504 78 507 81 
rect 504 81 507 84 
rect 504 84 507 87 
rect 504 87 507 90 
rect 504 90 507 93 
rect 504 93 507 96 
rect 504 96 507 99 
rect 504 99 507 102 
rect 504 102 507 105 
rect 504 105 507 108 
rect 504 108 507 111 
rect 504 111 507 114 
rect 504 114 507 117 
rect 504 117 507 120 
rect 504 120 507 123 
rect 504 123 507 126 
rect 504 126 507 129 
rect 504 129 507 132 
rect 504 132 507 135 
rect 504 135 507 138 
rect 504 138 507 141 
rect 504 141 507 144 
rect 504 144 507 147 
rect 504 147 507 150 
rect 504 150 507 153 
rect 504 153 507 156 
rect 504 156 507 159 
rect 504 159 507 162 
rect 504 162 507 165 
rect 504 165 507 168 
rect 504 168 507 171 
rect 504 171 507 174 
rect 504 174 507 177 
rect 504 177 507 180 
rect 504 180 507 183 
rect 504 183 507 186 
rect 504 186 507 189 
rect 504 189 507 192 
rect 504 192 507 195 
rect 504 195 507 198 
rect 504 198 507 201 
rect 504 201 507 204 
rect 504 204 507 207 
rect 504 207 507 210 
rect 504 210 507 213 
rect 504 213 507 216 
rect 504 216 507 219 
rect 504 219 507 222 
rect 504 222 507 225 
rect 504 225 507 228 
rect 504 228 507 231 
rect 504 231 507 234 
rect 504 234 507 237 
rect 504 237 507 240 
rect 504 240 507 243 
rect 504 243 507 246 
rect 504 246 507 249 
rect 504 249 507 252 
rect 504 252 507 255 
rect 504 255 507 258 
rect 504 258 507 261 
rect 504 261 507 264 
rect 504 264 507 267 
rect 504 267 507 270 
rect 504 270 507 273 
rect 504 273 507 276 
rect 504 276 507 279 
rect 504 279 507 282 
rect 504 282 507 285 
rect 504 285 507 288 
rect 504 288 507 291 
rect 504 291 507 294 
rect 504 294 507 297 
rect 504 297 507 300 
rect 504 300 507 303 
rect 504 303 507 306 
rect 504 306 507 309 
rect 504 309 507 312 
rect 504 312 507 315 
rect 504 315 507 318 
rect 504 318 507 321 
rect 504 321 507 324 
rect 504 324 507 327 
rect 504 327 507 330 
rect 504 330 507 333 
rect 504 333 507 336 
rect 504 336 507 339 
rect 504 339 507 342 
rect 504 342 507 345 
rect 504 345 507 348 
rect 504 348 507 351 
rect 504 351 507 354 
rect 504 354 507 357 
rect 504 357 507 360 
rect 504 360 507 363 
rect 504 363 507 366 
rect 504 366 507 369 
rect 504 369 507 372 
rect 504 372 507 375 
rect 504 375 507 378 
rect 504 378 507 381 
rect 504 381 507 384 
rect 504 384 507 387 
rect 504 387 507 390 
rect 504 390 507 393 
rect 504 393 507 396 
rect 504 396 507 399 
rect 504 399 507 402 
rect 504 402 507 405 
rect 504 405 507 408 
rect 504 408 507 411 
rect 504 411 507 414 
rect 504 414 507 417 
rect 504 417 507 420 
rect 504 420 507 423 
rect 504 423 507 426 
rect 504 426 507 429 
rect 504 429 507 432 
rect 504 432 507 435 
rect 504 435 507 438 
rect 504 438 507 441 
rect 504 441 507 444 
rect 504 444 507 447 
rect 504 447 507 450 
rect 504 450 507 453 
rect 504 453 507 456 
rect 504 456 507 459 
rect 504 459 507 462 
rect 504 462 507 465 
rect 504 465 507 468 
rect 504 468 507 471 
rect 504 471 507 474 
rect 504 474 507 477 
rect 504 477 507 480 
rect 504 480 507 483 
rect 504 483 507 486 
rect 504 486 507 489 
rect 504 489 507 492 
rect 504 492 507 495 
rect 504 495 507 498 
rect 504 498 507 501 
rect 504 501 507 504 
rect 504 504 507 507 
rect 504 507 507 510 
rect 507 0 510 3 
rect 507 3 510 6 
rect 507 6 510 9 
rect 507 9 510 12 
rect 507 12 510 15 
rect 507 15 510 18 
rect 507 18 510 21 
rect 507 21 510 24 
rect 507 24 510 27 
rect 507 27 510 30 
rect 507 30 510 33 
rect 507 33 510 36 
rect 507 36 510 39 
rect 507 39 510 42 
rect 507 42 510 45 
rect 507 45 510 48 
rect 507 48 510 51 
rect 507 51 510 54 
rect 507 54 510 57 
rect 507 57 510 60 
rect 507 60 510 63 
rect 507 63 510 66 
rect 507 66 510 69 
rect 507 69 510 72 
rect 507 72 510 75 
rect 507 75 510 78 
rect 507 78 510 81 
rect 507 81 510 84 
rect 507 84 510 87 
rect 507 87 510 90 
rect 507 90 510 93 
rect 507 93 510 96 
rect 507 96 510 99 
rect 507 99 510 102 
rect 507 102 510 105 
rect 507 105 510 108 
rect 507 108 510 111 
rect 507 111 510 114 
rect 507 114 510 117 
rect 507 117 510 120 
rect 507 120 510 123 
rect 507 123 510 126 
rect 507 126 510 129 
rect 507 129 510 132 
rect 507 132 510 135 
rect 507 135 510 138 
rect 507 138 510 141 
rect 507 141 510 144 
rect 507 144 510 147 
rect 507 147 510 150 
rect 507 150 510 153 
rect 507 153 510 156 
rect 507 156 510 159 
rect 507 159 510 162 
rect 507 162 510 165 
rect 507 165 510 168 
rect 507 168 510 171 
rect 507 171 510 174 
rect 507 174 510 177 
rect 507 177 510 180 
rect 507 180 510 183 
rect 507 183 510 186 
rect 507 186 510 189 
rect 507 189 510 192 
rect 507 192 510 195 
rect 507 195 510 198 
rect 507 198 510 201 
rect 507 201 510 204 
rect 507 204 510 207 
rect 507 207 510 210 
rect 507 210 510 213 
rect 507 213 510 216 
rect 507 216 510 219 
rect 507 219 510 222 
rect 507 222 510 225 
rect 507 225 510 228 
rect 507 228 510 231 
rect 507 231 510 234 
rect 507 234 510 237 
rect 507 237 510 240 
rect 507 240 510 243 
rect 507 243 510 246 
rect 507 246 510 249 
rect 507 249 510 252 
rect 507 252 510 255 
rect 507 255 510 258 
rect 507 258 510 261 
rect 507 261 510 264 
rect 507 264 510 267 
rect 507 267 510 270 
rect 507 270 510 273 
rect 507 273 510 276 
rect 507 276 510 279 
rect 507 279 510 282 
rect 507 282 510 285 
rect 507 285 510 288 
rect 507 288 510 291 
rect 507 291 510 294 
rect 507 294 510 297 
rect 507 297 510 300 
rect 507 300 510 303 
rect 507 303 510 306 
rect 507 306 510 309 
rect 507 309 510 312 
rect 507 312 510 315 
rect 507 315 510 318 
rect 507 318 510 321 
rect 507 321 510 324 
rect 507 324 510 327 
rect 507 327 510 330 
rect 507 330 510 333 
rect 507 333 510 336 
rect 507 336 510 339 
rect 507 339 510 342 
rect 507 342 510 345 
rect 507 345 510 348 
rect 507 348 510 351 
rect 507 351 510 354 
rect 507 354 510 357 
rect 507 357 510 360 
rect 507 360 510 363 
rect 507 363 510 366 
rect 507 366 510 369 
rect 507 369 510 372 
rect 507 372 510 375 
rect 507 375 510 378 
rect 507 378 510 381 
rect 507 381 510 384 
rect 507 384 510 387 
rect 507 387 510 390 
rect 507 390 510 393 
rect 507 393 510 396 
rect 507 396 510 399 
rect 507 399 510 402 
rect 507 402 510 405 
rect 507 405 510 408 
rect 507 408 510 411 
rect 507 411 510 414 
rect 507 414 510 417 
rect 507 417 510 420 
rect 507 420 510 423 
rect 507 423 510 426 
rect 507 426 510 429 
rect 507 429 510 432 
rect 507 432 510 435 
rect 507 435 510 438 
rect 507 438 510 441 
rect 507 441 510 444 
rect 507 444 510 447 
rect 507 447 510 450 
rect 507 450 510 453 
rect 507 453 510 456 
rect 507 456 510 459 
rect 507 459 510 462 
rect 507 462 510 465 
rect 507 465 510 468 
rect 507 468 510 471 
rect 507 471 510 474 
rect 507 474 510 477 
rect 507 477 510 480 
rect 507 480 510 483 
rect 507 483 510 486 
rect 507 486 510 489 
rect 507 489 510 492 
rect 507 492 510 495 
rect 507 495 510 498 
rect 507 498 510 501 
rect 507 501 510 504 
rect 507 504 510 507 
rect 507 507 510 510 
<< labels >>
<< metal1 >>
rect 0 0 3 3 
rect 0 3 3 6 
rect 0 6 3 9 
rect 0 9 3 12 
rect 0 12 3 15 
rect 0 15 3 18 
rect 0 18 3 21 
rect 0 21 3 24 
rect 0 24 3 27 
rect 0 27 3 30 
rect 0 30 3 33 
rect 0 33 3 36 
rect 0 36 3 39 
rect 0 39 3 42 
rect 0 42 3 45 
rect 0 45 3 48 
rect 0 48 3 51 
rect 0 51 3 54 
rect 0 54 3 57 
rect 0 57 3 60 
rect 0 60 3 63 
rect 0 63 3 66 
rect 0 66 3 69 
rect 0 69 3 72 
rect 0 72 3 75 
rect 0 75 3 78 
rect 0 78 3 81 
rect 0 81 3 84 
rect 0 84 3 87 
rect 0 87 3 90 
rect 0 90 3 93 
rect 0 93 3 96 
rect 0 96 3 99 
rect 0 99 3 102 
rect 0 102 3 105 
rect 0 105 3 108 
rect 0 108 3 111 
rect 0 111 3 114 
rect 0 114 3 117 
rect 0 117 3 120 
rect 0 120 3 123 
rect 0 123 3 126 
rect 0 126 3 129 
rect 0 129 3 132 
rect 0 132 3 135 
rect 0 135 3 138 
rect 0 138 3 141 
rect 0 141 3 144 
rect 0 144 3 147 
rect 0 147 3 150 
rect 0 150 3 153 
rect 0 153 3 156 
rect 0 156 3 159 
rect 0 159 3 162 
rect 0 162 3 165 
rect 0 165 3 168 
rect 0 168 3 171 
rect 0 171 3 174 
rect 0 174 3 177 
rect 0 177 3 180 
rect 0 180 3 183 
rect 0 183 3 186 
rect 0 186 3 189 
rect 0 189 3 192 
rect 0 192 3 195 
rect 0 195 3 198 
rect 0 198 3 201 
rect 0 201 3 204 
rect 0 204 3 207 
rect 0 207 3 210 
rect 0 210 3 213 
rect 0 213 3 216 
rect 0 216 3 219 
rect 0 219 3 222 
rect 0 222 3 225 
rect 0 225 3 228 
rect 0 228 3 231 
rect 0 231 3 234 
rect 0 234 3 237 
rect 0 237 3 240 
rect 0 240 3 243 
rect 0 243 3 246 
rect 0 246 3 249 
rect 0 249 3 252 
rect 0 252 3 255 
rect 0 255 3 258 
rect 0 258 3 261 
rect 0 261 3 264 
rect 0 264 3 267 
rect 0 267 3 270 
rect 0 270 3 273 
rect 0 273 3 276 
rect 0 276 3 279 
rect 0 279 3 282 
rect 0 282 3 285 
rect 0 285 3 288 
rect 0 288 3 291 
rect 0 291 3 294 
rect 0 294 3 297 
rect 0 297 3 300 
rect 0 300 3 303 
rect 0 303 3 306 
rect 0 306 3 309 
rect 0 309 3 312 
rect 0 312 3 315 
rect 0 315 3 318 
rect 0 318 3 321 
rect 0 321 3 324 
rect 0 324 3 327 
rect 0 327 3 330 
rect 0 330 3 333 
rect 0 333 3 336 
rect 0 336 3 339 
rect 0 339 3 342 
rect 0 342 3 345 
rect 0 345 3 348 
rect 0 348 3 351 
rect 0 351 3 354 
rect 0 354 3 357 
rect 0 357 3 360 
rect 0 360 3 363 
rect 0 363 3 366 
rect 0 366 3 369 
rect 0 369 3 372 
rect 0 372 3 375 
rect 0 375 3 378 
rect 0 378 3 381 
rect 0 381 3 384 
rect 0 384 3 387 
rect 0 387 3 390 
rect 0 390 3 393 
rect 0 393 3 396 
rect 0 396 3 399 
rect 0 399 3 402 
rect 0 402 3 405 
rect 0 405 3 408 
rect 0 408 3 411 
rect 0 411 3 414 
rect 0 414 3 417 
rect 0 417 3 420 
rect 0 420 3 423 
rect 0 423 3 426 
rect 0 426 3 429 
rect 0 429 3 432 
rect 0 432 3 435 
rect 0 435 3 438 
rect 0 438 3 441 
rect 0 441 3 444 
rect 0 444 3 447 
rect 0 447 3 450 
rect 0 450 3 453 
rect 0 453 3 456 
rect 0 456 3 459 
rect 0 459 3 462 
rect 0 462 3 465 
rect 0 465 3 468 
rect 0 468 3 471 
rect 0 471 3 474 
rect 0 474 3 477 
rect 0 477 3 480 
rect 0 480 3 483 
rect 0 483 3 486 
rect 0 486 3 489 
rect 0 489 3 492 
rect 0 492 3 495 
rect 0 495 3 498 
rect 0 498 3 501 
rect 0 501 3 504 
rect 0 504 3 507 
rect 0 507 3 510 
rect 3 0 6 3 
rect 3 3 6 6 
rect 3 6 6 9 
rect 3 9 6 12 
rect 3 12 6 15 
rect 3 15 6 18 
rect 3 18 6 21 
rect 3 21 6 24 
rect 3 24 6 27 
rect 3 27 6 30 
rect 3 30 6 33 
rect 3 33 6 36 
rect 3 36 6 39 
rect 3 39 6 42 
rect 3 42 6 45 
rect 3 45 6 48 
rect 3 48 6 51 
rect 3 51 6 54 
rect 3 54 6 57 
rect 3 57 6 60 
rect 3 60 6 63 
rect 3 63 6 66 
rect 3 66 6 69 
rect 3 69 6 72 
rect 3 72 6 75 
rect 3 75 6 78 
rect 3 78 6 81 
rect 3 81 6 84 
rect 3 84 6 87 
rect 3 87 6 90 
rect 3 90 6 93 
rect 3 93 6 96 
rect 3 96 6 99 
rect 3 99 6 102 
rect 3 102 6 105 
rect 3 105 6 108 
rect 3 108 6 111 
rect 3 111 6 114 
rect 3 114 6 117 
rect 3 117 6 120 
rect 3 120 6 123 
rect 3 123 6 126 
rect 3 126 6 129 
rect 3 129 6 132 
rect 3 132 6 135 
rect 3 135 6 138 
rect 3 138 6 141 
rect 3 141 6 144 
rect 3 144 6 147 
rect 3 147 6 150 
rect 3 150 6 153 
rect 3 153 6 156 
rect 3 156 6 159 
rect 3 159 6 162 
rect 3 162 6 165 
rect 3 165 6 168 
rect 3 168 6 171 
rect 3 171 6 174 
rect 3 174 6 177 
rect 3 177 6 180 
rect 3 180 6 183 
rect 3 183 6 186 
rect 3 186 6 189 
rect 3 189 6 192 
rect 3 192 6 195 
rect 3 195 6 198 
rect 3 198 6 201 
rect 3 201 6 204 
rect 3 204 6 207 
rect 3 207 6 210 
rect 3 210 6 213 
rect 3 213 6 216 
rect 3 216 6 219 
rect 3 219 6 222 
rect 3 222 6 225 
rect 3 225 6 228 
rect 3 228 6 231 
rect 3 231 6 234 
rect 3 234 6 237 
rect 3 237 6 240 
rect 3 240 6 243 
rect 3 243 6 246 
rect 3 246 6 249 
rect 3 249 6 252 
rect 3 252 6 255 
rect 3 255 6 258 
rect 3 258 6 261 
rect 3 261 6 264 
rect 3 264 6 267 
rect 3 267 6 270 
rect 3 270 6 273 
rect 3 273 6 276 
rect 3 276 6 279 
rect 3 279 6 282 
rect 3 282 6 285 
rect 3 285 6 288 
rect 3 288 6 291 
rect 3 291 6 294 
rect 3 294 6 297 
rect 3 297 6 300 
rect 3 300 6 303 
rect 3 303 6 306 
rect 3 306 6 309 
rect 3 309 6 312 
rect 3 312 6 315 
rect 3 315 6 318 
rect 3 318 6 321 
rect 3 321 6 324 
rect 3 324 6 327 
rect 3 327 6 330 
rect 3 330 6 333 
rect 3 333 6 336 
rect 3 336 6 339 
rect 3 339 6 342 
rect 3 342 6 345 
rect 3 345 6 348 
rect 3 348 6 351 
rect 3 351 6 354 
rect 3 354 6 357 
rect 3 357 6 360 
rect 3 360 6 363 
rect 3 363 6 366 
rect 3 366 6 369 
rect 3 369 6 372 
rect 3 372 6 375 
rect 3 375 6 378 
rect 3 378 6 381 
rect 3 381 6 384 
rect 3 384 6 387 
rect 3 387 6 390 
rect 3 390 6 393 
rect 3 393 6 396 
rect 3 396 6 399 
rect 3 399 6 402 
rect 3 402 6 405 
rect 3 405 6 408 
rect 3 408 6 411 
rect 3 411 6 414 
rect 3 414 6 417 
rect 3 417 6 420 
rect 3 420 6 423 
rect 3 423 6 426 
rect 3 426 6 429 
rect 3 429 6 432 
rect 3 432 6 435 
rect 3 435 6 438 
rect 3 438 6 441 
rect 3 441 6 444 
rect 3 444 6 447 
rect 3 447 6 450 
rect 3 450 6 453 
rect 3 453 6 456 
rect 3 456 6 459 
rect 3 459 6 462 
rect 3 462 6 465 
rect 3 465 6 468 
rect 3 468 6 471 
rect 3 471 6 474 
rect 3 474 6 477 
rect 3 477 6 480 
rect 3 480 6 483 
rect 3 483 6 486 
rect 3 486 6 489 
rect 3 489 6 492 
rect 3 492 6 495 
rect 3 495 6 498 
rect 3 498 6 501 
rect 3 501 6 504 
rect 3 504 6 507 
rect 3 507 6 510 
rect 6 0 9 3 
rect 6 3 9 6 
rect 6 6 9 9 
rect 6 9 9 12 
rect 6 12 9 15 
rect 6 15 9 18 
rect 6 18 9 21 
rect 6 21 9 24 
rect 6 24 9 27 
rect 6 27 9 30 
rect 6 30 9 33 
rect 6 33 9 36 
rect 6 36 9 39 
rect 6 39 9 42 
rect 6 42 9 45 
rect 6 45 9 48 
rect 6 48 9 51 
rect 6 51 9 54 
rect 6 54 9 57 
rect 6 57 9 60 
rect 6 60 9 63 
rect 6 63 9 66 
rect 6 66 9 69 
rect 6 69 9 72 
rect 6 72 9 75 
rect 6 75 9 78 
rect 6 78 9 81 
rect 6 81 9 84 
rect 6 84 9 87 
rect 6 87 9 90 
rect 6 90 9 93 
rect 6 93 9 96 
rect 6 96 9 99 
rect 6 99 9 102 
rect 6 102 9 105 
rect 6 105 9 108 
rect 6 108 9 111 
rect 6 111 9 114 
rect 6 114 9 117 
rect 6 117 9 120 
rect 6 120 9 123 
rect 6 123 9 126 
rect 6 126 9 129 
rect 6 129 9 132 
rect 6 132 9 135 
rect 6 135 9 138 
rect 6 138 9 141 
rect 6 141 9 144 
rect 6 144 9 147 
rect 6 147 9 150 
rect 6 150 9 153 
rect 6 153 9 156 
rect 6 156 9 159 
rect 6 159 9 162 
rect 6 162 9 165 
rect 6 165 9 168 
rect 6 168 9 171 
rect 6 171 9 174 
rect 6 174 9 177 
rect 6 177 9 180 
rect 6 180 9 183 
rect 6 183 9 186 
rect 6 186 9 189 
rect 6 189 9 192 
rect 6 192 9 195 
rect 6 195 9 198 
rect 6 198 9 201 
rect 6 201 9 204 
rect 6 204 9 207 
rect 6 207 9 210 
rect 6 210 9 213 
rect 6 213 9 216 
rect 6 216 9 219 
rect 6 219 9 222 
rect 6 222 9 225 
rect 6 225 9 228 
rect 6 228 9 231 
rect 6 231 9 234 
rect 6 234 9 237 
rect 6 237 9 240 
rect 6 240 9 243 
rect 6 243 9 246 
rect 6 246 9 249 
rect 6 249 9 252 
rect 6 252 9 255 
rect 6 255 9 258 
rect 6 258 9 261 
rect 6 261 9 264 
rect 6 264 9 267 
rect 6 267 9 270 
rect 6 270 9 273 
rect 6 273 9 276 
rect 6 276 9 279 
rect 6 279 9 282 
rect 6 282 9 285 
rect 6 285 9 288 
rect 6 288 9 291 
rect 6 291 9 294 
rect 6 294 9 297 
rect 6 297 9 300 
rect 6 300 9 303 
rect 6 303 9 306 
rect 6 306 9 309 
rect 6 309 9 312 
rect 6 312 9 315 
rect 6 315 9 318 
rect 6 318 9 321 
rect 6 321 9 324 
rect 6 324 9 327 
rect 6 327 9 330 
rect 6 330 9 333 
rect 6 333 9 336 
rect 6 336 9 339 
rect 6 339 9 342 
rect 6 342 9 345 
rect 6 345 9 348 
rect 6 348 9 351 
rect 6 351 9 354 
rect 6 354 9 357 
rect 6 357 9 360 
rect 6 360 9 363 
rect 6 363 9 366 
rect 6 366 9 369 
rect 6 369 9 372 
rect 6 372 9 375 
rect 6 375 9 378 
rect 6 378 9 381 
rect 6 381 9 384 
rect 6 384 9 387 
rect 6 387 9 390 
rect 6 390 9 393 
rect 6 393 9 396 
rect 6 396 9 399 
rect 6 399 9 402 
rect 6 402 9 405 
rect 6 405 9 408 
rect 6 408 9 411 
rect 6 411 9 414 
rect 6 414 9 417 
rect 6 417 9 420 
rect 6 420 9 423 
rect 6 423 9 426 
rect 6 426 9 429 
rect 6 429 9 432 
rect 6 432 9 435 
rect 6 435 9 438 
rect 6 438 9 441 
rect 6 441 9 444 
rect 6 444 9 447 
rect 6 447 9 450 
rect 6 450 9 453 
rect 6 453 9 456 
rect 6 456 9 459 
rect 6 459 9 462 
rect 6 462 9 465 
rect 6 465 9 468 
rect 6 468 9 471 
rect 6 471 9 474 
rect 6 474 9 477 
rect 6 477 9 480 
rect 6 480 9 483 
rect 6 483 9 486 
rect 6 486 9 489 
rect 6 489 9 492 
rect 6 492 9 495 
rect 6 495 9 498 
rect 6 498 9 501 
rect 6 501 9 504 
rect 6 504 9 507 
rect 6 507 9 510 
rect 9 0 12 3 
rect 9 3 12 6 
rect 9 6 12 9 
rect 9 9 12 12 
rect 9 12 12 15 
rect 9 15 12 18 
rect 9 18 12 21 
rect 9 21 12 24 
rect 9 24 12 27 
rect 9 27 12 30 
rect 9 30 12 33 
rect 9 33 12 36 
rect 9 36 12 39 
rect 9 39 12 42 
rect 9 42 12 45 
rect 9 45 12 48 
rect 9 48 12 51 
rect 9 51 12 54 
rect 9 54 12 57 
rect 9 57 12 60 
rect 9 60 12 63 
rect 9 63 12 66 
rect 9 66 12 69 
rect 9 69 12 72 
rect 9 72 12 75 
rect 9 75 12 78 
rect 9 78 12 81 
rect 9 81 12 84 
rect 9 84 12 87 
rect 9 87 12 90 
rect 9 90 12 93 
rect 9 93 12 96 
rect 9 96 12 99 
rect 9 99 12 102 
rect 9 102 12 105 
rect 9 105 12 108 
rect 9 108 12 111 
rect 9 111 12 114 
rect 9 114 12 117 
rect 9 117 12 120 
rect 9 120 12 123 
rect 9 123 12 126 
rect 9 126 12 129 
rect 9 129 12 132 
rect 9 132 12 135 
rect 9 135 12 138 
rect 9 138 12 141 
rect 9 141 12 144 
rect 9 144 12 147 
rect 9 147 12 150 
rect 9 150 12 153 
rect 9 153 12 156 
rect 9 156 12 159 
rect 9 159 12 162 
rect 9 162 12 165 
rect 9 165 12 168 
rect 9 168 12 171 
rect 9 171 12 174 
rect 9 174 12 177 
rect 9 177 12 180 
rect 9 180 12 183 
rect 9 183 12 186 
rect 9 186 12 189 
rect 9 189 12 192 
rect 9 192 12 195 
rect 9 195 12 198 
rect 9 198 12 201 
rect 9 201 12 204 
rect 9 204 12 207 
rect 9 207 12 210 
rect 9 210 12 213 
rect 9 213 12 216 
rect 9 216 12 219 
rect 9 219 12 222 
rect 9 222 12 225 
rect 9 225 12 228 
rect 9 228 12 231 
rect 9 231 12 234 
rect 9 234 12 237 
rect 9 237 12 240 
rect 9 240 12 243 
rect 9 243 12 246 
rect 9 246 12 249 
rect 9 249 12 252 
rect 9 252 12 255 
rect 9 255 12 258 
rect 9 258 12 261 
rect 9 261 12 264 
rect 9 264 12 267 
rect 9 267 12 270 
rect 9 270 12 273 
rect 9 273 12 276 
rect 9 276 12 279 
rect 9 279 12 282 
rect 9 282 12 285 
rect 9 285 12 288 
rect 9 288 12 291 
rect 9 291 12 294 
rect 9 294 12 297 
rect 9 297 12 300 
rect 9 300 12 303 
rect 9 303 12 306 
rect 9 306 12 309 
rect 9 309 12 312 
rect 9 312 12 315 
rect 9 315 12 318 
rect 9 318 12 321 
rect 9 321 12 324 
rect 9 324 12 327 
rect 9 327 12 330 
rect 9 330 12 333 
rect 9 333 12 336 
rect 9 336 12 339 
rect 9 339 12 342 
rect 9 342 12 345 
rect 9 345 12 348 
rect 9 348 12 351 
rect 9 351 12 354 
rect 9 354 12 357 
rect 9 357 12 360 
rect 9 360 12 363 
rect 9 363 12 366 
rect 9 366 12 369 
rect 9 369 12 372 
rect 9 372 12 375 
rect 9 375 12 378 
rect 9 378 12 381 
rect 9 381 12 384 
rect 9 384 12 387 
rect 9 387 12 390 
rect 9 390 12 393 
rect 9 393 12 396 
rect 9 396 12 399 
rect 9 399 12 402 
rect 9 402 12 405 
rect 9 405 12 408 
rect 9 408 12 411 
rect 9 411 12 414 
rect 9 414 12 417 
rect 9 417 12 420 
rect 9 420 12 423 
rect 9 423 12 426 
rect 9 426 12 429 
rect 9 429 12 432 
rect 9 432 12 435 
rect 9 435 12 438 
rect 9 438 12 441 
rect 9 441 12 444 
rect 9 444 12 447 
rect 9 447 12 450 
rect 9 450 12 453 
rect 9 453 12 456 
rect 9 456 12 459 
rect 9 459 12 462 
rect 9 462 12 465 
rect 9 465 12 468 
rect 9 468 12 471 
rect 9 471 12 474 
rect 9 474 12 477 
rect 9 477 12 480 
rect 9 480 12 483 
rect 9 483 12 486 
rect 9 486 12 489 
rect 9 489 12 492 
rect 9 492 12 495 
rect 9 495 12 498 
rect 9 498 12 501 
rect 9 501 12 504 
rect 9 504 12 507 
rect 9 507 12 510 
rect 12 0 15 3 
rect 12 3 15 6 
rect 12 6 15 9 
rect 12 9 15 12 
rect 12 12 15 15 
rect 12 15 15 18 
rect 12 18 15 21 
rect 12 21 15 24 
rect 12 24 15 27 
rect 12 27 15 30 
rect 12 30 15 33 
rect 12 33 15 36 
rect 12 36 15 39 
rect 12 39 15 42 
rect 12 42 15 45 
rect 12 45 15 48 
rect 12 48 15 51 
rect 12 51 15 54 
rect 12 54 15 57 
rect 12 57 15 60 
rect 12 60 15 63 
rect 12 63 15 66 
rect 12 66 15 69 
rect 12 69 15 72 
rect 12 72 15 75 
rect 12 75 15 78 
rect 12 78 15 81 
rect 12 81 15 84 
rect 12 84 15 87 
rect 12 87 15 90 
rect 12 90 15 93 
rect 12 93 15 96 
rect 12 96 15 99 
rect 12 99 15 102 
rect 12 102 15 105 
rect 12 105 15 108 
rect 12 108 15 111 
rect 12 111 15 114 
rect 12 114 15 117 
rect 12 117 15 120 
rect 12 120 15 123 
rect 12 123 15 126 
rect 12 126 15 129 
rect 12 129 15 132 
rect 12 132 15 135 
rect 12 135 15 138 
rect 12 138 15 141 
rect 12 141 15 144 
rect 12 144 15 147 
rect 12 147 15 150 
rect 12 150 15 153 
rect 12 153 15 156 
rect 12 156 15 159 
rect 12 159 15 162 
rect 12 162 15 165 
rect 12 165 15 168 
rect 12 168 15 171 
rect 12 171 15 174 
rect 12 174 15 177 
rect 12 177 15 180 
rect 12 180 15 183 
rect 12 183 15 186 
rect 12 186 15 189 
rect 12 189 15 192 
rect 12 192 15 195 
rect 12 195 15 198 
rect 12 198 15 201 
rect 12 201 15 204 
rect 12 204 15 207 
rect 12 207 15 210 
rect 12 210 15 213 
rect 12 213 15 216 
rect 12 216 15 219 
rect 12 219 15 222 
rect 12 222 15 225 
rect 12 225 15 228 
rect 12 228 15 231 
rect 12 231 15 234 
rect 12 234 15 237 
rect 12 237 15 240 
rect 12 240 15 243 
rect 12 243 15 246 
rect 12 246 15 249 
rect 12 249 15 252 
rect 12 252 15 255 
rect 12 255 15 258 
rect 12 258 15 261 
rect 12 261 15 264 
rect 12 264 15 267 
rect 12 267 15 270 
rect 12 270 15 273 
rect 12 273 15 276 
rect 12 276 15 279 
rect 12 279 15 282 
rect 12 282 15 285 
rect 12 285 15 288 
rect 12 288 15 291 
rect 12 291 15 294 
rect 12 294 15 297 
rect 12 297 15 300 
rect 12 300 15 303 
rect 12 303 15 306 
rect 12 306 15 309 
rect 12 309 15 312 
rect 12 312 15 315 
rect 12 315 15 318 
rect 12 318 15 321 
rect 12 321 15 324 
rect 12 324 15 327 
rect 12 327 15 330 
rect 12 330 15 333 
rect 12 333 15 336 
rect 12 336 15 339 
rect 12 339 15 342 
rect 12 342 15 345 
rect 12 345 15 348 
rect 12 348 15 351 
rect 12 351 15 354 
rect 12 354 15 357 
rect 12 357 15 360 
rect 12 360 15 363 
rect 12 363 15 366 
rect 12 366 15 369 
rect 12 369 15 372 
rect 12 372 15 375 
rect 12 375 15 378 
rect 12 378 15 381 
rect 12 381 15 384 
rect 12 384 15 387 
rect 12 387 15 390 
rect 12 390 15 393 
rect 12 393 15 396 
rect 12 396 15 399 
rect 12 399 15 402 
rect 12 402 15 405 
rect 12 405 15 408 
rect 12 408 15 411 
rect 12 411 15 414 
rect 12 414 15 417 
rect 12 417 15 420 
rect 12 420 15 423 
rect 12 423 15 426 
rect 12 426 15 429 
rect 12 429 15 432 
rect 12 432 15 435 
rect 12 435 15 438 
rect 12 438 15 441 
rect 12 441 15 444 
rect 12 444 15 447 
rect 12 447 15 450 
rect 12 450 15 453 
rect 12 453 15 456 
rect 12 456 15 459 
rect 12 459 15 462 
rect 12 462 15 465 
rect 12 465 15 468 
rect 12 468 15 471 
rect 12 471 15 474 
rect 12 474 15 477 
rect 12 477 15 480 
rect 12 480 15 483 
rect 12 483 15 486 
rect 12 486 15 489 
rect 12 489 15 492 
rect 12 492 15 495 
rect 12 495 15 498 
rect 12 498 15 501 
rect 12 501 15 504 
rect 12 504 15 507 
rect 12 507 15 510 
rect 15 0 18 3 
rect 15 3 18 6 
rect 15 6 18 9 
rect 15 9 18 12 
rect 15 12 18 15 
rect 15 15 18 18 
rect 15 18 18 21 
rect 15 21 18 24 
rect 15 24 18 27 
rect 15 27 18 30 
rect 15 30 18 33 
rect 15 33 18 36 
rect 15 36 18 39 
rect 15 39 18 42 
rect 15 42 18 45 
rect 15 45 18 48 
rect 15 48 18 51 
rect 15 51 18 54 
rect 15 54 18 57 
rect 15 57 18 60 
rect 15 60 18 63 
rect 15 63 18 66 
rect 15 66 18 69 
rect 15 69 18 72 
rect 15 72 18 75 
rect 15 75 18 78 
rect 15 78 18 81 
rect 15 81 18 84 
rect 15 84 18 87 
rect 15 87 18 90 
rect 15 90 18 93 
rect 15 93 18 96 
rect 15 96 18 99 
rect 15 99 18 102 
rect 15 102 18 105 
rect 15 105 18 108 
rect 15 108 18 111 
rect 15 111 18 114 
rect 15 114 18 117 
rect 15 117 18 120 
rect 15 120 18 123 
rect 15 123 18 126 
rect 15 126 18 129 
rect 15 129 18 132 
rect 15 132 18 135 
rect 15 135 18 138 
rect 15 138 18 141 
rect 15 141 18 144 
rect 15 144 18 147 
rect 15 147 18 150 
rect 15 150 18 153 
rect 15 153 18 156 
rect 15 156 18 159 
rect 15 159 18 162 
rect 15 162 18 165 
rect 15 165 18 168 
rect 15 168 18 171 
rect 15 171 18 174 
rect 15 174 18 177 
rect 15 177 18 180 
rect 15 180 18 183 
rect 15 183 18 186 
rect 15 186 18 189 
rect 15 189 18 192 
rect 15 192 18 195 
rect 15 195 18 198 
rect 15 198 18 201 
rect 15 201 18 204 
rect 15 204 18 207 
rect 15 207 18 210 
rect 15 210 18 213 
rect 15 213 18 216 
rect 15 216 18 219 
rect 15 219 18 222 
rect 15 222 18 225 
rect 15 225 18 228 
rect 15 228 18 231 
rect 15 231 18 234 
rect 15 234 18 237 
rect 15 237 18 240 
rect 15 240 18 243 
rect 15 243 18 246 
rect 15 246 18 249 
rect 15 249 18 252 
rect 15 252 18 255 
rect 15 255 18 258 
rect 15 258 18 261 
rect 15 261 18 264 
rect 15 264 18 267 
rect 15 267 18 270 
rect 15 270 18 273 
rect 15 273 18 276 
rect 15 276 18 279 
rect 15 279 18 282 
rect 15 282 18 285 
rect 15 285 18 288 
rect 15 288 18 291 
rect 15 291 18 294 
rect 15 294 18 297 
rect 15 297 18 300 
rect 15 300 18 303 
rect 15 303 18 306 
rect 15 306 18 309 
rect 15 309 18 312 
rect 15 312 18 315 
rect 15 315 18 318 
rect 15 318 18 321 
rect 15 321 18 324 
rect 15 324 18 327 
rect 15 327 18 330 
rect 15 330 18 333 
rect 15 333 18 336 
rect 15 336 18 339 
rect 15 339 18 342 
rect 15 342 18 345 
rect 15 345 18 348 
rect 15 348 18 351 
rect 15 351 18 354 
rect 15 354 18 357 
rect 15 357 18 360 
rect 15 360 18 363 
rect 15 363 18 366 
rect 15 366 18 369 
rect 15 369 18 372 
rect 15 372 18 375 
rect 15 375 18 378 
rect 15 378 18 381 
rect 15 381 18 384 
rect 15 384 18 387 
rect 15 387 18 390 
rect 15 390 18 393 
rect 15 393 18 396 
rect 15 396 18 399 
rect 15 399 18 402 
rect 15 402 18 405 
rect 15 405 18 408 
rect 15 408 18 411 
rect 15 411 18 414 
rect 15 414 18 417 
rect 15 417 18 420 
rect 15 420 18 423 
rect 15 423 18 426 
rect 15 426 18 429 
rect 15 429 18 432 
rect 15 432 18 435 
rect 15 435 18 438 
rect 15 438 18 441 
rect 15 441 18 444 
rect 15 444 18 447 
rect 15 447 18 450 
rect 15 450 18 453 
rect 15 453 18 456 
rect 15 456 18 459 
rect 15 459 18 462 
rect 15 462 18 465 
rect 15 465 18 468 
rect 15 468 18 471 
rect 15 471 18 474 
rect 15 474 18 477 
rect 15 477 18 480 
rect 15 480 18 483 
rect 15 483 18 486 
rect 15 486 18 489 
rect 15 489 18 492 
rect 15 492 18 495 
rect 15 495 18 498 
rect 15 498 18 501 
rect 15 501 18 504 
rect 15 504 18 507 
rect 15 507 18 510 
rect 18 0 21 3 
rect 18 3 21 6 
rect 18 6 21 9 
rect 18 9 21 12 
rect 18 12 21 15 
rect 18 15 21 18 
rect 18 18 21 21 
rect 18 21 21 24 
rect 18 24 21 27 
rect 18 27 21 30 
rect 18 30 21 33 
rect 18 33 21 36 
rect 18 36 21 39 
rect 18 39 21 42 
rect 18 42 21 45 
rect 18 45 21 48 
rect 18 48 21 51 
rect 18 51 21 54 
rect 18 54 21 57 
rect 18 57 21 60 
rect 18 60 21 63 
rect 18 63 21 66 
rect 18 66 21 69 
rect 18 69 21 72 
rect 18 72 21 75 
rect 18 75 21 78 
rect 18 78 21 81 
rect 18 81 21 84 
rect 18 84 21 87 
rect 18 87 21 90 
rect 18 90 21 93 
rect 18 93 21 96 
rect 18 96 21 99 
rect 18 99 21 102 
rect 18 102 21 105 
rect 18 105 21 108 
rect 18 108 21 111 
rect 18 111 21 114 
rect 18 114 21 117 
rect 18 117 21 120 
rect 18 120 21 123 
rect 18 123 21 126 
rect 18 126 21 129 
rect 18 129 21 132 
rect 18 132 21 135 
rect 18 135 21 138 
rect 18 138 21 141 
rect 18 141 21 144 
rect 18 144 21 147 
rect 18 147 21 150 
rect 18 150 21 153 
rect 18 153 21 156 
rect 18 156 21 159 
rect 18 159 21 162 
rect 18 162 21 165 
rect 18 165 21 168 
rect 18 168 21 171 
rect 18 171 21 174 
rect 18 174 21 177 
rect 18 177 21 180 
rect 18 180 21 183 
rect 18 183 21 186 
rect 18 186 21 189 
rect 18 189 21 192 
rect 18 192 21 195 
rect 18 195 21 198 
rect 18 198 21 201 
rect 18 201 21 204 
rect 18 204 21 207 
rect 18 207 21 210 
rect 18 210 21 213 
rect 18 213 21 216 
rect 18 216 21 219 
rect 18 219 21 222 
rect 18 222 21 225 
rect 18 225 21 228 
rect 18 228 21 231 
rect 18 231 21 234 
rect 18 234 21 237 
rect 18 237 21 240 
rect 18 240 21 243 
rect 18 243 21 246 
rect 18 246 21 249 
rect 18 249 21 252 
rect 18 252 21 255 
rect 18 255 21 258 
rect 18 258 21 261 
rect 18 261 21 264 
rect 18 264 21 267 
rect 18 267 21 270 
rect 18 270 21 273 
rect 18 273 21 276 
rect 18 276 21 279 
rect 18 279 21 282 
rect 18 282 21 285 
rect 18 285 21 288 
rect 18 288 21 291 
rect 18 291 21 294 
rect 18 294 21 297 
rect 18 297 21 300 
rect 18 300 21 303 
rect 18 303 21 306 
rect 18 306 21 309 
rect 18 309 21 312 
rect 18 312 21 315 
rect 18 315 21 318 
rect 18 318 21 321 
rect 18 321 21 324 
rect 18 324 21 327 
rect 18 327 21 330 
rect 18 330 21 333 
rect 18 333 21 336 
rect 18 336 21 339 
rect 18 339 21 342 
rect 18 342 21 345 
rect 18 345 21 348 
rect 18 348 21 351 
rect 18 351 21 354 
rect 18 354 21 357 
rect 18 357 21 360 
rect 18 360 21 363 
rect 18 363 21 366 
rect 18 366 21 369 
rect 18 369 21 372 
rect 18 372 21 375 
rect 18 375 21 378 
rect 18 378 21 381 
rect 18 381 21 384 
rect 18 384 21 387 
rect 18 387 21 390 
rect 18 390 21 393 
rect 18 393 21 396 
rect 18 396 21 399 
rect 18 399 21 402 
rect 18 402 21 405 
rect 18 405 21 408 
rect 18 408 21 411 
rect 18 411 21 414 
rect 18 414 21 417 
rect 18 417 21 420 
rect 18 420 21 423 
rect 18 423 21 426 
rect 18 426 21 429 
rect 18 429 21 432 
rect 18 432 21 435 
rect 18 435 21 438 
rect 18 438 21 441 
rect 18 441 21 444 
rect 18 444 21 447 
rect 18 447 21 450 
rect 18 450 21 453 
rect 18 453 21 456 
rect 18 456 21 459 
rect 18 459 21 462 
rect 18 462 21 465 
rect 18 465 21 468 
rect 18 468 21 471 
rect 18 471 21 474 
rect 18 474 21 477 
rect 18 477 21 480 
rect 18 480 21 483 
rect 18 483 21 486 
rect 18 486 21 489 
rect 18 489 21 492 
rect 18 492 21 495 
rect 18 495 21 498 
rect 18 498 21 501 
rect 18 501 21 504 
rect 18 504 21 507 
rect 18 507 21 510 
rect 21 0 24 3 
rect 21 3 24 6 
rect 21 6 24 9 
rect 21 9 24 12 
rect 21 12 24 15 
rect 21 15 24 18 
rect 21 18 24 21 
rect 21 21 24 24 
rect 21 24 24 27 
rect 21 27 24 30 
rect 21 30 24 33 
rect 21 33 24 36 
rect 21 36 24 39 
rect 21 39 24 42 
rect 21 42 24 45 
rect 21 45 24 48 
rect 21 48 24 51 
rect 21 51 24 54 
rect 21 54 24 57 
rect 21 57 24 60 
rect 21 60 24 63 
rect 21 63 24 66 
rect 21 66 24 69 
rect 21 69 24 72 
rect 21 72 24 75 
rect 21 75 24 78 
rect 21 78 24 81 
rect 21 81 24 84 
rect 21 84 24 87 
rect 21 87 24 90 
rect 21 90 24 93 
rect 21 93 24 96 
rect 21 96 24 99 
rect 21 99 24 102 
rect 21 102 24 105 
rect 21 105 24 108 
rect 21 108 24 111 
rect 21 111 24 114 
rect 21 114 24 117 
rect 21 117 24 120 
rect 21 120 24 123 
rect 21 123 24 126 
rect 21 126 24 129 
rect 21 129 24 132 
rect 21 132 24 135 
rect 21 135 24 138 
rect 21 138 24 141 
rect 21 141 24 144 
rect 21 144 24 147 
rect 21 147 24 150 
rect 21 150 24 153 
rect 21 153 24 156 
rect 21 156 24 159 
rect 21 159 24 162 
rect 21 162 24 165 
rect 21 165 24 168 
rect 21 168 24 171 
rect 21 171 24 174 
rect 21 174 24 177 
rect 21 177 24 180 
rect 21 180 24 183 
rect 21 183 24 186 
rect 21 186 24 189 
rect 21 189 24 192 
rect 21 192 24 195 
rect 21 195 24 198 
rect 21 198 24 201 
rect 21 201 24 204 
rect 21 204 24 207 
rect 21 207 24 210 
rect 21 210 24 213 
rect 21 213 24 216 
rect 21 216 24 219 
rect 21 219 24 222 
rect 21 222 24 225 
rect 21 225 24 228 
rect 21 228 24 231 
rect 21 231 24 234 
rect 21 234 24 237 
rect 21 237 24 240 
rect 21 240 24 243 
rect 21 243 24 246 
rect 21 246 24 249 
rect 21 249 24 252 
rect 21 252 24 255 
rect 21 255 24 258 
rect 21 258 24 261 
rect 21 261 24 264 
rect 21 264 24 267 
rect 21 267 24 270 
rect 21 270 24 273 
rect 21 273 24 276 
rect 21 276 24 279 
rect 21 279 24 282 
rect 21 282 24 285 
rect 21 285 24 288 
rect 21 288 24 291 
rect 21 291 24 294 
rect 21 294 24 297 
rect 21 297 24 300 
rect 21 300 24 303 
rect 21 303 24 306 
rect 21 306 24 309 
rect 21 309 24 312 
rect 21 312 24 315 
rect 21 315 24 318 
rect 21 318 24 321 
rect 21 321 24 324 
rect 21 324 24 327 
rect 21 327 24 330 
rect 21 330 24 333 
rect 21 333 24 336 
rect 21 336 24 339 
rect 21 339 24 342 
rect 21 342 24 345 
rect 21 345 24 348 
rect 21 348 24 351 
rect 21 351 24 354 
rect 21 354 24 357 
rect 21 357 24 360 
rect 21 360 24 363 
rect 21 363 24 366 
rect 21 366 24 369 
rect 21 369 24 372 
rect 21 372 24 375 
rect 21 375 24 378 
rect 21 378 24 381 
rect 21 381 24 384 
rect 21 384 24 387 
rect 21 387 24 390 
rect 21 390 24 393 
rect 21 393 24 396 
rect 21 396 24 399 
rect 21 399 24 402 
rect 21 402 24 405 
rect 21 405 24 408 
rect 21 408 24 411 
rect 21 411 24 414 
rect 21 414 24 417 
rect 21 417 24 420 
rect 21 420 24 423 
rect 21 423 24 426 
rect 21 426 24 429 
rect 21 429 24 432 
rect 21 432 24 435 
rect 21 435 24 438 
rect 21 438 24 441 
rect 21 441 24 444 
rect 21 444 24 447 
rect 21 447 24 450 
rect 21 450 24 453 
rect 21 453 24 456 
rect 21 456 24 459 
rect 21 459 24 462 
rect 21 462 24 465 
rect 21 465 24 468 
rect 21 468 24 471 
rect 21 471 24 474 
rect 21 474 24 477 
rect 21 477 24 480 
rect 21 480 24 483 
rect 21 483 24 486 
rect 21 486 24 489 
rect 21 489 24 492 
rect 21 492 24 495 
rect 21 495 24 498 
rect 21 498 24 501 
rect 21 501 24 504 
rect 21 504 24 507 
rect 21 507 24 510 
rect 24 0 27 3 
rect 24 3 27 6 
rect 24 6 27 9 
rect 24 9 27 12 
rect 24 12 27 15 
rect 24 15 27 18 
rect 24 18 27 21 
rect 24 21 27 24 
rect 24 24 27 27 
rect 24 27 27 30 
rect 24 30 27 33 
rect 24 33 27 36 
rect 24 36 27 39 
rect 24 39 27 42 
rect 24 42 27 45 
rect 24 45 27 48 
rect 24 48 27 51 
rect 24 51 27 54 
rect 24 54 27 57 
rect 24 57 27 60 
rect 24 60 27 63 
rect 24 63 27 66 
rect 24 66 27 69 
rect 24 69 27 72 
rect 24 72 27 75 
rect 24 75 27 78 
rect 24 78 27 81 
rect 24 81 27 84 
rect 24 84 27 87 
rect 24 87 27 90 
rect 24 90 27 93 
rect 24 93 27 96 
rect 24 96 27 99 
rect 24 99 27 102 
rect 24 102 27 105 
rect 24 105 27 108 
rect 24 108 27 111 
rect 24 111 27 114 
rect 24 114 27 117 
rect 24 117 27 120 
rect 24 120 27 123 
rect 24 123 27 126 
rect 24 126 27 129 
rect 24 129 27 132 
rect 24 132 27 135 
rect 24 135 27 138 
rect 24 138 27 141 
rect 24 141 27 144 
rect 24 144 27 147 
rect 24 147 27 150 
rect 24 150 27 153 
rect 24 153 27 156 
rect 24 156 27 159 
rect 24 159 27 162 
rect 24 162 27 165 
rect 24 165 27 168 
rect 24 168 27 171 
rect 24 171 27 174 
rect 24 174 27 177 
rect 24 177 27 180 
rect 24 180 27 183 
rect 24 183 27 186 
rect 24 186 27 189 
rect 24 189 27 192 
rect 24 192 27 195 
rect 24 195 27 198 
rect 24 198 27 201 
rect 24 201 27 204 
rect 24 204 27 207 
rect 24 207 27 210 
rect 24 210 27 213 
rect 24 213 27 216 
rect 24 216 27 219 
rect 24 219 27 222 
rect 24 222 27 225 
rect 24 225 27 228 
rect 24 228 27 231 
rect 24 231 27 234 
rect 24 234 27 237 
rect 24 237 27 240 
rect 24 240 27 243 
rect 24 243 27 246 
rect 24 246 27 249 
rect 24 249 27 252 
rect 24 252 27 255 
rect 24 255 27 258 
rect 24 258 27 261 
rect 24 261 27 264 
rect 24 264 27 267 
rect 24 267 27 270 
rect 24 270 27 273 
rect 24 273 27 276 
rect 24 276 27 279 
rect 24 279 27 282 
rect 24 282 27 285 
rect 24 285 27 288 
rect 24 288 27 291 
rect 24 291 27 294 
rect 24 294 27 297 
rect 24 297 27 300 
rect 24 300 27 303 
rect 24 303 27 306 
rect 24 306 27 309 
rect 24 309 27 312 
rect 24 312 27 315 
rect 24 315 27 318 
rect 24 318 27 321 
rect 24 321 27 324 
rect 24 324 27 327 
rect 24 327 27 330 
rect 24 330 27 333 
rect 24 333 27 336 
rect 24 336 27 339 
rect 24 339 27 342 
rect 24 342 27 345 
rect 24 345 27 348 
rect 24 348 27 351 
rect 24 351 27 354 
rect 24 354 27 357 
rect 24 357 27 360 
rect 24 360 27 363 
rect 24 363 27 366 
rect 24 366 27 369 
rect 24 369 27 372 
rect 24 372 27 375 
rect 24 375 27 378 
rect 24 378 27 381 
rect 24 381 27 384 
rect 24 384 27 387 
rect 24 387 27 390 
rect 24 390 27 393 
rect 24 393 27 396 
rect 24 396 27 399 
rect 24 399 27 402 
rect 24 402 27 405 
rect 24 405 27 408 
rect 24 408 27 411 
rect 24 411 27 414 
rect 24 414 27 417 
rect 24 417 27 420 
rect 24 420 27 423 
rect 24 423 27 426 
rect 24 426 27 429 
rect 24 429 27 432 
rect 24 432 27 435 
rect 24 435 27 438 
rect 24 438 27 441 
rect 24 441 27 444 
rect 24 444 27 447 
rect 24 447 27 450 
rect 24 450 27 453 
rect 24 453 27 456 
rect 24 456 27 459 
rect 24 459 27 462 
rect 24 462 27 465 
rect 24 465 27 468 
rect 24 468 27 471 
rect 24 471 27 474 
rect 24 474 27 477 
rect 24 477 27 480 
rect 24 480 27 483 
rect 24 483 27 486 
rect 24 486 27 489 
rect 24 489 27 492 
rect 24 492 27 495 
rect 24 495 27 498 
rect 24 498 27 501 
rect 24 501 27 504 
rect 24 504 27 507 
rect 24 507 27 510 
rect 27 0 30 3 
rect 27 3 30 6 
rect 27 6 30 9 
rect 27 9 30 12 
rect 27 12 30 15 
rect 27 15 30 18 
rect 27 18 30 21 
rect 27 21 30 24 
rect 27 24 30 27 
rect 27 27 30 30 
rect 27 30 30 33 
rect 27 33 30 36 
rect 27 36 30 39 
rect 27 39 30 42 
rect 27 42 30 45 
rect 27 45 30 48 
rect 27 48 30 51 
rect 27 51 30 54 
rect 27 54 30 57 
rect 27 57 30 60 
rect 27 60 30 63 
rect 27 63 30 66 
rect 27 66 30 69 
rect 27 69 30 72 
rect 27 72 30 75 
rect 27 75 30 78 
rect 27 78 30 81 
rect 27 81 30 84 
rect 27 84 30 87 
rect 27 87 30 90 
rect 27 90 30 93 
rect 27 93 30 96 
rect 27 96 30 99 
rect 27 99 30 102 
rect 27 102 30 105 
rect 27 105 30 108 
rect 27 108 30 111 
rect 27 111 30 114 
rect 27 114 30 117 
rect 27 117 30 120 
rect 27 120 30 123 
rect 27 123 30 126 
rect 27 126 30 129 
rect 27 129 30 132 
rect 27 132 30 135 
rect 27 135 30 138 
rect 27 138 30 141 
rect 27 141 30 144 
rect 27 144 30 147 
rect 27 147 30 150 
rect 27 150 30 153 
rect 27 153 30 156 
rect 27 156 30 159 
rect 27 159 30 162 
rect 27 162 30 165 
rect 27 165 30 168 
rect 27 168 30 171 
rect 27 171 30 174 
rect 27 174 30 177 
rect 27 177 30 180 
rect 27 180 30 183 
rect 27 183 30 186 
rect 27 186 30 189 
rect 27 189 30 192 
rect 27 192 30 195 
rect 27 195 30 198 
rect 27 198 30 201 
rect 27 201 30 204 
rect 27 204 30 207 
rect 27 207 30 210 
rect 27 210 30 213 
rect 27 213 30 216 
rect 27 216 30 219 
rect 27 219 30 222 
rect 27 222 30 225 
rect 27 225 30 228 
rect 27 228 30 231 
rect 27 231 30 234 
rect 27 234 30 237 
rect 27 237 30 240 
rect 27 240 30 243 
rect 27 243 30 246 
rect 27 246 30 249 
rect 27 249 30 252 
rect 27 252 30 255 
rect 27 255 30 258 
rect 27 258 30 261 
rect 27 261 30 264 
rect 27 264 30 267 
rect 27 267 30 270 
rect 27 270 30 273 
rect 27 273 30 276 
rect 27 276 30 279 
rect 27 279 30 282 
rect 27 282 30 285 
rect 27 285 30 288 
rect 27 288 30 291 
rect 27 291 30 294 
rect 27 294 30 297 
rect 27 297 30 300 
rect 27 300 30 303 
rect 27 303 30 306 
rect 27 306 30 309 
rect 27 309 30 312 
rect 27 312 30 315 
rect 27 315 30 318 
rect 27 318 30 321 
rect 27 321 30 324 
rect 27 324 30 327 
rect 27 327 30 330 
rect 27 330 30 333 
rect 27 333 30 336 
rect 27 336 30 339 
rect 27 339 30 342 
rect 27 342 30 345 
rect 27 345 30 348 
rect 27 348 30 351 
rect 27 351 30 354 
rect 27 354 30 357 
rect 27 357 30 360 
rect 27 360 30 363 
rect 27 363 30 366 
rect 27 366 30 369 
rect 27 369 30 372 
rect 27 372 30 375 
rect 27 375 30 378 
rect 27 378 30 381 
rect 27 381 30 384 
rect 27 384 30 387 
rect 27 387 30 390 
rect 27 390 30 393 
rect 27 393 30 396 
rect 27 396 30 399 
rect 27 399 30 402 
rect 27 402 30 405 
rect 27 405 30 408 
rect 27 408 30 411 
rect 27 411 30 414 
rect 27 414 30 417 
rect 27 417 30 420 
rect 27 420 30 423 
rect 27 423 30 426 
rect 27 426 30 429 
rect 27 429 30 432 
rect 27 432 30 435 
rect 27 435 30 438 
rect 27 438 30 441 
rect 27 441 30 444 
rect 27 444 30 447 
rect 27 447 30 450 
rect 27 450 30 453 
rect 27 453 30 456 
rect 27 456 30 459 
rect 27 459 30 462 
rect 27 462 30 465 
rect 27 465 30 468 
rect 27 468 30 471 
rect 27 471 30 474 
rect 27 474 30 477 
rect 27 477 30 480 
rect 27 480 30 483 
rect 27 483 30 486 
rect 27 486 30 489 
rect 27 489 30 492 
rect 27 492 30 495 
rect 27 495 30 498 
rect 27 498 30 501 
rect 27 501 30 504 
rect 27 504 30 507 
rect 27 507 30 510 
rect 30 0 33 3 
rect 30 3 33 6 
rect 30 6 33 9 
rect 30 9 33 12 
rect 30 12 33 15 
rect 30 15 33 18 
rect 30 18 33 21 
rect 30 21 33 24 
rect 30 24 33 27 
rect 30 27 33 30 
rect 30 30 33 33 
rect 30 33 33 36 
rect 30 36 33 39 
rect 30 39 33 42 
rect 30 42 33 45 
rect 30 45 33 48 
rect 30 48 33 51 
rect 30 51 33 54 
rect 30 54 33 57 
rect 30 57 33 60 
rect 30 60 33 63 
rect 30 63 33 66 
rect 30 66 33 69 
rect 30 69 33 72 
rect 30 72 33 75 
rect 30 75 33 78 
rect 30 78 33 81 
rect 30 81 33 84 
rect 30 84 33 87 
rect 30 87 33 90 
rect 30 90 33 93 
rect 30 93 33 96 
rect 30 96 33 99 
rect 30 99 33 102 
rect 30 102 33 105 
rect 30 105 33 108 
rect 30 108 33 111 
rect 30 111 33 114 
rect 30 114 33 117 
rect 30 117 33 120 
rect 30 120 33 123 
rect 30 123 33 126 
rect 30 126 33 129 
rect 30 129 33 132 
rect 30 132 33 135 
rect 30 135 33 138 
rect 30 138 33 141 
rect 30 141 33 144 
rect 30 144 33 147 
rect 30 147 33 150 
rect 30 150 33 153 
rect 30 153 33 156 
rect 30 156 33 159 
rect 30 159 33 162 
rect 30 162 33 165 
rect 30 165 33 168 
rect 30 168 33 171 
rect 30 171 33 174 
rect 30 174 33 177 
rect 30 177 33 180 
rect 30 180 33 183 
rect 30 183 33 186 
rect 30 186 33 189 
rect 30 189 33 192 
rect 30 192 33 195 
rect 30 195 33 198 
rect 30 198 33 201 
rect 30 201 33 204 
rect 30 204 33 207 
rect 30 207 33 210 
rect 30 210 33 213 
rect 30 213 33 216 
rect 30 216 33 219 
rect 30 219 33 222 
rect 30 222 33 225 
rect 30 225 33 228 
rect 30 228 33 231 
rect 30 231 33 234 
rect 30 234 33 237 
rect 30 237 33 240 
rect 30 240 33 243 
rect 30 243 33 246 
rect 30 246 33 249 
rect 30 249 33 252 
rect 30 252 33 255 
rect 30 255 33 258 
rect 30 258 33 261 
rect 30 261 33 264 
rect 30 264 33 267 
rect 30 267 33 270 
rect 30 270 33 273 
rect 30 273 33 276 
rect 30 276 33 279 
rect 30 279 33 282 
rect 30 282 33 285 
rect 30 285 33 288 
rect 30 288 33 291 
rect 30 291 33 294 
rect 30 294 33 297 
rect 30 297 33 300 
rect 30 300 33 303 
rect 30 303 33 306 
rect 30 306 33 309 
rect 30 309 33 312 
rect 30 312 33 315 
rect 30 315 33 318 
rect 30 318 33 321 
rect 30 321 33 324 
rect 30 324 33 327 
rect 30 327 33 330 
rect 30 330 33 333 
rect 30 333 33 336 
rect 30 336 33 339 
rect 30 339 33 342 
rect 30 342 33 345 
rect 30 345 33 348 
rect 30 348 33 351 
rect 30 351 33 354 
rect 30 354 33 357 
rect 30 357 33 360 
rect 30 360 33 363 
rect 30 363 33 366 
rect 30 366 33 369 
rect 30 369 33 372 
rect 30 372 33 375 
rect 30 375 33 378 
rect 30 378 33 381 
rect 30 381 33 384 
rect 30 384 33 387 
rect 30 387 33 390 
rect 30 390 33 393 
rect 30 393 33 396 
rect 30 396 33 399 
rect 30 399 33 402 
rect 30 402 33 405 
rect 30 405 33 408 
rect 30 408 33 411 
rect 30 411 33 414 
rect 30 414 33 417 
rect 30 417 33 420 
rect 30 420 33 423 
rect 30 423 33 426 
rect 30 426 33 429 
rect 30 429 33 432 
rect 30 432 33 435 
rect 30 435 33 438 
rect 30 438 33 441 
rect 30 441 33 444 
rect 30 444 33 447 
rect 30 447 33 450 
rect 30 450 33 453 
rect 30 453 33 456 
rect 30 456 33 459 
rect 30 459 33 462 
rect 30 462 33 465 
rect 30 465 33 468 
rect 30 468 33 471 
rect 30 471 33 474 
rect 30 474 33 477 
rect 30 477 33 480 
rect 30 480 33 483 
rect 30 483 33 486 
rect 30 486 33 489 
rect 30 489 33 492 
rect 30 492 33 495 
rect 30 495 33 498 
rect 30 498 33 501 
rect 30 501 33 504 
rect 30 504 33 507 
rect 30 507 33 510 
rect 33 0 36 3 
rect 33 3 36 6 
rect 33 6 36 9 
rect 33 9 36 12 
rect 33 12 36 15 
rect 33 15 36 18 
rect 33 18 36 21 
rect 33 21 36 24 
rect 33 24 36 27 
rect 33 27 36 30 
rect 33 30 36 33 
rect 33 33 36 36 
rect 33 36 36 39 
rect 33 39 36 42 
rect 33 42 36 45 
rect 33 45 36 48 
rect 33 48 36 51 
rect 33 51 36 54 
rect 33 54 36 57 
rect 33 57 36 60 
rect 33 60 36 63 
rect 33 63 36 66 
rect 33 66 36 69 
rect 33 69 36 72 
rect 33 72 36 75 
rect 33 75 36 78 
rect 33 78 36 81 
rect 33 81 36 84 
rect 33 84 36 87 
rect 33 87 36 90 
rect 33 90 36 93 
rect 33 93 36 96 
rect 33 96 36 99 
rect 33 99 36 102 
rect 33 102 36 105 
rect 33 105 36 108 
rect 33 108 36 111 
rect 33 111 36 114 
rect 33 114 36 117 
rect 33 117 36 120 
rect 33 120 36 123 
rect 33 123 36 126 
rect 33 126 36 129 
rect 33 129 36 132 
rect 33 132 36 135 
rect 33 135 36 138 
rect 33 138 36 141 
rect 33 141 36 144 
rect 33 144 36 147 
rect 33 147 36 150 
rect 33 150 36 153 
rect 33 153 36 156 
rect 33 156 36 159 
rect 33 159 36 162 
rect 33 162 36 165 
rect 33 165 36 168 
rect 33 168 36 171 
rect 33 171 36 174 
rect 33 174 36 177 
rect 33 177 36 180 
rect 33 180 36 183 
rect 33 183 36 186 
rect 33 186 36 189 
rect 33 189 36 192 
rect 33 192 36 195 
rect 33 195 36 198 
rect 33 198 36 201 
rect 33 201 36 204 
rect 33 204 36 207 
rect 33 207 36 210 
rect 33 210 36 213 
rect 33 213 36 216 
rect 33 216 36 219 
rect 33 219 36 222 
rect 33 222 36 225 
rect 33 225 36 228 
rect 33 228 36 231 
rect 33 231 36 234 
rect 33 234 36 237 
rect 33 237 36 240 
rect 33 240 36 243 
rect 33 243 36 246 
rect 33 246 36 249 
rect 33 249 36 252 
rect 33 252 36 255 
rect 33 255 36 258 
rect 33 258 36 261 
rect 33 261 36 264 
rect 33 264 36 267 
rect 33 267 36 270 
rect 33 270 36 273 
rect 33 273 36 276 
rect 33 276 36 279 
rect 33 279 36 282 
rect 33 282 36 285 
rect 33 285 36 288 
rect 33 288 36 291 
rect 33 291 36 294 
rect 33 294 36 297 
rect 33 297 36 300 
rect 33 300 36 303 
rect 33 303 36 306 
rect 33 306 36 309 
rect 33 309 36 312 
rect 33 312 36 315 
rect 33 315 36 318 
rect 33 318 36 321 
rect 33 321 36 324 
rect 33 324 36 327 
rect 33 327 36 330 
rect 33 330 36 333 
rect 33 333 36 336 
rect 33 336 36 339 
rect 33 339 36 342 
rect 33 342 36 345 
rect 33 345 36 348 
rect 33 348 36 351 
rect 33 351 36 354 
rect 33 354 36 357 
rect 33 357 36 360 
rect 33 360 36 363 
rect 33 363 36 366 
rect 33 366 36 369 
rect 33 369 36 372 
rect 33 372 36 375 
rect 33 375 36 378 
rect 33 378 36 381 
rect 33 381 36 384 
rect 33 384 36 387 
rect 33 387 36 390 
rect 33 390 36 393 
rect 33 393 36 396 
rect 33 396 36 399 
rect 33 399 36 402 
rect 33 402 36 405 
rect 33 405 36 408 
rect 33 408 36 411 
rect 33 411 36 414 
rect 33 414 36 417 
rect 33 417 36 420 
rect 33 420 36 423 
rect 33 423 36 426 
rect 33 426 36 429 
rect 33 429 36 432 
rect 33 432 36 435 
rect 33 435 36 438 
rect 33 438 36 441 
rect 33 441 36 444 
rect 33 444 36 447 
rect 33 447 36 450 
rect 33 450 36 453 
rect 33 453 36 456 
rect 33 456 36 459 
rect 33 459 36 462 
rect 33 462 36 465 
rect 33 465 36 468 
rect 33 468 36 471 
rect 33 471 36 474 
rect 33 474 36 477 
rect 33 477 36 480 
rect 33 480 36 483 
rect 33 483 36 486 
rect 33 486 36 489 
rect 33 489 36 492 
rect 33 492 36 495 
rect 33 495 36 498 
rect 33 498 36 501 
rect 33 501 36 504 
rect 33 504 36 507 
rect 33 507 36 510 
rect 36 0 39 3 
rect 36 3 39 6 
rect 36 6 39 9 
rect 36 9 39 12 
rect 36 12 39 15 
rect 36 15 39 18 
rect 36 18 39 21 
rect 36 21 39 24 
rect 36 24 39 27 
rect 36 27 39 30 
rect 36 30 39 33 
rect 36 33 39 36 
rect 36 36 39 39 
rect 36 39 39 42 
rect 36 42 39 45 
rect 36 45 39 48 
rect 36 48 39 51 
rect 36 51 39 54 
rect 36 54 39 57 
rect 36 57 39 60 
rect 36 60 39 63 
rect 36 63 39 66 
rect 36 66 39 69 
rect 36 69 39 72 
rect 36 72 39 75 
rect 36 75 39 78 
rect 36 78 39 81 
rect 36 81 39 84 
rect 36 84 39 87 
rect 36 87 39 90 
rect 36 90 39 93 
rect 36 93 39 96 
rect 36 96 39 99 
rect 36 99 39 102 
rect 36 102 39 105 
rect 36 105 39 108 
rect 36 108 39 111 
rect 36 111 39 114 
rect 36 114 39 117 
rect 36 117 39 120 
rect 36 120 39 123 
rect 36 123 39 126 
rect 36 126 39 129 
rect 36 129 39 132 
rect 36 132 39 135 
rect 36 135 39 138 
rect 36 138 39 141 
rect 36 141 39 144 
rect 36 144 39 147 
rect 36 147 39 150 
rect 36 150 39 153 
rect 36 153 39 156 
rect 36 156 39 159 
rect 36 159 39 162 
rect 36 162 39 165 
rect 36 165 39 168 
rect 36 168 39 171 
rect 36 171 39 174 
rect 36 174 39 177 
rect 36 177 39 180 
rect 36 180 39 183 
rect 36 183 39 186 
rect 36 186 39 189 
rect 36 189 39 192 
rect 36 192 39 195 
rect 36 195 39 198 
rect 36 198 39 201 
rect 36 201 39 204 
rect 36 204 39 207 
rect 36 207 39 210 
rect 36 210 39 213 
rect 36 213 39 216 
rect 36 216 39 219 
rect 36 219 39 222 
rect 36 222 39 225 
rect 36 225 39 228 
rect 36 228 39 231 
rect 36 231 39 234 
rect 36 234 39 237 
rect 36 237 39 240 
rect 36 240 39 243 
rect 36 243 39 246 
rect 36 246 39 249 
rect 36 249 39 252 
rect 36 252 39 255 
rect 36 255 39 258 
rect 36 258 39 261 
rect 36 261 39 264 
rect 36 264 39 267 
rect 36 267 39 270 
rect 36 270 39 273 
rect 36 273 39 276 
rect 36 276 39 279 
rect 36 279 39 282 
rect 36 282 39 285 
rect 36 285 39 288 
rect 36 288 39 291 
rect 36 291 39 294 
rect 36 294 39 297 
rect 36 297 39 300 
rect 36 300 39 303 
rect 36 303 39 306 
rect 36 306 39 309 
rect 36 309 39 312 
rect 36 312 39 315 
rect 36 315 39 318 
rect 36 318 39 321 
rect 36 321 39 324 
rect 36 324 39 327 
rect 36 327 39 330 
rect 36 330 39 333 
rect 36 333 39 336 
rect 36 336 39 339 
rect 36 339 39 342 
rect 36 342 39 345 
rect 36 345 39 348 
rect 36 348 39 351 
rect 36 351 39 354 
rect 36 354 39 357 
rect 36 357 39 360 
rect 36 360 39 363 
rect 36 363 39 366 
rect 36 366 39 369 
rect 36 369 39 372 
rect 36 372 39 375 
rect 36 375 39 378 
rect 36 378 39 381 
rect 36 381 39 384 
rect 36 384 39 387 
rect 36 387 39 390 
rect 36 390 39 393 
rect 36 393 39 396 
rect 36 396 39 399 
rect 36 399 39 402 
rect 36 402 39 405 
rect 36 405 39 408 
rect 36 408 39 411 
rect 36 411 39 414 
rect 36 414 39 417 
rect 36 417 39 420 
rect 36 420 39 423 
rect 36 423 39 426 
rect 36 426 39 429 
rect 36 429 39 432 
rect 36 432 39 435 
rect 36 435 39 438 
rect 36 438 39 441 
rect 36 441 39 444 
rect 36 444 39 447 
rect 36 447 39 450 
rect 36 450 39 453 
rect 36 453 39 456 
rect 36 456 39 459 
rect 36 459 39 462 
rect 36 462 39 465 
rect 36 465 39 468 
rect 36 468 39 471 
rect 36 471 39 474 
rect 36 474 39 477 
rect 36 477 39 480 
rect 36 480 39 483 
rect 36 483 39 486 
rect 36 486 39 489 
rect 36 489 39 492 
rect 36 492 39 495 
rect 36 495 39 498 
rect 36 498 39 501 
rect 36 501 39 504 
rect 36 504 39 507 
rect 36 507 39 510 
rect 39 0 42 3 
rect 39 3 42 6 
rect 39 6 42 9 
rect 39 9 42 12 
rect 39 12 42 15 
rect 39 15 42 18 
rect 39 18 42 21 
rect 39 21 42 24 
rect 39 24 42 27 
rect 39 27 42 30 
rect 39 30 42 33 
rect 39 33 42 36 
rect 39 36 42 39 
rect 39 39 42 42 
rect 39 42 42 45 
rect 39 45 42 48 
rect 39 48 42 51 
rect 39 51 42 54 
rect 39 54 42 57 
rect 39 57 42 60 
rect 39 60 42 63 
rect 39 63 42 66 
rect 39 66 42 69 
rect 39 69 42 72 
rect 39 72 42 75 
rect 39 75 42 78 
rect 39 78 42 81 
rect 39 81 42 84 
rect 39 84 42 87 
rect 39 87 42 90 
rect 39 90 42 93 
rect 39 93 42 96 
rect 39 96 42 99 
rect 39 99 42 102 
rect 39 102 42 105 
rect 39 105 42 108 
rect 39 108 42 111 
rect 39 111 42 114 
rect 39 114 42 117 
rect 39 117 42 120 
rect 39 120 42 123 
rect 39 123 42 126 
rect 39 126 42 129 
rect 39 129 42 132 
rect 39 132 42 135 
rect 39 135 42 138 
rect 39 138 42 141 
rect 39 141 42 144 
rect 39 144 42 147 
rect 39 147 42 150 
rect 39 150 42 153 
rect 39 153 42 156 
rect 39 156 42 159 
rect 39 159 42 162 
rect 39 162 42 165 
rect 39 165 42 168 
rect 39 168 42 171 
rect 39 171 42 174 
rect 39 174 42 177 
rect 39 177 42 180 
rect 39 180 42 183 
rect 39 183 42 186 
rect 39 186 42 189 
rect 39 189 42 192 
rect 39 192 42 195 
rect 39 195 42 198 
rect 39 198 42 201 
rect 39 201 42 204 
rect 39 204 42 207 
rect 39 207 42 210 
rect 39 210 42 213 
rect 39 213 42 216 
rect 39 216 42 219 
rect 39 219 42 222 
rect 39 222 42 225 
rect 39 225 42 228 
rect 39 228 42 231 
rect 39 231 42 234 
rect 39 234 42 237 
rect 39 237 42 240 
rect 39 240 42 243 
rect 39 243 42 246 
rect 39 246 42 249 
rect 39 249 42 252 
rect 39 252 42 255 
rect 39 255 42 258 
rect 39 258 42 261 
rect 39 261 42 264 
rect 39 264 42 267 
rect 39 267 42 270 
rect 39 270 42 273 
rect 39 273 42 276 
rect 39 276 42 279 
rect 39 279 42 282 
rect 39 282 42 285 
rect 39 285 42 288 
rect 39 288 42 291 
rect 39 291 42 294 
rect 39 294 42 297 
rect 39 297 42 300 
rect 39 300 42 303 
rect 39 303 42 306 
rect 39 306 42 309 
rect 39 309 42 312 
rect 39 312 42 315 
rect 39 315 42 318 
rect 39 318 42 321 
rect 39 321 42 324 
rect 39 324 42 327 
rect 39 327 42 330 
rect 39 330 42 333 
rect 39 333 42 336 
rect 39 336 42 339 
rect 39 339 42 342 
rect 39 342 42 345 
rect 39 345 42 348 
rect 39 348 42 351 
rect 39 351 42 354 
rect 39 354 42 357 
rect 39 357 42 360 
rect 39 360 42 363 
rect 39 363 42 366 
rect 39 366 42 369 
rect 39 369 42 372 
rect 39 372 42 375 
rect 39 375 42 378 
rect 39 378 42 381 
rect 39 381 42 384 
rect 39 384 42 387 
rect 39 387 42 390 
rect 39 390 42 393 
rect 39 393 42 396 
rect 39 396 42 399 
rect 39 399 42 402 
rect 39 402 42 405 
rect 39 405 42 408 
rect 39 408 42 411 
rect 39 411 42 414 
rect 39 414 42 417 
rect 39 417 42 420 
rect 39 420 42 423 
rect 39 423 42 426 
rect 39 426 42 429 
rect 39 429 42 432 
rect 39 432 42 435 
rect 39 435 42 438 
rect 39 438 42 441 
rect 39 441 42 444 
rect 39 444 42 447 
rect 39 447 42 450 
rect 39 450 42 453 
rect 39 453 42 456 
rect 39 456 42 459 
rect 39 459 42 462 
rect 39 462 42 465 
rect 39 465 42 468 
rect 39 468 42 471 
rect 39 471 42 474 
rect 39 474 42 477 
rect 39 477 42 480 
rect 39 480 42 483 
rect 39 483 42 486 
rect 39 486 42 489 
rect 39 489 42 492 
rect 39 492 42 495 
rect 39 495 42 498 
rect 39 498 42 501 
rect 39 501 42 504 
rect 39 504 42 507 
rect 39 507 42 510 
rect 42 0 45 3 
rect 42 3 45 6 
rect 42 6 45 9 
rect 42 9 45 12 
rect 42 12 45 15 
rect 42 15 45 18 
rect 42 18 45 21 
rect 42 21 45 24 
rect 42 24 45 27 
rect 42 27 45 30 
rect 42 30 45 33 
rect 42 33 45 36 
rect 42 36 45 39 
rect 42 39 45 42 
rect 42 42 45 45 
rect 42 45 45 48 
rect 42 48 45 51 
rect 42 51 45 54 
rect 42 54 45 57 
rect 42 57 45 60 
rect 42 60 45 63 
rect 42 63 45 66 
rect 42 66 45 69 
rect 42 69 45 72 
rect 42 72 45 75 
rect 42 75 45 78 
rect 42 78 45 81 
rect 42 81 45 84 
rect 42 84 45 87 
rect 42 87 45 90 
rect 42 90 45 93 
rect 42 93 45 96 
rect 42 96 45 99 
rect 42 99 45 102 
rect 42 102 45 105 
rect 42 105 45 108 
rect 42 108 45 111 
rect 42 111 45 114 
rect 42 114 45 117 
rect 42 117 45 120 
rect 42 120 45 123 
rect 42 123 45 126 
rect 42 126 45 129 
rect 42 129 45 132 
rect 42 132 45 135 
rect 42 135 45 138 
rect 42 138 45 141 
rect 42 141 45 144 
rect 42 144 45 147 
rect 42 147 45 150 
rect 42 150 45 153 
rect 42 153 45 156 
rect 42 156 45 159 
rect 42 159 45 162 
rect 42 162 45 165 
rect 42 165 45 168 
rect 42 168 45 171 
rect 42 171 45 174 
rect 42 174 45 177 
rect 42 177 45 180 
rect 42 180 45 183 
rect 42 183 45 186 
rect 42 186 45 189 
rect 42 189 45 192 
rect 42 192 45 195 
rect 42 195 45 198 
rect 42 198 45 201 
rect 42 201 45 204 
rect 42 204 45 207 
rect 42 207 45 210 
rect 42 210 45 213 
rect 42 213 45 216 
rect 42 216 45 219 
rect 42 219 45 222 
rect 42 222 45 225 
rect 42 225 45 228 
rect 42 228 45 231 
rect 42 231 45 234 
rect 42 234 45 237 
rect 42 237 45 240 
rect 42 240 45 243 
rect 42 243 45 246 
rect 42 246 45 249 
rect 42 249 45 252 
rect 42 252 45 255 
rect 42 255 45 258 
rect 42 258 45 261 
rect 42 261 45 264 
rect 42 264 45 267 
rect 42 267 45 270 
rect 42 270 45 273 
rect 42 273 45 276 
rect 42 276 45 279 
rect 42 279 45 282 
rect 42 282 45 285 
rect 42 285 45 288 
rect 42 288 45 291 
rect 42 291 45 294 
rect 42 294 45 297 
rect 42 297 45 300 
rect 42 300 45 303 
rect 42 303 45 306 
rect 42 306 45 309 
rect 42 309 45 312 
rect 42 312 45 315 
rect 42 315 45 318 
rect 42 318 45 321 
rect 42 321 45 324 
rect 42 324 45 327 
rect 42 327 45 330 
rect 42 330 45 333 
rect 42 333 45 336 
rect 42 336 45 339 
rect 42 339 45 342 
rect 42 342 45 345 
rect 42 345 45 348 
rect 42 348 45 351 
rect 42 351 45 354 
rect 42 354 45 357 
rect 42 357 45 360 
rect 42 360 45 363 
rect 42 363 45 366 
rect 42 366 45 369 
rect 42 369 45 372 
rect 42 372 45 375 
rect 42 375 45 378 
rect 42 378 45 381 
rect 42 381 45 384 
rect 42 384 45 387 
rect 42 387 45 390 
rect 42 390 45 393 
rect 42 393 45 396 
rect 42 396 45 399 
rect 42 399 45 402 
rect 42 402 45 405 
rect 42 405 45 408 
rect 42 408 45 411 
rect 42 411 45 414 
rect 42 414 45 417 
rect 42 417 45 420 
rect 42 420 45 423 
rect 42 423 45 426 
rect 42 426 45 429 
rect 42 429 45 432 
rect 42 432 45 435 
rect 42 435 45 438 
rect 42 438 45 441 
rect 42 441 45 444 
rect 42 444 45 447 
rect 42 447 45 450 
rect 42 450 45 453 
rect 42 453 45 456 
rect 42 456 45 459 
rect 42 459 45 462 
rect 42 462 45 465 
rect 42 465 45 468 
rect 42 468 45 471 
rect 42 471 45 474 
rect 42 474 45 477 
rect 42 477 45 480 
rect 42 480 45 483 
rect 42 483 45 486 
rect 42 486 45 489 
rect 42 489 45 492 
rect 42 492 45 495 
rect 42 495 45 498 
rect 42 498 45 501 
rect 42 501 45 504 
rect 42 504 45 507 
rect 42 507 45 510 
rect 45 0 48 3 
rect 45 3 48 6 
rect 45 6 48 9 
rect 45 9 48 12 
rect 45 12 48 15 
rect 45 15 48 18 
rect 45 18 48 21 
rect 45 21 48 24 
rect 45 24 48 27 
rect 45 27 48 30 
rect 45 30 48 33 
rect 45 33 48 36 
rect 45 36 48 39 
rect 45 39 48 42 
rect 45 42 48 45 
rect 45 45 48 48 
rect 45 48 48 51 
rect 45 51 48 54 
rect 45 54 48 57 
rect 45 57 48 60 
rect 45 60 48 63 
rect 45 63 48 66 
rect 45 66 48 69 
rect 45 69 48 72 
rect 45 72 48 75 
rect 45 75 48 78 
rect 45 78 48 81 
rect 45 81 48 84 
rect 45 84 48 87 
rect 45 87 48 90 
rect 45 90 48 93 
rect 45 93 48 96 
rect 45 96 48 99 
rect 45 99 48 102 
rect 45 102 48 105 
rect 45 105 48 108 
rect 45 108 48 111 
rect 45 111 48 114 
rect 45 114 48 117 
rect 45 117 48 120 
rect 45 120 48 123 
rect 45 123 48 126 
rect 45 126 48 129 
rect 45 129 48 132 
rect 45 132 48 135 
rect 45 135 48 138 
rect 45 138 48 141 
rect 45 141 48 144 
rect 45 144 48 147 
rect 45 147 48 150 
rect 45 150 48 153 
rect 45 153 48 156 
rect 45 156 48 159 
rect 45 159 48 162 
rect 45 162 48 165 
rect 45 165 48 168 
rect 45 168 48 171 
rect 45 171 48 174 
rect 45 174 48 177 
rect 45 177 48 180 
rect 45 180 48 183 
rect 45 183 48 186 
rect 45 186 48 189 
rect 45 189 48 192 
rect 45 192 48 195 
rect 45 195 48 198 
rect 45 198 48 201 
rect 45 201 48 204 
rect 45 204 48 207 
rect 45 207 48 210 
rect 45 210 48 213 
rect 45 213 48 216 
rect 45 216 48 219 
rect 45 219 48 222 
rect 45 222 48 225 
rect 45 225 48 228 
rect 45 228 48 231 
rect 45 231 48 234 
rect 45 234 48 237 
rect 45 237 48 240 
rect 45 240 48 243 
rect 45 243 48 246 
rect 45 246 48 249 
rect 45 249 48 252 
rect 45 252 48 255 
rect 45 255 48 258 
rect 45 258 48 261 
rect 45 261 48 264 
rect 45 264 48 267 
rect 45 267 48 270 
rect 45 270 48 273 
rect 45 273 48 276 
rect 45 276 48 279 
rect 45 279 48 282 
rect 45 282 48 285 
rect 45 285 48 288 
rect 45 288 48 291 
rect 45 291 48 294 
rect 45 294 48 297 
rect 45 297 48 300 
rect 45 300 48 303 
rect 45 303 48 306 
rect 45 306 48 309 
rect 45 309 48 312 
rect 45 312 48 315 
rect 45 315 48 318 
rect 45 318 48 321 
rect 45 321 48 324 
rect 45 324 48 327 
rect 45 327 48 330 
rect 45 330 48 333 
rect 45 333 48 336 
rect 45 336 48 339 
rect 45 339 48 342 
rect 45 342 48 345 
rect 45 345 48 348 
rect 45 348 48 351 
rect 45 351 48 354 
rect 45 354 48 357 
rect 45 357 48 360 
rect 45 360 48 363 
rect 45 363 48 366 
rect 45 366 48 369 
rect 45 369 48 372 
rect 45 372 48 375 
rect 45 375 48 378 
rect 45 378 48 381 
rect 45 381 48 384 
rect 45 384 48 387 
rect 45 387 48 390 
rect 45 390 48 393 
rect 45 393 48 396 
rect 45 396 48 399 
rect 45 399 48 402 
rect 45 402 48 405 
rect 45 405 48 408 
rect 45 408 48 411 
rect 45 411 48 414 
rect 45 414 48 417 
rect 45 417 48 420 
rect 45 420 48 423 
rect 45 423 48 426 
rect 45 426 48 429 
rect 45 429 48 432 
rect 45 432 48 435 
rect 45 435 48 438 
rect 45 438 48 441 
rect 45 441 48 444 
rect 45 444 48 447 
rect 45 447 48 450 
rect 45 450 48 453 
rect 45 453 48 456 
rect 45 456 48 459 
rect 45 459 48 462 
rect 45 462 48 465 
rect 45 465 48 468 
rect 45 468 48 471 
rect 45 471 48 474 
rect 45 474 48 477 
rect 45 477 48 480 
rect 45 480 48 483 
rect 45 483 48 486 
rect 45 486 48 489 
rect 45 489 48 492 
rect 45 492 48 495 
rect 45 495 48 498 
rect 45 498 48 501 
rect 45 501 48 504 
rect 45 504 48 507 
rect 45 507 48 510 
rect 48 0 51 3 
rect 48 3 51 6 
rect 48 6 51 9 
rect 48 9 51 12 
rect 48 12 51 15 
rect 48 15 51 18 
rect 48 18 51 21 
rect 48 21 51 24 
rect 48 24 51 27 
rect 48 27 51 30 
rect 48 30 51 33 
rect 48 33 51 36 
rect 48 36 51 39 
rect 48 39 51 42 
rect 48 42 51 45 
rect 48 45 51 48 
rect 48 48 51 51 
rect 48 51 51 54 
rect 48 54 51 57 
rect 48 57 51 60 
rect 48 60 51 63 
rect 48 63 51 66 
rect 48 66 51 69 
rect 48 69 51 72 
rect 48 72 51 75 
rect 48 75 51 78 
rect 48 78 51 81 
rect 48 81 51 84 
rect 48 84 51 87 
rect 48 87 51 90 
rect 48 90 51 93 
rect 48 93 51 96 
rect 48 96 51 99 
rect 48 99 51 102 
rect 48 102 51 105 
rect 48 105 51 108 
rect 48 108 51 111 
rect 48 111 51 114 
rect 48 114 51 117 
rect 48 117 51 120 
rect 48 120 51 123 
rect 48 123 51 126 
rect 48 126 51 129 
rect 48 129 51 132 
rect 48 132 51 135 
rect 48 135 51 138 
rect 48 138 51 141 
rect 48 141 51 144 
rect 48 144 51 147 
rect 48 147 51 150 
rect 48 150 51 153 
rect 48 153 51 156 
rect 48 156 51 159 
rect 48 159 51 162 
rect 48 162 51 165 
rect 48 165 51 168 
rect 48 168 51 171 
rect 48 171 51 174 
rect 48 174 51 177 
rect 48 177 51 180 
rect 48 180 51 183 
rect 48 183 51 186 
rect 48 186 51 189 
rect 48 189 51 192 
rect 48 192 51 195 
rect 48 195 51 198 
rect 48 198 51 201 
rect 48 201 51 204 
rect 48 204 51 207 
rect 48 207 51 210 
rect 48 210 51 213 
rect 48 213 51 216 
rect 48 216 51 219 
rect 48 219 51 222 
rect 48 222 51 225 
rect 48 225 51 228 
rect 48 228 51 231 
rect 48 231 51 234 
rect 48 234 51 237 
rect 48 237 51 240 
rect 48 240 51 243 
rect 48 243 51 246 
rect 48 246 51 249 
rect 48 249 51 252 
rect 48 252 51 255 
rect 48 255 51 258 
rect 48 258 51 261 
rect 48 261 51 264 
rect 48 264 51 267 
rect 48 267 51 270 
rect 48 270 51 273 
rect 48 273 51 276 
rect 48 276 51 279 
rect 48 279 51 282 
rect 48 282 51 285 
rect 48 285 51 288 
rect 48 288 51 291 
rect 48 291 51 294 
rect 48 294 51 297 
rect 48 297 51 300 
rect 48 300 51 303 
rect 48 303 51 306 
rect 48 306 51 309 
rect 48 309 51 312 
rect 48 312 51 315 
rect 48 315 51 318 
rect 48 318 51 321 
rect 48 321 51 324 
rect 48 324 51 327 
rect 48 327 51 330 
rect 48 330 51 333 
rect 48 333 51 336 
rect 48 336 51 339 
rect 48 339 51 342 
rect 48 342 51 345 
rect 48 345 51 348 
rect 48 348 51 351 
rect 48 351 51 354 
rect 48 354 51 357 
rect 48 357 51 360 
rect 48 360 51 363 
rect 48 363 51 366 
rect 48 366 51 369 
rect 48 369 51 372 
rect 48 372 51 375 
rect 48 375 51 378 
rect 48 378 51 381 
rect 48 381 51 384 
rect 48 384 51 387 
rect 48 387 51 390 
rect 48 390 51 393 
rect 48 393 51 396 
rect 48 396 51 399 
rect 48 399 51 402 
rect 48 402 51 405 
rect 48 405 51 408 
rect 48 408 51 411 
rect 48 411 51 414 
rect 48 414 51 417 
rect 48 417 51 420 
rect 48 420 51 423 
rect 48 423 51 426 
rect 48 426 51 429 
rect 48 429 51 432 
rect 48 432 51 435 
rect 48 435 51 438 
rect 48 438 51 441 
rect 48 441 51 444 
rect 48 444 51 447 
rect 48 447 51 450 
rect 48 450 51 453 
rect 48 453 51 456 
rect 48 456 51 459 
rect 48 459 51 462 
rect 48 462 51 465 
rect 48 465 51 468 
rect 48 468 51 471 
rect 48 471 51 474 
rect 48 474 51 477 
rect 48 477 51 480 
rect 48 480 51 483 
rect 48 483 51 486 
rect 48 486 51 489 
rect 48 489 51 492 
rect 48 492 51 495 
rect 48 495 51 498 
rect 48 498 51 501 
rect 48 501 51 504 
rect 48 504 51 507 
rect 48 507 51 510 
rect 51 0 54 3 
rect 51 3 54 6 
rect 51 6 54 9 
rect 51 9 54 12 
rect 51 12 54 15 
rect 51 15 54 18 
rect 51 18 54 21 
rect 51 21 54 24 
rect 51 24 54 27 
rect 51 27 54 30 
rect 51 30 54 33 
rect 51 33 54 36 
rect 51 36 54 39 
rect 51 39 54 42 
rect 51 42 54 45 
rect 51 45 54 48 
rect 51 48 54 51 
rect 51 51 54 54 
rect 51 54 54 57 
rect 51 57 54 60 
rect 51 60 54 63 
rect 51 63 54 66 
rect 51 66 54 69 
rect 51 69 54 72 
rect 51 72 54 75 
rect 51 75 54 78 
rect 51 78 54 81 
rect 51 81 54 84 
rect 51 84 54 87 
rect 51 87 54 90 
rect 51 90 54 93 
rect 51 93 54 96 
rect 51 96 54 99 
rect 51 99 54 102 
rect 51 102 54 105 
rect 51 105 54 108 
rect 51 108 54 111 
rect 51 111 54 114 
rect 51 114 54 117 
rect 51 117 54 120 
rect 51 120 54 123 
rect 51 123 54 126 
rect 51 126 54 129 
rect 51 129 54 132 
rect 51 132 54 135 
rect 51 135 54 138 
rect 51 138 54 141 
rect 51 141 54 144 
rect 51 144 54 147 
rect 51 147 54 150 
rect 51 150 54 153 
rect 51 153 54 156 
rect 51 156 54 159 
rect 51 159 54 162 
rect 51 162 54 165 
rect 51 165 54 168 
rect 51 168 54 171 
rect 51 171 54 174 
rect 51 174 54 177 
rect 51 177 54 180 
rect 51 180 54 183 
rect 51 183 54 186 
rect 51 186 54 189 
rect 51 189 54 192 
rect 51 192 54 195 
rect 51 195 54 198 
rect 51 198 54 201 
rect 51 201 54 204 
rect 51 204 54 207 
rect 51 207 54 210 
rect 51 210 54 213 
rect 51 213 54 216 
rect 51 216 54 219 
rect 51 219 54 222 
rect 51 222 54 225 
rect 51 225 54 228 
rect 51 228 54 231 
rect 51 231 54 234 
rect 51 234 54 237 
rect 51 237 54 240 
rect 51 240 54 243 
rect 51 243 54 246 
rect 51 246 54 249 
rect 51 249 54 252 
rect 51 252 54 255 
rect 51 255 54 258 
rect 51 258 54 261 
rect 51 261 54 264 
rect 51 264 54 267 
rect 51 267 54 270 
rect 51 270 54 273 
rect 51 273 54 276 
rect 51 276 54 279 
rect 51 279 54 282 
rect 51 282 54 285 
rect 51 285 54 288 
rect 51 288 54 291 
rect 51 291 54 294 
rect 51 294 54 297 
rect 51 297 54 300 
rect 51 300 54 303 
rect 51 303 54 306 
rect 51 306 54 309 
rect 51 309 54 312 
rect 51 312 54 315 
rect 51 315 54 318 
rect 51 318 54 321 
rect 51 321 54 324 
rect 51 324 54 327 
rect 51 327 54 330 
rect 51 330 54 333 
rect 51 333 54 336 
rect 51 336 54 339 
rect 51 339 54 342 
rect 51 342 54 345 
rect 51 345 54 348 
rect 51 348 54 351 
rect 51 351 54 354 
rect 51 354 54 357 
rect 51 357 54 360 
rect 51 360 54 363 
rect 51 363 54 366 
rect 51 366 54 369 
rect 51 369 54 372 
rect 51 372 54 375 
rect 51 375 54 378 
rect 51 378 54 381 
rect 51 381 54 384 
rect 51 384 54 387 
rect 51 387 54 390 
rect 51 390 54 393 
rect 51 393 54 396 
rect 51 396 54 399 
rect 51 399 54 402 
rect 51 402 54 405 
rect 51 405 54 408 
rect 51 408 54 411 
rect 51 411 54 414 
rect 51 414 54 417 
rect 51 417 54 420 
rect 51 420 54 423 
rect 51 423 54 426 
rect 51 426 54 429 
rect 51 429 54 432 
rect 51 432 54 435 
rect 51 435 54 438 
rect 51 438 54 441 
rect 51 441 54 444 
rect 51 444 54 447 
rect 51 447 54 450 
rect 51 450 54 453 
rect 51 453 54 456 
rect 51 456 54 459 
rect 51 459 54 462 
rect 51 462 54 465 
rect 51 465 54 468 
rect 51 468 54 471 
rect 51 471 54 474 
rect 51 474 54 477 
rect 51 477 54 480 
rect 51 480 54 483 
rect 51 483 54 486 
rect 51 486 54 489 
rect 51 489 54 492 
rect 51 492 54 495 
rect 51 495 54 498 
rect 51 498 54 501 
rect 51 501 54 504 
rect 51 504 54 507 
rect 51 507 54 510 
rect 54 0 57 3 
rect 54 3 57 6 
rect 54 6 57 9 
rect 54 9 57 12 
rect 54 12 57 15 
rect 54 15 57 18 
rect 54 18 57 21 
rect 54 21 57 24 
rect 54 24 57 27 
rect 54 27 57 30 
rect 54 30 57 33 
rect 54 33 57 36 
rect 54 36 57 39 
rect 54 39 57 42 
rect 54 42 57 45 
rect 54 45 57 48 
rect 54 48 57 51 
rect 54 51 57 54 
rect 54 54 57 57 
rect 54 57 57 60 
rect 54 60 57 63 
rect 54 63 57 66 
rect 54 66 57 69 
rect 54 69 57 72 
rect 54 72 57 75 
rect 54 75 57 78 
rect 54 78 57 81 
rect 54 81 57 84 
rect 54 84 57 87 
rect 54 87 57 90 
rect 54 90 57 93 
rect 54 93 57 96 
rect 54 96 57 99 
rect 54 99 57 102 
rect 54 102 57 105 
rect 54 105 57 108 
rect 54 108 57 111 
rect 54 111 57 114 
rect 54 114 57 117 
rect 54 117 57 120 
rect 54 120 57 123 
rect 54 123 57 126 
rect 54 126 57 129 
rect 54 129 57 132 
rect 54 132 57 135 
rect 54 135 57 138 
rect 54 138 57 141 
rect 54 141 57 144 
rect 54 144 57 147 
rect 54 147 57 150 
rect 54 150 57 153 
rect 54 153 57 156 
rect 54 156 57 159 
rect 54 159 57 162 
rect 54 162 57 165 
rect 54 165 57 168 
rect 54 168 57 171 
rect 54 171 57 174 
rect 54 174 57 177 
rect 54 177 57 180 
rect 54 180 57 183 
rect 54 183 57 186 
rect 54 186 57 189 
rect 54 189 57 192 
rect 54 192 57 195 
rect 54 195 57 198 
rect 54 198 57 201 
rect 54 201 57 204 
rect 54 204 57 207 
rect 54 207 57 210 
rect 54 210 57 213 
rect 54 213 57 216 
rect 54 216 57 219 
rect 54 219 57 222 
rect 54 222 57 225 
rect 54 225 57 228 
rect 54 228 57 231 
rect 54 231 57 234 
rect 54 234 57 237 
rect 54 237 57 240 
rect 54 240 57 243 
rect 54 243 57 246 
rect 54 246 57 249 
rect 54 249 57 252 
rect 54 252 57 255 
rect 54 255 57 258 
rect 54 258 57 261 
rect 54 261 57 264 
rect 54 264 57 267 
rect 54 267 57 270 
rect 54 270 57 273 
rect 54 273 57 276 
rect 54 276 57 279 
rect 54 279 57 282 
rect 54 282 57 285 
rect 54 285 57 288 
rect 54 288 57 291 
rect 54 291 57 294 
rect 54 294 57 297 
rect 54 297 57 300 
rect 54 300 57 303 
rect 54 303 57 306 
rect 54 306 57 309 
rect 54 309 57 312 
rect 54 312 57 315 
rect 54 315 57 318 
rect 54 318 57 321 
rect 54 321 57 324 
rect 54 324 57 327 
rect 54 327 57 330 
rect 54 330 57 333 
rect 54 333 57 336 
rect 54 336 57 339 
rect 54 339 57 342 
rect 54 342 57 345 
rect 54 345 57 348 
rect 54 348 57 351 
rect 54 351 57 354 
rect 54 354 57 357 
rect 54 357 57 360 
rect 54 360 57 363 
rect 54 363 57 366 
rect 54 366 57 369 
rect 54 369 57 372 
rect 54 372 57 375 
rect 54 375 57 378 
rect 54 378 57 381 
rect 54 381 57 384 
rect 54 384 57 387 
rect 54 387 57 390 
rect 54 390 57 393 
rect 54 393 57 396 
rect 54 396 57 399 
rect 54 399 57 402 
rect 54 402 57 405 
rect 54 405 57 408 
rect 54 408 57 411 
rect 54 411 57 414 
rect 54 414 57 417 
rect 54 417 57 420 
rect 54 420 57 423 
rect 54 423 57 426 
rect 54 426 57 429 
rect 54 429 57 432 
rect 54 432 57 435 
rect 54 435 57 438 
rect 54 438 57 441 
rect 54 441 57 444 
rect 54 444 57 447 
rect 54 447 57 450 
rect 54 450 57 453 
rect 54 453 57 456 
rect 54 456 57 459 
rect 54 459 57 462 
rect 54 462 57 465 
rect 54 465 57 468 
rect 54 468 57 471 
rect 54 471 57 474 
rect 54 474 57 477 
rect 54 477 57 480 
rect 54 480 57 483 
rect 54 483 57 486 
rect 54 486 57 489 
rect 54 489 57 492 
rect 54 492 57 495 
rect 54 495 57 498 
rect 54 498 57 501 
rect 54 501 57 504 
rect 54 504 57 507 
rect 54 507 57 510 
rect 57 0 60 3 
rect 57 3 60 6 
rect 57 6 60 9 
rect 57 9 60 12 
rect 57 12 60 15 
rect 57 15 60 18 
rect 57 18 60 21 
rect 57 21 60 24 
rect 57 24 60 27 
rect 57 27 60 30 
rect 57 30 60 33 
rect 57 33 60 36 
rect 57 36 60 39 
rect 57 39 60 42 
rect 57 42 60 45 
rect 57 45 60 48 
rect 57 48 60 51 
rect 57 51 60 54 
rect 57 54 60 57 
rect 57 57 60 60 
rect 57 60 60 63 
rect 57 63 60 66 
rect 57 66 60 69 
rect 57 69 60 72 
rect 57 72 60 75 
rect 57 75 60 78 
rect 57 78 60 81 
rect 57 81 60 84 
rect 57 84 60 87 
rect 57 87 60 90 
rect 57 90 60 93 
rect 57 93 60 96 
rect 57 96 60 99 
rect 57 99 60 102 
rect 57 102 60 105 
rect 57 105 60 108 
rect 57 108 60 111 
rect 57 111 60 114 
rect 57 114 60 117 
rect 57 117 60 120 
rect 57 120 60 123 
rect 57 123 60 126 
rect 57 126 60 129 
rect 57 129 60 132 
rect 57 132 60 135 
rect 57 135 60 138 
rect 57 138 60 141 
rect 57 141 60 144 
rect 57 144 60 147 
rect 57 147 60 150 
rect 57 150 60 153 
rect 57 153 60 156 
rect 57 156 60 159 
rect 57 159 60 162 
rect 57 162 60 165 
rect 57 165 60 168 
rect 57 168 60 171 
rect 57 171 60 174 
rect 57 174 60 177 
rect 57 177 60 180 
rect 57 180 60 183 
rect 57 183 60 186 
rect 57 186 60 189 
rect 57 189 60 192 
rect 57 192 60 195 
rect 57 195 60 198 
rect 57 198 60 201 
rect 57 201 60 204 
rect 57 204 60 207 
rect 57 207 60 210 
rect 57 210 60 213 
rect 57 213 60 216 
rect 57 216 60 219 
rect 57 219 60 222 
rect 57 222 60 225 
rect 57 225 60 228 
rect 57 228 60 231 
rect 57 231 60 234 
rect 57 234 60 237 
rect 57 237 60 240 
rect 57 240 60 243 
rect 57 243 60 246 
rect 57 246 60 249 
rect 57 249 60 252 
rect 57 252 60 255 
rect 57 255 60 258 
rect 57 258 60 261 
rect 57 261 60 264 
rect 57 264 60 267 
rect 57 267 60 270 
rect 57 270 60 273 
rect 57 273 60 276 
rect 57 276 60 279 
rect 57 279 60 282 
rect 57 282 60 285 
rect 57 285 60 288 
rect 57 288 60 291 
rect 57 291 60 294 
rect 57 294 60 297 
rect 57 297 60 300 
rect 57 300 60 303 
rect 57 303 60 306 
rect 57 306 60 309 
rect 57 309 60 312 
rect 57 312 60 315 
rect 57 315 60 318 
rect 57 318 60 321 
rect 57 321 60 324 
rect 57 324 60 327 
rect 57 327 60 330 
rect 57 330 60 333 
rect 57 333 60 336 
rect 57 336 60 339 
rect 57 339 60 342 
rect 57 342 60 345 
rect 57 345 60 348 
rect 57 348 60 351 
rect 57 351 60 354 
rect 57 354 60 357 
rect 57 357 60 360 
rect 57 360 60 363 
rect 57 363 60 366 
rect 57 366 60 369 
rect 57 369 60 372 
rect 57 372 60 375 
rect 57 375 60 378 
rect 57 378 60 381 
rect 57 381 60 384 
rect 57 384 60 387 
rect 57 387 60 390 
rect 57 390 60 393 
rect 57 393 60 396 
rect 57 396 60 399 
rect 57 399 60 402 
rect 57 402 60 405 
rect 57 405 60 408 
rect 57 408 60 411 
rect 57 411 60 414 
rect 57 414 60 417 
rect 57 417 60 420 
rect 57 420 60 423 
rect 57 423 60 426 
rect 57 426 60 429 
rect 57 429 60 432 
rect 57 432 60 435 
rect 57 435 60 438 
rect 57 438 60 441 
rect 57 441 60 444 
rect 57 444 60 447 
rect 57 447 60 450 
rect 57 450 60 453 
rect 57 453 60 456 
rect 57 456 60 459 
rect 57 459 60 462 
rect 57 462 60 465 
rect 57 465 60 468 
rect 57 468 60 471 
rect 57 471 60 474 
rect 57 474 60 477 
rect 57 477 60 480 
rect 57 480 60 483 
rect 57 483 60 486 
rect 57 486 60 489 
rect 57 489 60 492 
rect 57 492 60 495 
rect 57 495 60 498 
rect 57 498 60 501 
rect 57 501 60 504 
rect 57 504 60 507 
rect 57 507 60 510 
rect 60 0 63 3 
rect 60 3 63 6 
rect 60 6 63 9 
rect 60 9 63 12 
rect 60 12 63 15 
rect 60 15 63 18 
rect 60 18 63 21 
rect 60 21 63 24 
rect 60 24 63 27 
rect 60 27 63 30 
rect 60 30 63 33 
rect 60 33 63 36 
rect 60 36 63 39 
rect 60 39 63 42 
rect 60 42 63 45 
rect 60 45 63 48 
rect 60 48 63 51 
rect 60 51 63 54 
rect 60 54 63 57 
rect 60 57 63 60 
rect 60 60 63 63 
rect 60 63 63 66 
rect 60 66 63 69 
rect 60 69 63 72 
rect 60 72 63 75 
rect 60 75 63 78 
rect 60 78 63 81 
rect 60 81 63 84 
rect 60 84 63 87 
rect 60 87 63 90 
rect 60 90 63 93 
rect 60 93 63 96 
rect 60 96 63 99 
rect 60 99 63 102 
rect 60 102 63 105 
rect 60 105 63 108 
rect 60 108 63 111 
rect 60 111 63 114 
rect 60 114 63 117 
rect 60 117 63 120 
rect 60 120 63 123 
rect 60 123 63 126 
rect 60 126 63 129 
rect 60 129 63 132 
rect 60 132 63 135 
rect 60 135 63 138 
rect 60 138 63 141 
rect 60 141 63 144 
rect 60 144 63 147 
rect 60 147 63 150 
rect 60 150 63 153 
rect 60 153 63 156 
rect 60 156 63 159 
rect 60 159 63 162 
rect 60 162 63 165 
rect 60 165 63 168 
rect 60 168 63 171 
rect 60 171 63 174 
rect 60 174 63 177 
rect 60 177 63 180 
rect 60 180 63 183 
rect 60 183 63 186 
rect 60 186 63 189 
rect 60 189 63 192 
rect 60 192 63 195 
rect 60 195 63 198 
rect 60 198 63 201 
rect 60 201 63 204 
rect 60 204 63 207 
rect 60 207 63 210 
rect 60 210 63 213 
rect 60 213 63 216 
rect 60 216 63 219 
rect 60 219 63 222 
rect 60 222 63 225 
rect 60 225 63 228 
rect 60 228 63 231 
rect 60 231 63 234 
rect 60 234 63 237 
rect 60 237 63 240 
rect 60 240 63 243 
rect 60 243 63 246 
rect 60 246 63 249 
rect 60 249 63 252 
rect 60 252 63 255 
rect 60 255 63 258 
rect 60 258 63 261 
rect 60 261 63 264 
rect 60 264 63 267 
rect 60 267 63 270 
rect 60 270 63 273 
rect 60 273 63 276 
rect 60 276 63 279 
rect 60 279 63 282 
rect 60 282 63 285 
rect 60 285 63 288 
rect 60 288 63 291 
rect 60 291 63 294 
rect 60 294 63 297 
rect 60 297 63 300 
rect 60 300 63 303 
rect 60 303 63 306 
rect 60 306 63 309 
rect 60 309 63 312 
rect 60 312 63 315 
rect 60 315 63 318 
rect 60 318 63 321 
rect 60 321 63 324 
rect 60 324 63 327 
rect 60 327 63 330 
rect 60 330 63 333 
rect 60 333 63 336 
rect 60 336 63 339 
rect 60 339 63 342 
rect 60 342 63 345 
rect 60 345 63 348 
rect 60 348 63 351 
rect 60 351 63 354 
rect 60 354 63 357 
rect 60 357 63 360 
rect 60 360 63 363 
rect 60 363 63 366 
rect 60 366 63 369 
rect 60 369 63 372 
rect 60 372 63 375 
rect 60 375 63 378 
rect 60 378 63 381 
rect 60 381 63 384 
rect 60 384 63 387 
rect 60 387 63 390 
rect 60 390 63 393 
rect 60 393 63 396 
rect 60 396 63 399 
rect 60 399 63 402 
rect 60 402 63 405 
rect 60 405 63 408 
rect 60 408 63 411 
rect 60 411 63 414 
rect 60 414 63 417 
rect 60 417 63 420 
rect 60 420 63 423 
rect 60 423 63 426 
rect 60 426 63 429 
rect 60 429 63 432 
rect 60 432 63 435 
rect 60 435 63 438 
rect 60 438 63 441 
rect 60 441 63 444 
rect 60 444 63 447 
rect 60 447 63 450 
rect 60 450 63 453 
rect 60 453 63 456 
rect 60 456 63 459 
rect 60 459 63 462 
rect 60 462 63 465 
rect 60 465 63 468 
rect 60 468 63 471 
rect 60 471 63 474 
rect 60 474 63 477 
rect 60 477 63 480 
rect 60 480 63 483 
rect 60 483 63 486 
rect 60 486 63 489 
rect 60 489 63 492 
rect 60 492 63 495 
rect 60 495 63 498 
rect 60 498 63 501 
rect 60 501 63 504 
rect 60 504 63 507 
rect 60 507 63 510 
rect 63 0 66 3 
rect 63 3 66 6 
rect 63 6 66 9 
rect 63 9 66 12 
rect 63 12 66 15 
rect 63 15 66 18 
rect 63 18 66 21 
rect 63 21 66 24 
rect 63 24 66 27 
rect 63 27 66 30 
rect 63 30 66 33 
rect 63 33 66 36 
rect 63 36 66 39 
rect 63 39 66 42 
rect 63 42 66 45 
rect 63 45 66 48 
rect 63 48 66 51 
rect 63 51 66 54 
rect 63 54 66 57 
rect 63 57 66 60 
rect 63 60 66 63 
rect 63 63 66 66 
rect 63 66 66 69 
rect 63 69 66 72 
rect 63 72 66 75 
rect 63 75 66 78 
rect 63 78 66 81 
rect 63 81 66 84 
rect 63 84 66 87 
rect 63 87 66 90 
rect 63 90 66 93 
rect 63 93 66 96 
rect 63 96 66 99 
rect 63 99 66 102 
rect 63 102 66 105 
rect 63 105 66 108 
rect 63 108 66 111 
rect 63 111 66 114 
rect 63 114 66 117 
rect 63 117 66 120 
rect 63 120 66 123 
rect 63 123 66 126 
rect 63 126 66 129 
rect 63 129 66 132 
rect 63 132 66 135 
rect 63 135 66 138 
rect 63 138 66 141 
rect 63 141 66 144 
rect 63 144 66 147 
rect 63 147 66 150 
rect 63 150 66 153 
rect 63 153 66 156 
rect 63 156 66 159 
rect 63 159 66 162 
rect 63 162 66 165 
rect 63 165 66 168 
rect 63 168 66 171 
rect 63 171 66 174 
rect 63 174 66 177 
rect 63 177 66 180 
rect 63 180 66 183 
rect 63 183 66 186 
rect 63 186 66 189 
rect 63 189 66 192 
rect 63 192 66 195 
rect 63 195 66 198 
rect 63 198 66 201 
rect 63 201 66 204 
rect 63 204 66 207 
rect 63 207 66 210 
rect 63 210 66 213 
rect 63 213 66 216 
rect 63 216 66 219 
rect 63 219 66 222 
rect 63 222 66 225 
rect 63 225 66 228 
rect 63 228 66 231 
rect 63 231 66 234 
rect 63 234 66 237 
rect 63 237 66 240 
rect 63 240 66 243 
rect 63 243 66 246 
rect 63 246 66 249 
rect 63 249 66 252 
rect 63 252 66 255 
rect 63 255 66 258 
rect 63 258 66 261 
rect 63 261 66 264 
rect 63 264 66 267 
rect 63 267 66 270 
rect 63 270 66 273 
rect 63 273 66 276 
rect 63 276 66 279 
rect 63 279 66 282 
rect 63 282 66 285 
rect 63 285 66 288 
rect 63 288 66 291 
rect 63 291 66 294 
rect 63 294 66 297 
rect 63 297 66 300 
rect 63 300 66 303 
rect 63 303 66 306 
rect 63 306 66 309 
rect 63 309 66 312 
rect 63 312 66 315 
rect 63 315 66 318 
rect 63 318 66 321 
rect 63 321 66 324 
rect 63 324 66 327 
rect 63 327 66 330 
rect 63 330 66 333 
rect 63 333 66 336 
rect 63 336 66 339 
rect 63 339 66 342 
rect 63 342 66 345 
rect 63 345 66 348 
rect 63 348 66 351 
rect 63 351 66 354 
rect 63 354 66 357 
rect 63 357 66 360 
rect 63 360 66 363 
rect 63 363 66 366 
rect 63 366 66 369 
rect 63 369 66 372 
rect 63 372 66 375 
rect 63 375 66 378 
rect 63 378 66 381 
rect 63 381 66 384 
rect 63 384 66 387 
rect 63 387 66 390 
rect 63 390 66 393 
rect 63 393 66 396 
rect 63 396 66 399 
rect 63 399 66 402 
rect 63 402 66 405 
rect 63 405 66 408 
rect 63 408 66 411 
rect 63 411 66 414 
rect 63 414 66 417 
rect 63 417 66 420 
rect 63 420 66 423 
rect 63 423 66 426 
rect 63 426 66 429 
rect 63 429 66 432 
rect 63 432 66 435 
rect 63 435 66 438 
rect 63 438 66 441 
rect 63 441 66 444 
rect 63 444 66 447 
rect 63 447 66 450 
rect 63 450 66 453 
rect 63 453 66 456 
rect 63 456 66 459 
rect 63 459 66 462 
rect 63 462 66 465 
rect 63 465 66 468 
rect 63 468 66 471 
rect 63 471 66 474 
rect 63 474 66 477 
rect 63 477 66 480 
rect 63 480 66 483 
rect 63 483 66 486 
rect 63 486 66 489 
rect 63 489 66 492 
rect 63 492 66 495 
rect 63 495 66 498 
rect 63 498 66 501 
rect 63 501 66 504 
rect 63 504 66 507 
rect 63 507 66 510 
rect 66 0 69 3 
rect 66 3 69 6 
rect 66 6 69 9 
rect 66 9 69 12 
rect 66 12 69 15 
rect 66 15 69 18 
rect 66 18 69 21 
rect 66 21 69 24 
rect 66 24 69 27 
rect 66 27 69 30 
rect 66 30 69 33 
rect 66 33 69 36 
rect 66 36 69 39 
rect 66 39 69 42 
rect 66 42 69 45 
rect 66 45 69 48 
rect 66 48 69 51 
rect 66 51 69 54 
rect 66 54 69 57 
rect 66 57 69 60 
rect 66 60 69 63 
rect 66 63 69 66 
rect 66 66 69 69 
rect 66 69 69 72 
rect 66 72 69 75 
rect 66 75 69 78 
rect 66 78 69 81 
rect 66 81 69 84 
rect 66 84 69 87 
rect 66 87 69 90 
rect 66 90 69 93 
rect 66 93 69 96 
rect 66 96 69 99 
rect 66 99 69 102 
rect 66 102 69 105 
rect 66 105 69 108 
rect 66 108 69 111 
rect 66 111 69 114 
rect 66 114 69 117 
rect 66 117 69 120 
rect 66 120 69 123 
rect 66 123 69 126 
rect 66 126 69 129 
rect 66 129 69 132 
rect 66 132 69 135 
rect 66 135 69 138 
rect 66 138 69 141 
rect 66 141 69 144 
rect 66 144 69 147 
rect 66 147 69 150 
rect 66 150 69 153 
rect 66 153 69 156 
rect 66 156 69 159 
rect 66 159 69 162 
rect 66 162 69 165 
rect 66 165 69 168 
rect 66 168 69 171 
rect 66 171 69 174 
rect 66 174 69 177 
rect 66 177 69 180 
rect 66 180 69 183 
rect 66 183 69 186 
rect 66 186 69 189 
rect 66 189 69 192 
rect 66 192 69 195 
rect 66 195 69 198 
rect 66 198 69 201 
rect 66 201 69 204 
rect 66 204 69 207 
rect 66 207 69 210 
rect 66 210 69 213 
rect 66 213 69 216 
rect 66 216 69 219 
rect 66 219 69 222 
rect 66 222 69 225 
rect 66 225 69 228 
rect 66 228 69 231 
rect 66 231 69 234 
rect 66 234 69 237 
rect 66 237 69 240 
rect 66 240 69 243 
rect 66 243 69 246 
rect 66 246 69 249 
rect 66 249 69 252 
rect 66 252 69 255 
rect 66 255 69 258 
rect 66 258 69 261 
rect 66 261 69 264 
rect 66 264 69 267 
rect 66 267 69 270 
rect 66 270 69 273 
rect 66 273 69 276 
rect 66 276 69 279 
rect 66 279 69 282 
rect 66 282 69 285 
rect 66 285 69 288 
rect 66 288 69 291 
rect 66 291 69 294 
rect 66 294 69 297 
rect 66 297 69 300 
rect 66 300 69 303 
rect 66 303 69 306 
rect 66 306 69 309 
rect 66 309 69 312 
rect 66 312 69 315 
rect 66 315 69 318 
rect 66 318 69 321 
rect 66 321 69 324 
rect 66 324 69 327 
rect 66 327 69 330 
rect 66 330 69 333 
rect 66 333 69 336 
rect 66 336 69 339 
rect 66 339 69 342 
rect 66 342 69 345 
rect 66 345 69 348 
rect 66 348 69 351 
rect 66 351 69 354 
rect 66 354 69 357 
rect 66 357 69 360 
rect 66 360 69 363 
rect 66 363 69 366 
rect 66 366 69 369 
rect 66 369 69 372 
rect 66 372 69 375 
rect 66 375 69 378 
rect 66 378 69 381 
rect 66 381 69 384 
rect 66 384 69 387 
rect 66 387 69 390 
rect 66 390 69 393 
rect 66 393 69 396 
rect 66 396 69 399 
rect 66 399 69 402 
rect 66 402 69 405 
rect 66 405 69 408 
rect 66 408 69 411 
rect 66 411 69 414 
rect 66 414 69 417 
rect 66 417 69 420 
rect 66 420 69 423 
rect 66 423 69 426 
rect 66 426 69 429 
rect 66 429 69 432 
rect 66 432 69 435 
rect 66 435 69 438 
rect 66 438 69 441 
rect 66 441 69 444 
rect 66 444 69 447 
rect 66 447 69 450 
rect 66 450 69 453 
rect 66 453 69 456 
rect 66 456 69 459 
rect 66 459 69 462 
rect 66 462 69 465 
rect 66 465 69 468 
rect 66 468 69 471 
rect 66 471 69 474 
rect 66 474 69 477 
rect 66 477 69 480 
rect 66 480 69 483 
rect 66 483 69 486 
rect 66 486 69 489 
rect 66 489 69 492 
rect 66 492 69 495 
rect 66 495 69 498 
rect 66 498 69 501 
rect 66 501 69 504 
rect 66 504 69 507 
rect 66 507 69 510 
rect 69 0 72 3 
rect 69 3 72 6 
rect 69 6 72 9 
rect 69 9 72 12 
rect 69 12 72 15 
rect 69 15 72 18 
rect 69 18 72 21 
rect 69 21 72 24 
rect 69 24 72 27 
rect 69 27 72 30 
rect 69 30 72 33 
rect 69 33 72 36 
rect 69 36 72 39 
rect 69 39 72 42 
rect 69 42 72 45 
rect 69 45 72 48 
rect 69 48 72 51 
rect 69 51 72 54 
rect 69 54 72 57 
rect 69 57 72 60 
rect 69 60 72 63 
rect 69 63 72 66 
rect 69 66 72 69 
rect 69 69 72 72 
rect 69 72 72 75 
rect 69 75 72 78 
rect 69 78 72 81 
rect 69 81 72 84 
rect 69 84 72 87 
rect 69 87 72 90 
rect 69 90 72 93 
rect 69 93 72 96 
rect 69 96 72 99 
rect 69 99 72 102 
rect 69 102 72 105 
rect 69 105 72 108 
rect 69 108 72 111 
rect 69 111 72 114 
rect 69 114 72 117 
rect 69 117 72 120 
rect 69 120 72 123 
rect 69 123 72 126 
rect 69 126 72 129 
rect 69 129 72 132 
rect 69 132 72 135 
rect 69 135 72 138 
rect 69 138 72 141 
rect 69 141 72 144 
rect 69 144 72 147 
rect 69 147 72 150 
rect 69 150 72 153 
rect 69 153 72 156 
rect 69 156 72 159 
rect 69 159 72 162 
rect 69 162 72 165 
rect 69 165 72 168 
rect 69 168 72 171 
rect 69 171 72 174 
rect 69 174 72 177 
rect 69 177 72 180 
rect 69 180 72 183 
rect 69 183 72 186 
rect 69 186 72 189 
rect 69 189 72 192 
rect 69 192 72 195 
rect 69 195 72 198 
rect 69 198 72 201 
rect 69 201 72 204 
rect 69 204 72 207 
rect 69 207 72 210 
rect 69 210 72 213 
rect 69 213 72 216 
rect 69 216 72 219 
rect 69 219 72 222 
rect 69 222 72 225 
rect 69 225 72 228 
rect 69 228 72 231 
rect 69 231 72 234 
rect 69 234 72 237 
rect 69 237 72 240 
rect 69 240 72 243 
rect 69 243 72 246 
rect 69 246 72 249 
rect 69 249 72 252 
rect 69 252 72 255 
rect 69 255 72 258 
rect 69 258 72 261 
rect 69 261 72 264 
rect 69 264 72 267 
rect 69 267 72 270 
rect 69 270 72 273 
rect 69 273 72 276 
rect 69 276 72 279 
rect 69 279 72 282 
rect 69 282 72 285 
rect 69 285 72 288 
rect 69 288 72 291 
rect 69 291 72 294 
rect 69 294 72 297 
rect 69 297 72 300 
rect 69 300 72 303 
rect 69 303 72 306 
rect 69 306 72 309 
rect 69 309 72 312 
rect 69 312 72 315 
rect 69 315 72 318 
rect 69 318 72 321 
rect 69 321 72 324 
rect 69 324 72 327 
rect 69 327 72 330 
rect 69 330 72 333 
rect 69 333 72 336 
rect 69 336 72 339 
rect 69 339 72 342 
rect 69 342 72 345 
rect 69 345 72 348 
rect 69 348 72 351 
rect 69 351 72 354 
rect 69 354 72 357 
rect 69 357 72 360 
rect 69 360 72 363 
rect 69 363 72 366 
rect 69 366 72 369 
rect 69 369 72 372 
rect 69 372 72 375 
rect 69 375 72 378 
rect 69 378 72 381 
rect 69 381 72 384 
rect 69 384 72 387 
rect 69 387 72 390 
rect 69 390 72 393 
rect 69 393 72 396 
rect 69 396 72 399 
rect 69 399 72 402 
rect 69 402 72 405 
rect 69 405 72 408 
rect 69 408 72 411 
rect 69 411 72 414 
rect 69 414 72 417 
rect 69 417 72 420 
rect 69 420 72 423 
rect 69 423 72 426 
rect 69 426 72 429 
rect 69 429 72 432 
rect 69 432 72 435 
rect 69 435 72 438 
rect 69 438 72 441 
rect 69 441 72 444 
rect 69 444 72 447 
rect 69 447 72 450 
rect 69 450 72 453 
rect 69 453 72 456 
rect 69 456 72 459 
rect 69 459 72 462 
rect 69 462 72 465 
rect 69 465 72 468 
rect 69 468 72 471 
rect 69 471 72 474 
rect 69 474 72 477 
rect 69 477 72 480 
rect 69 480 72 483 
rect 69 483 72 486 
rect 69 486 72 489 
rect 69 489 72 492 
rect 69 492 72 495 
rect 69 495 72 498 
rect 69 498 72 501 
rect 69 501 72 504 
rect 69 504 72 507 
rect 69 507 72 510 
rect 72 0 75 3 
rect 72 3 75 6 
rect 72 6 75 9 
rect 72 9 75 12 
rect 72 12 75 15 
rect 72 15 75 18 
rect 72 18 75 21 
rect 72 21 75 24 
rect 72 24 75 27 
rect 72 27 75 30 
rect 72 30 75 33 
rect 72 33 75 36 
rect 72 36 75 39 
rect 72 39 75 42 
rect 72 42 75 45 
rect 72 45 75 48 
rect 72 48 75 51 
rect 72 51 75 54 
rect 72 54 75 57 
rect 72 57 75 60 
rect 72 60 75 63 
rect 72 63 75 66 
rect 72 66 75 69 
rect 72 69 75 72 
rect 72 72 75 75 
rect 72 75 75 78 
rect 72 78 75 81 
rect 72 81 75 84 
rect 72 84 75 87 
rect 72 87 75 90 
rect 72 90 75 93 
rect 72 93 75 96 
rect 72 96 75 99 
rect 72 99 75 102 
rect 72 102 75 105 
rect 72 105 75 108 
rect 72 108 75 111 
rect 72 111 75 114 
rect 72 114 75 117 
rect 72 117 75 120 
rect 72 120 75 123 
rect 72 123 75 126 
rect 72 126 75 129 
rect 72 129 75 132 
rect 72 132 75 135 
rect 72 135 75 138 
rect 72 138 75 141 
rect 72 141 75 144 
rect 72 144 75 147 
rect 72 147 75 150 
rect 72 150 75 153 
rect 72 153 75 156 
rect 72 156 75 159 
rect 72 159 75 162 
rect 72 162 75 165 
rect 72 165 75 168 
rect 72 168 75 171 
rect 72 171 75 174 
rect 72 174 75 177 
rect 72 177 75 180 
rect 72 180 75 183 
rect 72 183 75 186 
rect 72 186 75 189 
rect 72 189 75 192 
rect 72 192 75 195 
rect 72 195 75 198 
rect 72 198 75 201 
rect 72 201 75 204 
rect 72 204 75 207 
rect 72 207 75 210 
rect 72 210 75 213 
rect 72 213 75 216 
rect 72 216 75 219 
rect 72 219 75 222 
rect 72 222 75 225 
rect 72 225 75 228 
rect 72 228 75 231 
rect 72 231 75 234 
rect 72 234 75 237 
rect 72 237 75 240 
rect 72 240 75 243 
rect 72 243 75 246 
rect 72 246 75 249 
rect 72 249 75 252 
rect 72 252 75 255 
rect 72 255 75 258 
rect 72 258 75 261 
rect 72 261 75 264 
rect 72 264 75 267 
rect 72 267 75 270 
rect 72 270 75 273 
rect 72 273 75 276 
rect 72 276 75 279 
rect 72 279 75 282 
rect 72 282 75 285 
rect 72 285 75 288 
rect 72 288 75 291 
rect 72 291 75 294 
rect 72 294 75 297 
rect 72 297 75 300 
rect 72 300 75 303 
rect 72 303 75 306 
rect 72 306 75 309 
rect 72 309 75 312 
rect 72 312 75 315 
rect 72 315 75 318 
rect 72 318 75 321 
rect 72 321 75 324 
rect 72 324 75 327 
rect 72 327 75 330 
rect 72 330 75 333 
rect 72 333 75 336 
rect 72 336 75 339 
rect 72 339 75 342 
rect 72 342 75 345 
rect 72 345 75 348 
rect 72 348 75 351 
rect 72 351 75 354 
rect 72 354 75 357 
rect 72 357 75 360 
rect 72 360 75 363 
rect 72 363 75 366 
rect 72 366 75 369 
rect 72 369 75 372 
rect 72 372 75 375 
rect 72 375 75 378 
rect 72 378 75 381 
rect 72 381 75 384 
rect 72 384 75 387 
rect 72 387 75 390 
rect 72 390 75 393 
rect 72 393 75 396 
rect 72 396 75 399 
rect 72 399 75 402 
rect 72 402 75 405 
rect 72 405 75 408 
rect 72 408 75 411 
rect 72 411 75 414 
rect 72 414 75 417 
rect 72 417 75 420 
rect 72 420 75 423 
rect 72 423 75 426 
rect 72 426 75 429 
rect 72 429 75 432 
rect 72 432 75 435 
rect 72 435 75 438 
rect 72 438 75 441 
rect 72 441 75 444 
rect 72 444 75 447 
rect 72 447 75 450 
rect 72 450 75 453 
rect 72 453 75 456 
rect 72 456 75 459 
rect 72 459 75 462 
rect 72 462 75 465 
rect 72 465 75 468 
rect 72 468 75 471 
rect 72 471 75 474 
rect 72 474 75 477 
rect 72 477 75 480 
rect 72 480 75 483 
rect 72 483 75 486 
rect 72 486 75 489 
rect 72 489 75 492 
rect 72 492 75 495 
rect 72 495 75 498 
rect 72 498 75 501 
rect 72 501 75 504 
rect 72 504 75 507 
rect 72 507 75 510 
rect 75 0 78 3 
rect 75 3 78 6 
rect 75 6 78 9 
rect 75 9 78 12 
rect 75 12 78 15 
rect 75 15 78 18 
rect 75 18 78 21 
rect 75 21 78 24 
rect 75 24 78 27 
rect 75 27 78 30 
rect 75 30 78 33 
rect 75 33 78 36 
rect 75 36 78 39 
rect 75 39 78 42 
rect 75 42 78 45 
rect 75 45 78 48 
rect 75 48 78 51 
rect 75 51 78 54 
rect 75 54 78 57 
rect 75 57 78 60 
rect 75 60 78 63 
rect 75 63 78 66 
rect 75 66 78 69 
rect 75 69 78 72 
rect 75 72 78 75 
rect 75 75 78 78 
rect 75 78 78 81 
rect 75 81 78 84 
rect 75 84 78 87 
rect 75 87 78 90 
rect 75 90 78 93 
rect 75 93 78 96 
rect 75 96 78 99 
rect 75 99 78 102 
rect 75 102 78 105 
rect 75 105 78 108 
rect 75 108 78 111 
rect 75 111 78 114 
rect 75 114 78 117 
rect 75 117 78 120 
rect 75 120 78 123 
rect 75 123 78 126 
rect 75 126 78 129 
rect 75 129 78 132 
rect 75 132 78 135 
rect 75 135 78 138 
rect 75 138 78 141 
rect 75 141 78 144 
rect 75 144 78 147 
rect 75 147 78 150 
rect 75 150 78 153 
rect 75 153 78 156 
rect 75 156 78 159 
rect 75 159 78 162 
rect 75 162 78 165 
rect 75 165 78 168 
rect 75 168 78 171 
rect 75 171 78 174 
rect 75 174 78 177 
rect 75 177 78 180 
rect 75 180 78 183 
rect 75 183 78 186 
rect 75 186 78 189 
rect 75 189 78 192 
rect 75 192 78 195 
rect 75 195 78 198 
rect 75 198 78 201 
rect 75 201 78 204 
rect 75 204 78 207 
rect 75 207 78 210 
rect 75 210 78 213 
rect 75 213 78 216 
rect 75 216 78 219 
rect 75 219 78 222 
rect 75 222 78 225 
rect 75 225 78 228 
rect 75 228 78 231 
rect 75 231 78 234 
rect 75 234 78 237 
rect 75 237 78 240 
rect 75 240 78 243 
rect 75 243 78 246 
rect 75 246 78 249 
rect 75 249 78 252 
rect 75 252 78 255 
rect 75 255 78 258 
rect 75 258 78 261 
rect 75 261 78 264 
rect 75 264 78 267 
rect 75 267 78 270 
rect 75 270 78 273 
rect 75 273 78 276 
rect 75 276 78 279 
rect 75 279 78 282 
rect 75 282 78 285 
rect 75 285 78 288 
rect 75 288 78 291 
rect 75 291 78 294 
rect 75 294 78 297 
rect 75 297 78 300 
rect 75 300 78 303 
rect 75 303 78 306 
rect 75 306 78 309 
rect 75 309 78 312 
rect 75 312 78 315 
rect 75 315 78 318 
rect 75 318 78 321 
rect 75 321 78 324 
rect 75 324 78 327 
rect 75 327 78 330 
rect 75 330 78 333 
rect 75 333 78 336 
rect 75 336 78 339 
rect 75 339 78 342 
rect 75 342 78 345 
rect 75 345 78 348 
rect 75 348 78 351 
rect 75 351 78 354 
rect 75 354 78 357 
rect 75 357 78 360 
rect 75 360 78 363 
rect 75 363 78 366 
rect 75 366 78 369 
rect 75 369 78 372 
rect 75 372 78 375 
rect 75 375 78 378 
rect 75 378 78 381 
rect 75 381 78 384 
rect 75 384 78 387 
rect 75 387 78 390 
rect 75 390 78 393 
rect 75 393 78 396 
rect 75 396 78 399 
rect 75 399 78 402 
rect 75 402 78 405 
rect 75 405 78 408 
rect 75 408 78 411 
rect 75 411 78 414 
rect 75 414 78 417 
rect 75 417 78 420 
rect 75 420 78 423 
rect 75 423 78 426 
rect 75 426 78 429 
rect 75 429 78 432 
rect 75 432 78 435 
rect 75 435 78 438 
rect 75 438 78 441 
rect 75 441 78 444 
rect 75 444 78 447 
rect 75 447 78 450 
rect 75 450 78 453 
rect 75 453 78 456 
rect 75 456 78 459 
rect 75 459 78 462 
rect 75 462 78 465 
rect 75 465 78 468 
rect 75 468 78 471 
rect 75 471 78 474 
rect 75 474 78 477 
rect 75 477 78 480 
rect 75 480 78 483 
rect 75 483 78 486 
rect 75 486 78 489 
rect 75 489 78 492 
rect 75 492 78 495 
rect 75 495 78 498 
rect 75 498 78 501 
rect 75 501 78 504 
rect 75 504 78 507 
rect 75 507 78 510 
rect 78 0 81 3 
rect 78 3 81 6 
rect 78 6 81 9 
rect 78 9 81 12 
rect 78 12 81 15 
rect 78 15 81 18 
rect 78 18 81 21 
rect 78 21 81 24 
rect 78 24 81 27 
rect 78 27 81 30 
rect 78 30 81 33 
rect 78 33 81 36 
rect 78 36 81 39 
rect 78 39 81 42 
rect 78 42 81 45 
rect 78 45 81 48 
rect 78 48 81 51 
rect 78 51 81 54 
rect 78 54 81 57 
rect 78 57 81 60 
rect 78 60 81 63 
rect 78 63 81 66 
rect 78 66 81 69 
rect 78 69 81 72 
rect 78 72 81 75 
rect 78 75 81 78 
rect 78 78 81 81 
rect 78 81 81 84 
rect 78 84 81 87 
rect 78 87 81 90 
rect 78 90 81 93 
rect 78 93 81 96 
rect 78 96 81 99 
rect 78 99 81 102 
rect 78 102 81 105 
rect 78 105 81 108 
rect 78 108 81 111 
rect 78 111 81 114 
rect 78 114 81 117 
rect 78 117 81 120 
rect 78 120 81 123 
rect 78 123 81 126 
rect 78 126 81 129 
rect 78 129 81 132 
rect 78 132 81 135 
rect 78 135 81 138 
rect 78 138 81 141 
rect 78 141 81 144 
rect 78 144 81 147 
rect 78 147 81 150 
rect 78 150 81 153 
rect 78 153 81 156 
rect 78 156 81 159 
rect 78 159 81 162 
rect 78 162 81 165 
rect 78 165 81 168 
rect 78 168 81 171 
rect 78 171 81 174 
rect 78 174 81 177 
rect 78 177 81 180 
rect 78 180 81 183 
rect 78 183 81 186 
rect 78 186 81 189 
rect 78 189 81 192 
rect 78 192 81 195 
rect 78 195 81 198 
rect 78 198 81 201 
rect 78 201 81 204 
rect 78 204 81 207 
rect 78 207 81 210 
rect 78 210 81 213 
rect 78 213 81 216 
rect 78 216 81 219 
rect 78 219 81 222 
rect 78 222 81 225 
rect 78 225 81 228 
rect 78 228 81 231 
rect 78 231 81 234 
rect 78 234 81 237 
rect 78 237 81 240 
rect 78 240 81 243 
rect 78 243 81 246 
rect 78 246 81 249 
rect 78 249 81 252 
rect 78 252 81 255 
rect 78 255 81 258 
rect 78 258 81 261 
rect 78 261 81 264 
rect 78 264 81 267 
rect 78 267 81 270 
rect 78 270 81 273 
rect 78 273 81 276 
rect 78 276 81 279 
rect 78 279 81 282 
rect 78 282 81 285 
rect 78 285 81 288 
rect 78 288 81 291 
rect 78 291 81 294 
rect 78 294 81 297 
rect 78 297 81 300 
rect 78 300 81 303 
rect 78 303 81 306 
rect 78 306 81 309 
rect 78 309 81 312 
rect 78 312 81 315 
rect 78 315 81 318 
rect 78 318 81 321 
rect 78 321 81 324 
rect 78 324 81 327 
rect 78 327 81 330 
rect 78 330 81 333 
rect 78 333 81 336 
rect 78 336 81 339 
rect 78 339 81 342 
rect 78 342 81 345 
rect 78 345 81 348 
rect 78 348 81 351 
rect 78 351 81 354 
rect 78 354 81 357 
rect 78 357 81 360 
rect 78 360 81 363 
rect 78 363 81 366 
rect 78 366 81 369 
rect 78 369 81 372 
rect 78 372 81 375 
rect 78 375 81 378 
rect 78 378 81 381 
rect 78 381 81 384 
rect 78 384 81 387 
rect 78 387 81 390 
rect 78 390 81 393 
rect 78 393 81 396 
rect 78 396 81 399 
rect 78 399 81 402 
rect 78 402 81 405 
rect 78 405 81 408 
rect 78 408 81 411 
rect 78 411 81 414 
rect 78 414 81 417 
rect 78 417 81 420 
rect 78 420 81 423 
rect 78 423 81 426 
rect 78 426 81 429 
rect 78 429 81 432 
rect 78 432 81 435 
rect 78 435 81 438 
rect 78 438 81 441 
rect 78 441 81 444 
rect 78 444 81 447 
rect 78 447 81 450 
rect 78 450 81 453 
rect 78 453 81 456 
rect 78 456 81 459 
rect 78 459 81 462 
rect 78 462 81 465 
rect 78 465 81 468 
rect 78 468 81 471 
rect 78 471 81 474 
rect 78 474 81 477 
rect 78 477 81 480 
rect 78 480 81 483 
rect 78 483 81 486 
rect 78 486 81 489 
rect 78 489 81 492 
rect 78 492 81 495 
rect 78 495 81 498 
rect 78 498 81 501 
rect 78 501 81 504 
rect 78 504 81 507 
rect 78 507 81 510 
rect 81 0 84 3 
rect 81 3 84 6 
rect 81 6 84 9 
rect 81 9 84 12 
rect 81 12 84 15 
rect 81 15 84 18 
rect 81 18 84 21 
rect 81 21 84 24 
rect 81 24 84 27 
rect 81 27 84 30 
rect 81 30 84 33 
rect 81 33 84 36 
rect 81 36 84 39 
rect 81 39 84 42 
rect 81 42 84 45 
rect 81 45 84 48 
rect 81 48 84 51 
rect 81 51 84 54 
rect 81 54 84 57 
rect 81 57 84 60 
rect 81 60 84 63 
rect 81 63 84 66 
rect 81 66 84 69 
rect 81 69 84 72 
rect 81 72 84 75 
rect 81 75 84 78 
rect 81 78 84 81 
rect 81 81 84 84 
rect 81 84 84 87 
rect 81 87 84 90 
rect 81 90 84 93 
rect 81 93 84 96 
rect 81 96 84 99 
rect 81 99 84 102 
rect 81 102 84 105 
rect 81 105 84 108 
rect 81 108 84 111 
rect 81 111 84 114 
rect 81 114 84 117 
rect 81 117 84 120 
rect 81 120 84 123 
rect 81 123 84 126 
rect 81 126 84 129 
rect 81 129 84 132 
rect 81 132 84 135 
rect 81 135 84 138 
rect 81 138 84 141 
rect 81 141 84 144 
rect 81 144 84 147 
rect 81 147 84 150 
rect 81 150 84 153 
rect 81 153 84 156 
rect 81 156 84 159 
rect 81 159 84 162 
rect 81 162 84 165 
rect 81 165 84 168 
rect 81 168 84 171 
rect 81 171 84 174 
rect 81 174 84 177 
rect 81 177 84 180 
rect 81 180 84 183 
rect 81 183 84 186 
rect 81 186 84 189 
rect 81 189 84 192 
rect 81 192 84 195 
rect 81 195 84 198 
rect 81 198 84 201 
rect 81 201 84 204 
rect 81 204 84 207 
rect 81 207 84 210 
rect 81 210 84 213 
rect 81 213 84 216 
rect 81 216 84 219 
rect 81 219 84 222 
rect 81 222 84 225 
rect 81 225 84 228 
rect 81 228 84 231 
rect 81 231 84 234 
rect 81 234 84 237 
rect 81 237 84 240 
rect 81 240 84 243 
rect 81 243 84 246 
rect 81 246 84 249 
rect 81 249 84 252 
rect 81 252 84 255 
rect 81 255 84 258 
rect 81 258 84 261 
rect 81 261 84 264 
rect 81 264 84 267 
rect 81 267 84 270 
rect 81 270 84 273 
rect 81 273 84 276 
rect 81 276 84 279 
rect 81 279 84 282 
rect 81 282 84 285 
rect 81 285 84 288 
rect 81 288 84 291 
rect 81 291 84 294 
rect 81 294 84 297 
rect 81 297 84 300 
rect 81 300 84 303 
rect 81 303 84 306 
rect 81 306 84 309 
rect 81 309 84 312 
rect 81 312 84 315 
rect 81 315 84 318 
rect 81 318 84 321 
rect 81 321 84 324 
rect 81 324 84 327 
rect 81 327 84 330 
rect 81 330 84 333 
rect 81 333 84 336 
rect 81 336 84 339 
rect 81 339 84 342 
rect 81 342 84 345 
rect 81 345 84 348 
rect 81 348 84 351 
rect 81 351 84 354 
rect 81 354 84 357 
rect 81 357 84 360 
rect 81 360 84 363 
rect 81 363 84 366 
rect 81 366 84 369 
rect 81 369 84 372 
rect 81 372 84 375 
rect 81 375 84 378 
rect 81 378 84 381 
rect 81 381 84 384 
rect 81 384 84 387 
rect 81 387 84 390 
rect 81 390 84 393 
rect 81 393 84 396 
rect 81 396 84 399 
rect 81 399 84 402 
rect 81 402 84 405 
rect 81 405 84 408 
rect 81 408 84 411 
rect 81 411 84 414 
rect 81 414 84 417 
rect 81 417 84 420 
rect 81 420 84 423 
rect 81 423 84 426 
rect 81 426 84 429 
rect 81 429 84 432 
rect 81 432 84 435 
rect 81 435 84 438 
rect 81 438 84 441 
rect 81 441 84 444 
rect 81 444 84 447 
rect 81 447 84 450 
rect 81 450 84 453 
rect 81 453 84 456 
rect 81 456 84 459 
rect 81 459 84 462 
rect 81 462 84 465 
rect 81 465 84 468 
rect 81 468 84 471 
rect 81 471 84 474 
rect 81 474 84 477 
rect 81 477 84 480 
rect 81 480 84 483 
rect 81 483 84 486 
rect 81 486 84 489 
rect 81 489 84 492 
rect 81 492 84 495 
rect 81 495 84 498 
rect 81 498 84 501 
rect 81 501 84 504 
rect 81 504 84 507 
rect 81 507 84 510 
rect 84 0 87 3 
rect 84 3 87 6 
rect 84 6 87 9 
rect 84 9 87 12 
rect 84 12 87 15 
rect 84 15 87 18 
rect 84 18 87 21 
rect 84 21 87 24 
rect 84 24 87 27 
rect 84 27 87 30 
rect 84 30 87 33 
rect 84 33 87 36 
rect 84 36 87 39 
rect 84 39 87 42 
rect 84 42 87 45 
rect 84 45 87 48 
rect 84 48 87 51 
rect 84 51 87 54 
rect 84 54 87 57 
rect 84 57 87 60 
rect 84 60 87 63 
rect 84 63 87 66 
rect 84 66 87 69 
rect 84 69 87 72 
rect 84 72 87 75 
rect 84 75 87 78 
rect 84 78 87 81 
rect 84 81 87 84 
rect 84 84 87 87 
rect 84 87 87 90 
rect 84 90 87 93 
rect 84 93 87 96 
rect 84 96 87 99 
rect 84 99 87 102 
rect 84 102 87 105 
rect 84 105 87 108 
rect 84 108 87 111 
rect 84 111 87 114 
rect 84 114 87 117 
rect 84 117 87 120 
rect 84 120 87 123 
rect 84 123 87 126 
rect 84 126 87 129 
rect 84 129 87 132 
rect 84 132 87 135 
rect 84 135 87 138 
rect 84 138 87 141 
rect 84 141 87 144 
rect 84 144 87 147 
rect 84 147 87 150 
rect 84 150 87 153 
rect 84 153 87 156 
rect 84 156 87 159 
rect 84 159 87 162 
rect 84 162 87 165 
rect 84 165 87 168 
rect 84 168 87 171 
rect 84 171 87 174 
rect 84 174 87 177 
rect 84 177 87 180 
rect 84 180 87 183 
rect 84 183 87 186 
rect 84 186 87 189 
rect 84 189 87 192 
rect 84 192 87 195 
rect 84 195 87 198 
rect 84 198 87 201 
rect 84 201 87 204 
rect 84 204 87 207 
rect 84 207 87 210 
rect 84 210 87 213 
rect 84 213 87 216 
rect 84 216 87 219 
rect 84 219 87 222 
rect 84 222 87 225 
rect 84 225 87 228 
rect 84 228 87 231 
rect 84 231 87 234 
rect 84 234 87 237 
rect 84 237 87 240 
rect 84 240 87 243 
rect 84 243 87 246 
rect 84 246 87 249 
rect 84 249 87 252 
rect 84 252 87 255 
rect 84 255 87 258 
rect 84 258 87 261 
rect 84 261 87 264 
rect 84 264 87 267 
rect 84 267 87 270 
rect 84 270 87 273 
rect 84 273 87 276 
rect 84 276 87 279 
rect 84 279 87 282 
rect 84 282 87 285 
rect 84 285 87 288 
rect 84 288 87 291 
rect 84 291 87 294 
rect 84 294 87 297 
rect 84 297 87 300 
rect 84 300 87 303 
rect 84 303 87 306 
rect 84 306 87 309 
rect 84 309 87 312 
rect 84 312 87 315 
rect 84 315 87 318 
rect 84 318 87 321 
rect 84 321 87 324 
rect 84 324 87 327 
rect 84 327 87 330 
rect 84 330 87 333 
rect 84 333 87 336 
rect 84 336 87 339 
rect 84 339 87 342 
rect 84 342 87 345 
rect 84 345 87 348 
rect 84 348 87 351 
rect 84 351 87 354 
rect 84 354 87 357 
rect 84 357 87 360 
rect 84 360 87 363 
rect 84 363 87 366 
rect 84 366 87 369 
rect 84 369 87 372 
rect 84 372 87 375 
rect 84 375 87 378 
rect 84 378 87 381 
rect 84 381 87 384 
rect 84 384 87 387 
rect 84 387 87 390 
rect 84 390 87 393 
rect 84 393 87 396 
rect 84 396 87 399 
rect 84 399 87 402 
rect 84 402 87 405 
rect 84 405 87 408 
rect 84 408 87 411 
rect 84 411 87 414 
rect 84 414 87 417 
rect 84 417 87 420 
rect 84 420 87 423 
rect 84 423 87 426 
rect 84 426 87 429 
rect 84 429 87 432 
rect 84 432 87 435 
rect 84 435 87 438 
rect 84 438 87 441 
rect 84 441 87 444 
rect 84 444 87 447 
rect 84 447 87 450 
rect 84 450 87 453 
rect 84 453 87 456 
rect 84 456 87 459 
rect 84 459 87 462 
rect 84 462 87 465 
rect 84 465 87 468 
rect 84 468 87 471 
rect 84 471 87 474 
rect 84 474 87 477 
rect 84 477 87 480 
rect 84 480 87 483 
rect 84 483 87 486 
rect 84 486 87 489 
rect 84 489 87 492 
rect 84 492 87 495 
rect 84 495 87 498 
rect 84 498 87 501 
rect 84 501 87 504 
rect 84 504 87 507 
rect 84 507 87 510 
rect 87 0 90 3 
rect 87 3 90 6 
rect 87 6 90 9 
rect 87 9 90 12 
rect 87 12 90 15 
rect 87 15 90 18 
rect 87 18 90 21 
rect 87 21 90 24 
rect 87 24 90 27 
rect 87 27 90 30 
rect 87 30 90 33 
rect 87 33 90 36 
rect 87 36 90 39 
rect 87 39 90 42 
rect 87 42 90 45 
rect 87 45 90 48 
rect 87 48 90 51 
rect 87 51 90 54 
rect 87 54 90 57 
rect 87 57 90 60 
rect 87 60 90 63 
rect 87 63 90 66 
rect 87 66 90 69 
rect 87 69 90 72 
rect 87 72 90 75 
rect 87 75 90 78 
rect 87 78 90 81 
rect 87 81 90 84 
rect 87 84 90 87 
rect 87 87 90 90 
rect 87 90 90 93 
rect 87 93 90 96 
rect 87 96 90 99 
rect 87 99 90 102 
rect 87 102 90 105 
rect 87 105 90 108 
rect 87 108 90 111 
rect 87 111 90 114 
rect 87 114 90 117 
rect 87 117 90 120 
rect 87 120 90 123 
rect 87 123 90 126 
rect 87 126 90 129 
rect 87 129 90 132 
rect 87 132 90 135 
rect 87 135 90 138 
rect 87 138 90 141 
rect 87 141 90 144 
rect 87 144 90 147 
rect 87 147 90 150 
rect 87 150 90 153 
rect 87 153 90 156 
rect 87 156 90 159 
rect 87 159 90 162 
rect 87 162 90 165 
rect 87 165 90 168 
rect 87 168 90 171 
rect 87 171 90 174 
rect 87 174 90 177 
rect 87 177 90 180 
rect 87 180 90 183 
rect 87 183 90 186 
rect 87 186 90 189 
rect 87 189 90 192 
rect 87 192 90 195 
rect 87 195 90 198 
rect 87 198 90 201 
rect 87 201 90 204 
rect 87 204 90 207 
rect 87 207 90 210 
rect 87 210 90 213 
rect 87 213 90 216 
rect 87 216 90 219 
rect 87 219 90 222 
rect 87 222 90 225 
rect 87 225 90 228 
rect 87 228 90 231 
rect 87 231 90 234 
rect 87 234 90 237 
rect 87 237 90 240 
rect 87 240 90 243 
rect 87 243 90 246 
rect 87 246 90 249 
rect 87 249 90 252 
rect 87 252 90 255 
rect 87 255 90 258 
rect 87 258 90 261 
rect 87 261 90 264 
rect 87 264 90 267 
rect 87 267 90 270 
rect 87 270 90 273 
rect 87 273 90 276 
rect 87 276 90 279 
rect 87 279 90 282 
rect 87 282 90 285 
rect 87 285 90 288 
rect 87 288 90 291 
rect 87 291 90 294 
rect 87 294 90 297 
rect 87 297 90 300 
rect 87 300 90 303 
rect 87 303 90 306 
rect 87 306 90 309 
rect 87 309 90 312 
rect 87 312 90 315 
rect 87 315 90 318 
rect 87 318 90 321 
rect 87 321 90 324 
rect 87 324 90 327 
rect 87 327 90 330 
rect 87 330 90 333 
rect 87 333 90 336 
rect 87 336 90 339 
rect 87 339 90 342 
rect 87 342 90 345 
rect 87 345 90 348 
rect 87 348 90 351 
rect 87 351 90 354 
rect 87 354 90 357 
rect 87 357 90 360 
rect 87 360 90 363 
rect 87 363 90 366 
rect 87 366 90 369 
rect 87 369 90 372 
rect 87 372 90 375 
rect 87 375 90 378 
rect 87 378 90 381 
rect 87 381 90 384 
rect 87 384 90 387 
rect 87 387 90 390 
rect 87 390 90 393 
rect 87 393 90 396 
rect 87 396 90 399 
rect 87 399 90 402 
rect 87 402 90 405 
rect 87 405 90 408 
rect 87 408 90 411 
rect 87 411 90 414 
rect 87 414 90 417 
rect 87 417 90 420 
rect 87 420 90 423 
rect 87 423 90 426 
rect 87 426 90 429 
rect 87 429 90 432 
rect 87 432 90 435 
rect 87 435 90 438 
rect 87 438 90 441 
rect 87 441 90 444 
rect 87 444 90 447 
rect 87 447 90 450 
rect 87 450 90 453 
rect 87 453 90 456 
rect 87 456 90 459 
rect 87 459 90 462 
rect 87 462 90 465 
rect 87 465 90 468 
rect 87 468 90 471 
rect 87 471 90 474 
rect 87 474 90 477 
rect 87 477 90 480 
rect 87 480 90 483 
rect 87 483 90 486 
rect 87 486 90 489 
rect 87 489 90 492 
rect 87 492 90 495 
rect 87 495 90 498 
rect 87 498 90 501 
rect 87 501 90 504 
rect 87 504 90 507 
rect 87 507 90 510 
rect 90 0 93 3 
rect 90 3 93 6 
rect 90 6 93 9 
rect 90 9 93 12 
rect 90 12 93 15 
rect 90 15 93 18 
rect 90 18 93 21 
rect 90 21 93 24 
rect 90 24 93 27 
rect 90 27 93 30 
rect 90 30 93 33 
rect 90 33 93 36 
rect 90 36 93 39 
rect 90 39 93 42 
rect 90 42 93 45 
rect 90 45 93 48 
rect 90 48 93 51 
rect 90 51 93 54 
rect 90 54 93 57 
rect 90 57 93 60 
rect 90 60 93 63 
rect 90 63 93 66 
rect 90 66 93 69 
rect 90 69 93 72 
rect 90 72 93 75 
rect 90 75 93 78 
rect 90 78 93 81 
rect 90 81 93 84 
rect 90 84 93 87 
rect 90 87 93 90 
rect 90 90 93 93 
rect 90 93 93 96 
rect 90 96 93 99 
rect 90 99 93 102 
rect 90 102 93 105 
rect 90 105 93 108 
rect 90 108 93 111 
rect 90 111 93 114 
rect 90 114 93 117 
rect 90 117 93 120 
rect 90 120 93 123 
rect 90 123 93 126 
rect 90 126 93 129 
rect 90 129 93 132 
rect 90 132 93 135 
rect 90 135 93 138 
rect 90 138 93 141 
rect 90 141 93 144 
rect 90 144 93 147 
rect 90 147 93 150 
rect 90 150 93 153 
rect 90 153 93 156 
rect 90 156 93 159 
rect 90 159 93 162 
rect 90 162 93 165 
rect 90 165 93 168 
rect 90 168 93 171 
rect 90 171 93 174 
rect 90 174 93 177 
rect 90 177 93 180 
rect 90 180 93 183 
rect 90 183 93 186 
rect 90 186 93 189 
rect 90 189 93 192 
rect 90 192 93 195 
rect 90 195 93 198 
rect 90 198 93 201 
rect 90 201 93 204 
rect 90 204 93 207 
rect 90 207 93 210 
rect 90 210 93 213 
rect 90 213 93 216 
rect 90 216 93 219 
rect 90 219 93 222 
rect 90 222 93 225 
rect 90 225 93 228 
rect 90 228 93 231 
rect 90 231 93 234 
rect 90 234 93 237 
rect 90 237 93 240 
rect 90 240 93 243 
rect 90 243 93 246 
rect 90 246 93 249 
rect 90 249 93 252 
rect 90 252 93 255 
rect 90 255 93 258 
rect 90 258 93 261 
rect 90 261 93 264 
rect 90 264 93 267 
rect 90 267 93 270 
rect 90 270 93 273 
rect 90 273 93 276 
rect 90 276 93 279 
rect 90 279 93 282 
rect 90 282 93 285 
rect 90 285 93 288 
rect 90 288 93 291 
rect 90 291 93 294 
rect 90 294 93 297 
rect 90 297 93 300 
rect 90 300 93 303 
rect 90 303 93 306 
rect 90 306 93 309 
rect 90 309 93 312 
rect 90 312 93 315 
rect 90 315 93 318 
rect 90 318 93 321 
rect 90 321 93 324 
rect 90 324 93 327 
rect 90 327 93 330 
rect 90 330 93 333 
rect 90 333 93 336 
rect 90 336 93 339 
rect 90 339 93 342 
rect 90 342 93 345 
rect 90 345 93 348 
rect 90 348 93 351 
rect 90 351 93 354 
rect 90 354 93 357 
rect 90 357 93 360 
rect 90 360 93 363 
rect 90 363 93 366 
rect 90 366 93 369 
rect 90 369 93 372 
rect 90 372 93 375 
rect 90 375 93 378 
rect 90 378 93 381 
rect 90 381 93 384 
rect 90 384 93 387 
rect 90 387 93 390 
rect 90 390 93 393 
rect 90 393 93 396 
rect 90 396 93 399 
rect 90 399 93 402 
rect 90 402 93 405 
rect 90 405 93 408 
rect 90 408 93 411 
rect 90 411 93 414 
rect 90 414 93 417 
rect 90 417 93 420 
rect 90 420 93 423 
rect 90 423 93 426 
rect 90 426 93 429 
rect 90 429 93 432 
rect 90 432 93 435 
rect 90 435 93 438 
rect 90 438 93 441 
rect 90 441 93 444 
rect 90 444 93 447 
rect 90 447 93 450 
rect 90 450 93 453 
rect 90 453 93 456 
rect 90 456 93 459 
rect 90 459 93 462 
rect 90 462 93 465 
rect 90 465 93 468 
rect 90 468 93 471 
rect 90 471 93 474 
rect 90 474 93 477 
rect 90 477 93 480 
rect 90 480 93 483 
rect 90 483 93 486 
rect 90 486 93 489 
rect 90 489 93 492 
rect 90 492 93 495 
rect 90 495 93 498 
rect 90 498 93 501 
rect 90 501 93 504 
rect 90 504 93 507 
rect 90 507 93 510 
rect 93 0 96 3 
rect 93 3 96 6 
rect 93 6 96 9 
rect 93 9 96 12 
rect 93 12 96 15 
rect 93 15 96 18 
rect 93 18 96 21 
rect 93 21 96 24 
rect 93 24 96 27 
rect 93 27 96 30 
rect 93 30 96 33 
rect 93 33 96 36 
rect 93 36 96 39 
rect 93 39 96 42 
rect 93 42 96 45 
rect 93 45 96 48 
rect 93 48 96 51 
rect 93 51 96 54 
rect 93 54 96 57 
rect 93 57 96 60 
rect 93 60 96 63 
rect 93 63 96 66 
rect 93 66 96 69 
rect 93 69 96 72 
rect 93 72 96 75 
rect 93 75 96 78 
rect 93 78 96 81 
rect 93 81 96 84 
rect 93 84 96 87 
rect 93 87 96 90 
rect 93 90 96 93 
rect 93 93 96 96 
rect 93 96 96 99 
rect 93 99 96 102 
rect 93 102 96 105 
rect 93 105 96 108 
rect 93 108 96 111 
rect 93 111 96 114 
rect 93 114 96 117 
rect 93 117 96 120 
rect 93 120 96 123 
rect 93 123 96 126 
rect 93 126 96 129 
rect 93 129 96 132 
rect 93 132 96 135 
rect 93 135 96 138 
rect 93 138 96 141 
rect 93 141 96 144 
rect 93 144 96 147 
rect 93 147 96 150 
rect 93 150 96 153 
rect 93 153 96 156 
rect 93 156 96 159 
rect 93 159 96 162 
rect 93 162 96 165 
rect 93 165 96 168 
rect 93 168 96 171 
rect 93 171 96 174 
rect 93 174 96 177 
rect 93 177 96 180 
rect 93 180 96 183 
rect 93 183 96 186 
rect 93 186 96 189 
rect 93 189 96 192 
rect 93 192 96 195 
rect 93 195 96 198 
rect 93 198 96 201 
rect 93 201 96 204 
rect 93 204 96 207 
rect 93 207 96 210 
rect 93 210 96 213 
rect 93 213 96 216 
rect 93 216 96 219 
rect 93 219 96 222 
rect 93 222 96 225 
rect 93 225 96 228 
rect 93 228 96 231 
rect 93 231 96 234 
rect 93 234 96 237 
rect 93 237 96 240 
rect 93 240 96 243 
rect 93 243 96 246 
rect 93 246 96 249 
rect 93 249 96 252 
rect 93 252 96 255 
rect 93 255 96 258 
rect 93 258 96 261 
rect 93 261 96 264 
rect 93 264 96 267 
rect 93 267 96 270 
rect 93 270 96 273 
rect 93 273 96 276 
rect 93 276 96 279 
rect 93 279 96 282 
rect 93 282 96 285 
rect 93 285 96 288 
rect 93 288 96 291 
rect 93 291 96 294 
rect 93 294 96 297 
rect 93 297 96 300 
rect 93 300 96 303 
rect 93 303 96 306 
rect 93 306 96 309 
rect 93 309 96 312 
rect 93 312 96 315 
rect 93 315 96 318 
rect 93 318 96 321 
rect 93 321 96 324 
rect 93 324 96 327 
rect 93 327 96 330 
rect 93 330 96 333 
rect 93 333 96 336 
rect 93 336 96 339 
rect 93 339 96 342 
rect 93 342 96 345 
rect 93 345 96 348 
rect 93 348 96 351 
rect 93 351 96 354 
rect 93 354 96 357 
rect 93 357 96 360 
rect 93 360 96 363 
rect 93 363 96 366 
rect 93 366 96 369 
rect 93 369 96 372 
rect 93 372 96 375 
rect 93 375 96 378 
rect 93 378 96 381 
rect 93 381 96 384 
rect 93 384 96 387 
rect 93 387 96 390 
rect 93 390 96 393 
rect 93 393 96 396 
rect 93 396 96 399 
rect 93 399 96 402 
rect 93 402 96 405 
rect 93 405 96 408 
rect 93 408 96 411 
rect 93 411 96 414 
rect 93 414 96 417 
rect 93 417 96 420 
rect 93 420 96 423 
rect 93 423 96 426 
rect 93 426 96 429 
rect 93 429 96 432 
rect 93 432 96 435 
rect 93 435 96 438 
rect 93 438 96 441 
rect 93 441 96 444 
rect 93 444 96 447 
rect 93 447 96 450 
rect 93 450 96 453 
rect 93 453 96 456 
rect 93 456 96 459 
rect 93 459 96 462 
rect 93 462 96 465 
rect 93 465 96 468 
rect 93 468 96 471 
rect 93 471 96 474 
rect 93 474 96 477 
rect 93 477 96 480 
rect 93 480 96 483 
rect 93 483 96 486 
rect 93 486 96 489 
rect 93 489 96 492 
rect 93 492 96 495 
rect 93 495 96 498 
rect 93 498 96 501 
rect 93 501 96 504 
rect 93 504 96 507 
rect 93 507 96 510 
rect 96 0 99 3 
rect 96 3 99 6 
rect 96 6 99 9 
rect 96 9 99 12 
rect 96 12 99 15 
rect 96 15 99 18 
rect 96 18 99 21 
rect 96 21 99 24 
rect 96 24 99 27 
rect 96 27 99 30 
rect 96 30 99 33 
rect 96 33 99 36 
rect 96 36 99 39 
rect 96 39 99 42 
rect 96 42 99 45 
rect 96 45 99 48 
rect 96 48 99 51 
rect 96 51 99 54 
rect 96 54 99 57 
rect 96 57 99 60 
rect 96 60 99 63 
rect 96 63 99 66 
rect 96 66 99 69 
rect 96 69 99 72 
rect 96 72 99 75 
rect 96 75 99 78 
rect 96 78 99 81 
rect 96 81 99 84 
rect 96 84 99 87 
rect 96 87 99 90 
rect 96 90 99 93 
rect 96 93 99 96 
rect 96 96 99 99 
rect 96 99 99 102 
rect 96 102 99 105 
rect 96 105 99 108 
rect 96 108 99 111 
rect 96 111 99 114 
rect 96 114 99 117 
rect 96 117 99 120 
rect 96 120 99 123 
rect 96 123 99 126 
rect 96 126 99 129 
rect 96 129 99 132 
rect 96 132 99 135 
rect 96 135 99 138 
rect 96 138 99 141 
rect 96 141 99 144 
rect 96 144 99 147 
rect 96 147 99 150 
rect 96 150 99 153 
rect 96 153 99 156 
rect 96 156 99 159 
rect 96 159 99 162 
rect 96 162 99 165 
rect 96 165 99 168 
rect 96 168 99 171 
rect 96 171 99 174 
rect 96 174 99 177 
rect 96 177 99 180 
rect 96 180 99 183 
rect 96 183 99 186 
rect 96 186 99 189 
rect 96 189 99 192 
rect 96 192 99 195 
rect 96 195 99 198 
rect 96 198 99 201 
rect 96 201 99 204 
rect 96 204 99 207 
rect 96 207 99 210 
rect 96 210 99 213 
rect 96 213 99 216 
rect 96 216 99 219 
rect 96 219 99 222 
rect 96 222 99 225 
rect 96 225 99 228 
rect 96 228 99 231 
rect 96 231 99 234 
rect 96 234 99 237 
rect 96 237 99 240 
rect 96 240 99 243 
rect 96 243 99 246 
rect 96 246 99 249 
rect 96 249 99 252 
rect 96 252 99 255 
rect 96 255 99 258 
rect 96 258 99 261 
rect 96 261 99 264 
rect 96 264 99 267 
rect 96 267 99 270 
rect 96 270 99 273 
rect 96 273 99 276 
rect 96 276 99 279 
rect 96 279 99 282 
rect 96 282 99 285 
rect 96 285 99 288 
rect 96 288 99 291 
rect 96 291 99 294 
rect 96 294 99 297 
rect 96 297 99 300 
rect 96 300 99 303 
rect 96 303 99 306 
rect 96 306 99 309 
rect 96 309 99 312 
rect 96 312 99 315 
rect 96 315 99 318 
rect 96 318 99 321 
rect 96 321 99 324 
rect 96 324 99 327 
rect 96 327 99 330 
rect 96 330 99 333 
rect 96 333 99 336 
rect 96 336 99 339 
rect 96 339 99 342 
rect 96 342 99 345 
rect 96 345 99 348 
rect 96 348 99 351 
rect 96 351 99 354 
rect 96 354 99 357 
rect 96 357 99 360 
rect 96 360 99 363 
rect 96 363 99 366 
rect 96 366 99 369 
rect 96 369 99 372 
rect 96 372 99 375 
rect 96 375 99 378 
rect 96 378 99 381 
rect 96 381 99 384 
rect 96 384 99 387 
rect 96 387 99 390 
rect 96 390 99 393 
rect 96 393 99 396 
rect 96 396 99 399 
rect 96 399 99 402 
rect 96 402 99 405 
rect 96 405 99 408 
rect 96 408 99 411 
rect 96 411 99 414 
rect 96 414 99 417 
rect 96 417 99 420 
rect 96 420 99 423 
rect 96 423 99 426 
rect 96 426 99 429 
rect 96 429 99 432 
rect 96 432 99 435 
rect 96 435 99 438 
rect 96 438 99 441 
rect 96 441 99 444 
rect 96 444 99 447 
rect 96 447 99 450 
rect 96 450 99 453 
rect 96 453 99 456 
rect 96 456 99 459 
rect 96 459 99 462 
rect 96 462 99 465 
rect 96 465 99 468 
rect 96 468 99 471 
rect 96 471 99 474 
rect 96 474 99 477 
rect 96 477 99 480 
rect 96 480 99 483 
rect 96 483 99 486 
rect 96 486 99 489 
rect 96 489 99 492 
rect 96 492 99 495 
rect 96 495 99 498 
rect 96 498 99 501 
rect 96 501 99 504 
rect 96 504 99 507 
rect 96 507 99 510 
rect 99 0 102 3 
rect 99 3 102 6 
rect 99 6 102 9 
rect 99 9 102 12 
rect 99 12 102 15 
rect 99 15 102 18 
rect 99 18 102 21 
rect 99 21 102 24 
rect 99 24 102 27 
rect 99 27 102 30 
rect 99 30 102 33 
rect 99 33 102 36 
rect 99 36 102 39 
rect 99 39 102 42 
rect 99 42 102 45 
rect 99 45 102 48 
rect 99 48 102 51 
rect 99 51 102 54 
rect 99 54 102 57 
rect 99 57 102 60 
rect 99 60 102 63 
rect 99 63 102 66 
rect 99 66 102 69 
rect 99 69 102 72 
rect 99 72 102 75 
rect 99 75 102 78 
rect 99 78 102 81 
rect 99 81 102 84 
rect 99 84 102 87 
rect 99 87 102 90 
rect 99 90 102 93 
rect 99 93 102 96 
rect 99 96 102 99 
rect 99 99 102 102 
rect 99 102 102 105 
rect 99 105 102 108 
rect 99 108 102 111 
rect 99 111 102 114 
rect 99 114 102 117 
rect 99 117 102 120 
rect 99 120 102 123 
rect 99 123 102 126 
rect 99 126 102 129 
rect 99 129 102 132 
rect 99 132 102 135 
rect 99 135 102 138 
rect 99 138 102 141 
rect 99 141 102 144 
rect 99 144 102 147 
rect 99 147 102 150 
rect 99 150 102 153 
rect 99 153 102 156 
rect 99 156 102 159 
rect 99 159 102 162 
rect 99 162 102 165 
rect 99 165 102 168 
rect 99 168 102 171 
rect 99 171 102 174 
rect 99 174 102 177 
rect 99 177 102 180 
rect 99 180 102 183 
rect 99 183 102 186 
rect 99 186 102 189 
rect 99 189 102 192 
rect 99 192 102 195 
rect 99 195 102 198 
rect 99 198 102 201 
rect 99 201 102 204 
rect 99 204 102 207 
rect 99 207 102 210 
rect 99 210 102 213 
rect 99 213 102 216 
rect 99 216 102 219 
rect 99 219 102 222 
rect 99 222 102 225 
rect 99 225 102 228 
rect 99 228 102 231 
rect 99 231 102 234 
rect 99 234 102 237 
rect 99 237 102 240 
rect 99 240 102 243 
rect 99 243 102 246 
rect 99 246 102 249 
rect 99 249 102 252 
rect 99 252 102 255 
rect 99 255 102 258 
rect 99 258 102 261 
rect 99 261 102 264 
rect 99 264 102 267 
rect 99 267 102 270 
rect 99 270 102 273 
rect 99 273 102 276 
rect 99 276 102 279 
rect 99 279 102 282 
rect 99 282 102 285 
rect 99 285 102 288 
rect 99 288 102 291 
rect 99 291 102 294 
rect 99 294 102 297 
rect 99 297 102 300 
rect 99 300 102 303 
rect 99 303 102 306 
rect 99 306 102 309 
rect 99 309 102 312 
rect 99 312 102 315 
rect 99 315 102 318 
rect 99 318 102 321 
rect 99 321 102 324 
rect 99 324 102 327 
rect 99 327 102 330 
rect 99 330 102 333 
rect 99 333 102 336 
rect 99 336 102 339 
rect 99 339 102 342 
rect 99 342 102 345 
rect 99 345 102 348 
rect 99 348 102 351 
rect 99 351 102 354 
rect 99 354 102 357 
rect 99 357 102 360 
rect 99 360 102 363 
rect 99 363 102 366 
rect 99 366 102 369 
rect 99 369 102 372 
rect 99 372 102 375 
rect 99 375 102 378 
rect 99 378 102 381 
rect 99 381 102 384 
rect 99 384 102 387 
rect 99 387 102 390 
rect 99 390 102 393 
rect 99 393 102 396 
rect 99 396 102 399 
rect 99 399 102 402 
rect 99 402 102 405 
rect 99 405 102 408 
rect 99 408 102 411 
rect 99 411 102 414 
rect 99 414 102 417 
rect 99 417 102 420 
rect 99 420 102 423 
rect 99 423 102 426 
rect 99 426 102 429 
rect 99 429 102 432 
rect 99 432 102 435 
rect 99 435 102 438 
rect 99 438 102 441 
rect 99 441 102 444 
rect 99 444 102 447 
rect 99 447 102 450 
rect 99 450 102 453 
rect 99 453 102 456 
rect 99 456 102 459 
rect 99 459 102 462 
rect 99 462 102 465 
rect 99 465 102 468 
rect 99 468 102 471 
rect 99 471 102 474 
rect 99 474 102 477 
rect 99 477 102 480 
rect 99 480 102 483 
rect 99 483 102 486 
rect 99 486 102 489 
rect 99 489 102 492 
rect 99 492 102 495 
rect 99 495 102 498 
rect 99 498 102 501 
rect 99 501 102 504 
rect 99 504 102 507 
rect 99 507 102 510 
rect 102 0 105 3 
rect 102 3 105 6 
rect 102 6 105 9 
rect 102 9 105 12 
rect 102 12 105 15 
rect 102 15 105 18 
rect 102 18 105 21 
rect 102 21 105 24 
rect 102 24 105 27 
rect 102 27 105 30 
rect 102 30 105 33 
rect 102 33 105 36 
rect 102 36 105 39 
rect 102 39 105 42 
rect 102 42 105 45 
rect 102 45 105 48 
rect 102 48 105 51 
rect 102 51 105 54 
rect 102 54 105 57 
rect 102 57 105 60 
rect 102 60 105 63 
rect 102 63 105 66 
rect 102 66 105 69 
rect 102 69 105 72 
rect 102 72 105 75 
rect 102 75 105 78 
rect 102 78 105 81 
rect 102 81 105 84 
rect 102 84 105 87 
rect 102 87 105 90 
rect 102 90 105 93 
rect 102 93 105 96 
rect 102 96 105 99 
rect 102 99 105 102 
rect 102 102 105 105 
rect 102 105 105 108 
rect 102 108 105 111 
rect 102 111 105 114 
rect 102 114 105 117 
rect 102 117 105 120 
rect 102 120 105 123 
rect 102 123 105 126 
rect 102 126 105 129 
rect 102 129 105 132 
rect 102 132 105 135 
rect 102 135 105 138 
rect 102 138 105 141 
rect 102 141 105 144 
rect 102 144 105 147 
rect 102 147 105 150 
rect 102 150 105 153 
rect 102 153 105 156 
rect 102 156 105 159 
rect 102 159 105 162 
rect 102 162 105 165 
rect 102 165 105 168 
rect 102 168 105 171 
rect 102 171 105 174 
rect 102 174 105 177 
rect 102 177 105 180 
rect 102 180 105 183 
rect 102 183 105 186 
rect 102 186 105 189 
rect 102 189 105 192 
rect 102 192 105 195 
rect 102 195 105 198 
rect 102 198 105 201 
rect 102 201 105 204 
rect 102 204 105 207 
rect 102 207 105 210 
rect 102 210 105 213 
rect 102 213 105 216 
rect 102 216 105 219 
rect 102 219 105 222 
rect 102 222 105 225 
rect 102 225 105 228 
rect 102 228 105 231 
rect 102 231 105 234 
rect 102 234 105 237 
rect 102 237 105 240 
rect 102 240 105 243 
rect 102 243 105 246 
rect 102 246 105 249 
rect 102 249 105 252 
rect 102 252 105 255 
rect 102 255 105 258 
rect 102 258 105 261 
rect 102 261 105 264 
rect 102 264 105 267 
rect 102 267 105 270 
rect 102 270 105 273 
rect 102 273 105 276 
rect 102 276 105 279 
rect 102 279 105 282 
rect 102 282 105 285 
rect 102 285 105 288 
rect 102 288 105 291 
rect 102 291 105 294 
rect 102 294 105 297 
rect 102 297 105 300 
rect 102 300 105 303 
rect 102 303 105 306 
rect 102 306 105 309 
rect 102 309 105 312 
rect 102 312 105 315 
rect 102 315 105 318 
rect 102 318 105 321 
rect 102 321 105 324 
rect 102 324 105 327 
rect 102 327 105 330 
rect 102 330 105 333 
rect 102 333 105 336 
rect 102 336 105 339 
rect 102 339 105 342 
rect 102 342 105 345 
rect 102 345 105 348 
rect 102 348 105 351 
rect 102 351 105 354 
rect 102 354 105 357 
rect 102 357 105 360 
rect 102 360 105 363 
rect 102 363 105 366 
rect 102 366 105 369 
rect 102 369 105 372 
rect 102 372 105 375 
rect 102 375 105 378 
rect 102 378 105 381 
rect 102 381 105 384 
rect 102 384 105 387 
rect 102 387 105 390 
rect 102 390 105 393 
rect 102 393 105 396 
rect 102 396 105 399 
rect 102 399 105 402 
rect 102 402 105 405 
rect 102 405 105 408 
rect 102 408 105 411 
rect 102 411 105 414 
rect 102 414 105 417 
rect 102 417 105 420 
rect 102 420 105 423 
rect 102 423 105 426 
rect 102 426 105 429 
rect 102 429 105 432 
rect 102 432 105 435 
rect 102 435 105 438 
rect 102 438 105 441 
rect 102 441 105 444 
rect 102 444 105 447 
rect 102 447 105 450 
rect 102 450 105 453 
rect 102 453 105 456 
rect 102 456 105 459 
rect 102 459 105 462 
rect 102 462 105 465 
rect 102 465 105 468 
rect 102 468 105 471 
rect 102 471 105 474 
rect 102 474 105 477 
rect 102 477 105 480 
rect 102 480 105 483 
rect 102 483 105 486 
rect 102 486 105 489 
rect 102 489 105 492 
rect 102 492 105 495 
rect 102 495 105 498 
rect 102 498 105 501 
rect 102 501 105 504 
rect 102 504 105 507 
rect 102 507 105 510 
rect 105 0 108 3 
rect 105 3 108 6 
rect 105 6 108 9 
rect 105 9 108 12 
rect 105 12 108 15 
rect 105 15 108 18 
rect 105 18 108 21 
rect 105 21 108 24 
rect 105 24 108 27 
rect 105 27 108 30 
rect 105 30 108 33 
rect 105 33 108 36 
rect 105 36 108 39 
rect 105 39 108 42 
rect 105 42 108 45 
rect 105 45 108 48 
rect 105 48 108 51 
rect 105 51 108 54 
rect 105 54 108 57 
rect 105 57 108 60 
rect 105 60 108 63 
rect 105 63 108 66 
rect 105 66 108 69 
rect 105 69 108 72 
rect 105 72 108 75 
rect 105 75 108 78 
rect 105 78 108 81 
rect 105 81 108 84 
rect 105 84 108 87 
rect 105 87 108 90 
rect 105 90 108 93 
rect 105 93 108 96 
rect 105 96 108 99 
rect 105 99 108 102 
rect 105 102 108 105 
rect 105 105 108 108 
rect 105 108 108 111 
rect 105 111 108 114 
rect 105 114 108 117 
rect 105 117 108 120 
rect 105 120 108 123 
rect 105 123 108 126 
rect 105 126 108 129 
rect 105 129 108 132 
rect 105 132 108 135 
rect 105 135 108 138 
rect 105 138 108 141 
rect 105 141 108 144 
rect 105 144 108 147 
rect 105 147 108 150 
rect 105 150 108 153 
rect 105 153 108 156 
rect 105 156 108 159 
rect 105 159 108 162 
rect 105 162 108 165 
rect 105 165 108 168 
rect 105 168 108 171 
rect 105 171 108 174 
rect 105 174 108 177 
rect 105 177 108 180 
rect 105 180 108 183 
rect 105 183 108 186 
rect 105 186 108 189 
rect 105 189 108 192 
rect 105 192 108 195 
rect 105 195 108 198 
rect 105 198 108 201 
rect 105 201 108 204 
rect 105 204 108 207 
rect 105 207 108 210 
rect 105 210 108 213 
rect 105 213 108 216 
rect 105 216 108 219 
rect 105 219 108 222 
rect 105 222 108 225 
rect 105 225 108 228 
rect 105 228 108 231 
rect 105 231 108 234 
rect 105 234 108 237 
rect 105 237 108 240 
rect 105 240 108 243 
rect 105 243 108 246 
rect 105 246 108 249 
rect 105 249 108 252 
rect 105 252 108 255 
rect 105 255 108 258 
rect 105 258 108 261 
rect 105 261 108 264 
rect 105 264 108 267 
rect 105 267 108 270 
rect 105 270 108 273 
rect 105 273 108 276 
rect 105 276 108 279 
rect 105 279 108 282 
rect 105 282 108 285 
rect 105 285 108 288 
rect 105 288 108 291 
rect 105 291 108 294 
rect 105 294 108 297 
rect 105 297 108 300 
rect 105 300 108 303 
rect 105 303 108 306 
rect 105 306 108 309 
rect 105 309 108 312 
rect 105 312 108 315 
rect 105 315 108 318 
rect 105 318 108 321 
rect 105 321 108 324 
rect 105 324 108 327 
rect 105 327 108 330 
rect 105 330 108 333 
rect 105 333 108 336 
rect 105 336 108 339 
rect 105 339 108 342 
rect 105 342 108 345 
rect 105 345 108 348 
rect 105 348 108 351 
rect 105 351 108 354 
rect 105 354 108 357 
rect 105 357 108 360 
rect 105 360 108 363 
rect 105 363 108 366 
rect 105 366 108 369 
rect 105 369 108 372 
rect 105 372 108 375 
rect 105 375 108 378 
rect 105 378 108 381 
rect 105 381 108 384 
rect 105 384 108 387 
rect 105 387 108 390 
rect 105 390 108 393 
rect 105 393 108 396 
rect 105 396 108 399 
rect 105 399 108 402 
rect 105 402 108 405 
rect 105 405 108 408 
rect 105 408 108 411 
rect 105 411 108 414 
rect 105 414 108 417 
rect 105 417 108 420 
rect 105 420 108 423 
rect 105 423 108 426 
rect 105 426 108 429 
rect 105 429 108 432 
rect 105 432 108 435 
rect 105 435 108 438 
rect 105 438 108 441 
rect 105 441 108 444 
rect 105 444 108 447 
rect 105 447 108 450 
rect 105 450 108 453 
rect 105 453 108 456 
rect 105 456 108 459 
rect 105 459 108 462 
rect 105 462 108 465 
rect 105 465 108 468 
rect 105 468 108 471 
rect 105 471 108 474 
rect 105 474 108 477 
rect 105 477 108 480 
rect 105 480 108 483 
rect 105 483 108 486 
rect 105 486 108 489 
rect 105 489 108 492 
rect 105 492 108 495 
rect 105 495 108 498 
rect 105 498 108 501 
rect 105 501 108 504 
rect 105 504 108 507 
rect 105 507 108 510 
rect 108 0 111 3 
rect 108 3 111 6 
rect 108 6 111 9 
rect 108 9 111 12 
rect 108 12 111 15 
rect 108 15 111 18 
rect 108 18 111 21 
rect 108 21 111 24 
rect 108 24 111 27 
rect 108 27 111 30 
rect 108 30 111 33 
rect 108 33 111 36 
rect 108 36 111 39 
rect 108 39 111 42 
rect 108 42 111 45 
rect 108 45 111 48 
rect 108 48 111 51 
rect 108 51 111 54 
rect 108 54 111 57 
rect 108 57 111 60 
rect 108 60 111 63 
rect 108 63 111 66 
rect 108 66 111 69 
rect 108 69 111 72 
rect 108 72 111 75 
rect 108 75 111 78 
rect 108 78 111 81 
rect 108 81 111 84 
rect 108 84 111 87 
rect 108 87 111 90 
rect 108 90 111 93 
rect 108 93 111 96 
rect 108 96 111 99 
rect 108 99 111 102 
rect 108 102 111 105 
rect 108 105 111 108 
rect 108 108 111 111 
rect 108 111 111 114 
rect 108 114 111 117 
rect 108 117 111 120 
rect 108 120 111 123 
rect 108 123 111 126 
rect 108 126 111 129 
rect 108 129 111 132 
rect 108 132 111 135 
rect 108 135 111 138 
rect 108 138 111 141 
rect 108 141 111 144 
rect 108 144 111 147 
rect 108 147 111 150 
rect 108 150 111 153 
rect 108 153 111 156 
rect 108 156 111 159 
rect 108 159 111 162 
rect 108 162 111 165 
rect 108 165 111 168 
rect 108 168 111 171 
rect 108 171 111 174 
rect 108 174 111 177 
rect 108 177 111 180 
rect 108 180 111 183 
rect 108 183 111 186 
rect 108 186 111 189 
rect 108 189 111 192 
rect 108 192 111 195 
rect 108 195 111 198 
rect 108 198 111 201 
rect 108 201 111 204 
rect 108 204 111 207 
rect 108 207 111 210 
rect 108 210 111 213 
rect 108 213 111 216 
rect 108 216 111 219 
rect 108 219 111 222 
rect 108 222 111 225 
rect 108 225 111 228 
rect 108 228 111 231 
rect 108 231 111 234 
rect 108 234 111 237 
rect 108 237 111 240 
rect 108 240 111 243 
rect 108 243 111 246 
rect 108 246 111 249 
rect 108 249 111 252 
rect 108 252 111 255 
rect 108 255 111 258 
rect 108 258 111 261 
rect 108 261 111 264 
rect 108 264 111 267 
rect 108 267 111 270 
rect 108 270 111 273 
rect 108 273 111 276 
rect 108 276 111 279 
rect 108 279 111 282 
rect 108 282 111 285 
rect 108 285 111 288 
rect 108 288 111 291 
rect 108 291 111 294 
rect 108 294 111 297 
rect 108 297 111 300 
rect 108 300 111 303 
rect 108 303 111 306 
rect 108 306 111 309 
rect 108 309 111 312 
rect 108 312 111 315 
rect 108 315 111 318 
rect 108 318 111 321 
rect 108 321 111 324 
rect 108 324 111 327 
rect 108 327 111 330 
rect 108 330 111 333 
rect 108 333 111 336 
rect 108 336 111 339 
rect 108 339 111 342 
rect 108 342 111 345 
rect 108 345 111 348 
rect 108 348 111 351 
rect 108 351 111 354 
rect 108 354 111 357 
rect 108 357 111 360 
rect 108 360 111 363 
rect 108 363 111 366 
rect 108 366 111 369 
rect 108 369 111 372 
rect 108 372 111 375 
rect 108 375 111 378 
rect 108 378 111 381 
rect 108 381 111 384 
rect 108 384 111 387 
rect 108 387 111 390 
rect 108 390 111 393 
rect 108 393 111 396 
rect 108 396 111 399 
rect 108 399 111 402 
rect 108 402 111 405 
rect 108 405 111 408 
rect 108 408 111 411 
rect 108 411 111 414 
rect 108 414 111 417 
rect 108 417 111 420 
rect 108 420 111 423 
rect 108 423 111 426 
rect 108 426 111 429 
rect 108 429 111 432 
rect 108 432 111 435 
rect 108 435 111 438 
rect 108 438 111 441 
rect 108 441 111 444 
rect 108 444 111 447 
rect 108 447 111 450 
rect 108 450 111 453 
rect 108 453 111 456 
rect 108 456 111 459 
rect 108 459 111 462 
rect 108 462 111 465 
rect 108 465 111 468 
rect 108 468 111 471 
rect 108 471 111 474 
rect 108 474 111 477 
rect 108 477 111 480 
rect 108 480 111 483 
rect 108 483 111 486 
rect 108 486 111 489 
rect 108 489 111 492 
rect 108 492 111 495 
rect 108 495 111 498 
rect 108 498 111 501 
rect 108 501 111 504 
rect 108 504 111 507 
rect 108 507 111 510 
rect 111 0 114 3 
rect 111 3 114 6 
rect 111 6 114 9 
rect 111 9 114 12 
rect 111 12 114 15 
rect 111 15 114 18 
rect 111 18 114 21 
rect 111 21 114 24 
rect 111 24 114 27 
rect 111 27 114 30 
rect 111 30 114 33 
rect 111 33 114 36 
rect 111 36 114 39 
rect 111 39 114 42 
rect 111 42 114 45 
rect 111 45 114 48 
rect 111 48 114 51 
rect 111 51 114 54 
rect 111 54 114 57 
rect 111 57 114 60 
rect 111 60 114 63 
rect 111 63 114 66 
rect 111 66 114 69 
rect 111 69 114 72 
rect 111 72 114 75 
rect 111 75 114 78 
rect 111 78 114 81 
rect 111 81 114 84 
rect 111 84 114 87 
rect 111 87 114 90 
rect 111 90 114 93 
rect 111 93 114 96 
rect 111 96 114 99 
rect 111 99 114 102 
rect 111 102 114 105 
rect 111 105 114 108 
rect 111 108 114 111 
rect 111 111 114 114 
rect 111 114 114 117 
rect 111 117 114 120 
rect 111 120 114 123 
rect 111 123 114 126 
rect 111 126 114 129 
rect 111 129 114 132 
rect 111 132 114 135 
rect 111 135 114 138 
rect 111 138 114 141 
rect 111 141 114 144 
rect 111 144 114 147 
rect 111 147 114 150 
rect 111 150 114 153 
rect 111 153 114 156 
rect 111 156 114 159 
rect 111 159 114 162 
rect 111 162 114 165 
rect 111 165 114 168 
rect 111 168 114 171 
rect 111 171 114 174 
rect 111 174 114 177 
rect 111 177 114 180 
rect 111 180 114 183 
rect 111 183 114 186 
rect 111 186 114 189 
rect 111 189 114 192 
rect 111 192 114 195 
rect 111 195 114 198 
rect 111 198 114 201 
rect 111 201 114 204 
rect 111 204 114 207 
rect 111 207 114 210 
rect 111 210 114 213 
rect 111 213 114 216 
rect 111 216 114 219 
rect 111 219 114 222 
rect 111 222 114 225 
rect 111 225 114 228 
rect 111 228 114 231 
rect 111 231 114 234 
rect 111 234 114 237 
rect 111 237 114 240 
rect 111 240 114 243 
rect 111 243 114 246 
rect 111 246 114 249 
rect 111 249 114 252 
rect 111 252 114 255 
rect 111 255 114 258 
rect 111 258 114 261 
rect 111 261 114 264 
rect 111 264 114 267 
rect 111 267 114 270 
rect 111 270 114 273 
rect 111 273 114 276 
rect 111 276 114 279 
rect 111 279 114 282 
rect 111 282 114 285 
rect 111 285 114 288 
rect 111 288 114 291 
rect 111 291 114 294 
rect 111 294 114 297 
rect 111 297 114 300 
rect 111 300 114 303 
rect 111 303 114 306 
rect 111 306 114 309 
rect 111 309 114 312 
rect 111 312 114 315 
rect 111 315 114 318 
rect 111 318 114 321 
rect 111 321 114 324 
rect 111 324 114 327 
rect 111 327 114 330 
rect 111 330 114 333 
rect 111 333 114 336 
rect 111 336 114 339 
rect 111 339 114 342 
rect 111 342 114 345 
rect 111 345 114 348 
rect 111 348 114 351 
rect 111 351 114 354 
rect 111 354 114 357 
rect 111 357 114 360 
rect 111 360 114 363 
rect 111 363 114 366 
rect 111 366 114 369 
rect 111 369 114 372 
rect 111 372 114 375 
rect 111 375 114 378 
rect 111 378 114 381 
rect 111 381 114 384 
rect 111 384 114 387 
rect 111 387 114 390 
rect 111 390 114 393 
rect 111 393 114 396 
rect 111 396 114 399 
rect 111 399 114 402 
rect 111 402 114 405 
rect 111 405 114 408 
rect 111 408 114 411 
rect 111 411 114 414 
rect 111 414 114 417 
rect 111 417 114 420 
rect 111 420 114 423 
rect 111 423 114 426 
rect 111 426 114 429 
rect 111 429 114 432 
rect 111 432 114 435 
rect 111 435 114 438 
rect 111 438 114 441 
rect 111 441 114 444 
rect 111 444 114 447 
rect 111 447 114 450 
rect 111 450 114 453 
rect 111 453 114 456 
rect 111 456 114 459 
rect 111 459 114 462 
rect 111 462 114 465 
rect 111 465 114 468 
rect 111 468 114 471 
rect 111 471 114 474 
rect 111 474 114 477 
rect 111 477 114 480 
rect 111 480 114 483 
rect 111 483 114 486 
rect 111 486 114 489 
rect 111 489 114 492 
rect 111 492 114 495 
rect 111 495 114 498 
rect 111 498 114 501 
rect 111 501 114 504 
rect 111 504 114 507 
rect 111 507 114 510 
rect 114 0 117 3 
rect 114 3 117 6 
rect 114 6 117 9 
rect 114 9 117 12 
rect 114 12 117 15 
rect 114 15 117 18 
rect 114 18 117 21 
rect 114 21 117 24 
rect 114 24 117 27 
rect 114 27 117 30 
rect 114 30 117 33 
rect 114 33 117 36 
rect 114 36 117 39 
rect 114 39 117 42 
rect 114 42 117 45 
rect 114 45 117 48 
rect 114 48 117 51 
rect 114 51 117 54 
rect 114 54 117 57 
rect 114 57 117 60 
rect 114 60 117 63 
rect 114 63 117 66 
rect 114 66 117 69 
rect 114 69 117 72 
rect 114 72 117 75 
rect 114 75 117 78 
rect 114 78 117 81 
rect 114 81 117 84 
rect 114 84 117 87 
rect 114 87 117 90 
rect 114 90 117 93 
rect 114 93 117 96 
rect 114 96 117 99 
rect 114 99 117 102 
rect 114 102 117 105 
rect 114 105 117 108 
rect 114 108 117 111 
rect 114 111 117 114 
rect 114 114 117 117 
rect 114 117 117 120 
rect 114 120 117 123 
rect 114 123 117 126 
rect 114 126 117 129 
rect 114 129 117 132 
rect 114 132 117 135 
rect 114 135 117 138 
rect 114 138 117 141 
rect 114 141 117 144 
rect 114 144 117 147 
rect 114 147 117 150 
rect 114 150 117 153 
rect 114 153 117 156 
rect 114 156 117 159 
rect 114 159 117 162 
rect 114 162 117 165 
rect 114 165 117 168 
rect 114 168 117 171 
rect 114 171 117 174 
rect 114 174 117 177 
rect 114 177 117 180 
rect 114 180 117 183 
rect 114 183 117 186 
rect 114 186 117 189 
rect 114 189 117 192 
rect 114 192 117 195 
rect 114 195 117 198 
rect 114 198 117 201 
rect 114 201 117 204 
rect 114 204 117 207 
rect 114 207 117 210 
rect 114 210 117 213 
rect 114 213 117 216 
rect 114 216 117 219 
rect 114 219 117 222 
rect 114 222 117 225 
rect 114 225 117 228 
rect 114 228 117 231 
rect 114 231 117 234 
rect 114 234 117 237 
rect 114 237 117 240 
rect 114 240 117 243 
rect 114 243 117 246 
rect 114 246 117 249 
rect 114 249 117 252 
rect 114 252 117 255 
rect 114 255 117 258 
rect 114 258 117 261 
rect 114 261 117 264 
rect 114 264 117 267 
rect 114 267 117 270 
rect 114 270 117 273 
rect 114 273 117 276 
rect 114 276 117 279 
rect 114 279 117 282 
rect 114 282 117 285 
rect 114 285 117 288 
rect 114 288 117 291 
rect 114 291 117 294 
rect 114 294 117 297 
rect 114 297 117 300 
rect 114 300 117 303 
rect 114 303 117 306 
rect 114 306 117 309 
rect 114 309 117 312 
rect 114 312 117 315 
rect 114 315 117 318 
rect 114 318 117 321 
rect 114 321 117 324 
rect 114 324 117 327 
rect 114 327 117 330 
rect 114 330 117 333 
rect 114 333 117 336 
rect 114 336 117 339 
rect 114 339 117 342 
rect 114 342 117 345 
rect 114 345 117 348 
rect 114 348 117 351 
rect 114 351 117 354 
rect 114 354 117 357 
rect 114 357 117 360 
rect 114 360 117 363 
rect 114 363 117 366 
rect 114 366 117 369 
rect 114 369 117 372 
rect 114 372 117 375 
rect 114 375 117 378 
rect 114 378 117 381 
rect 114 381 117 384 
rect 114 384 117 387 
rect 114 387 117 390 
rect 114 390 117 393 
rect 114 393 117 396 
rect 114 396 117 399 
rect 114 399 117 402 
rect 114 402 117 405 
rect 114 405 117 408 
rect 114 408 117 411 
rect 114 411 117 414 
rect 114 414 117 417 
rect 114 417 117 420 
rect 114 420 117 423 
rect 114 423 117 426 
rect 114 426 117 429 
rect 114 429 117 432 
rect 114 432 117 435 
rect 114 435 117 438 
rect 114 438 117 441 
rect 114 441 117 444 
rect 114 444 117 447 
rect 114 447 117 450 
rect 114 450 117 453 
rect 114 453 117 456 
rect 114 456 117 459 
rect 114 459 117 462 
rect 114 462 117 465 
rect 114 465 117 468 
rect 114 468 117 471 
rect 114 471 117 474 
rect 114 474 117 477 
rect 114 477 117 480 
rect 114 480 117 483 
rect 114 483 117 486 
rect 114 486 117 489 
rect 114 489 117 492 
rect 114 492 117 495 
rect 114 495 117 498 
rect 114 498 117 501 
rect 114 501 117 504 
rect 114 504 117 507 
rect 114 507 117 510 
rect 117 0 120 3 
rect 117 3 120 6 
rect 117 6 120 9 
rect 117 9 120 12 
rect 117 12 120 15 
rect 117 15 120 18 
rect 117 18 120 21 
rect 117 21 120 24 
rect 117 24 120 27 
rect 117 27 120 30 
rect 117 30 120 33 
rect 117 33 120 36 
rect 117 36 120 39 
rect 117 39 120 42 
rect 117 42 120 45 
rect 117 45 120 48 
rect 117 48 120 51 
rect 117 51 120 54 
rect 117 54 120 57 
rect 117 57 120 60 
rect 117 60 120 63 
rect 117 63 120 66 
rect 117 66 120 69 
rect 117 69 120 72 
rect 117 72 120 75 
rect 117 75 120 78 
rect 117 78 120 81 
rect 117 81 120 84 
rect 117 84 120 87 
rect 117 87 120 90 
rect 117 90 120 93 
rect 117 93 120 96 
rect 117 96 120 99 
rect 117 99 120 102 
rect 117 102 120 105 
rect 117 105 120 108 
rect 117 108 120 111 
rect 117 111 120 114 
rect 117 114 120 117 
rect 117 117 120 120 
rect 117 120 120 123 
rect 117 123 120 126 
rect 117 126 120 129 
rect 117 129 120 132 
rect 117 132 120 135 
rect 117 135 120 138 
rect 117 138 120 141 
rect 117 141 120 144 
rect 117 144 120 147 
rect 117 147 120 150 
rect 117 150 120 153 
rect 117 153 120 156 
rect 117 156 120 159 
rect 117 159 120 162 
rect 117 162 120 165 
rect 117 165 120 168 
rect 117 168 120 171 
rect 117 171 120 174 
rect 117 174 120 177 
rect 117 177 120 180 
rect 117 180 120 183 
rect 117 183 120 186 
rect 117 186 120 189 
rect 117 189 120 192 
rect 117 192 120 195 
rect 117 195 120 198 
rect 117 198 120 201 
rect 117 201 120 204 
rect 117 204 120 207 
rect 117 207 120 210 
rect 117 210 120 213 
rect 117 213 120 216 
rect 117 216 120 219 
rect 117 219 120 222 
rect 117 222 120 225 
rect 117 225 120 228 
rect 117 228 120 231 
rect 117 231 120 234 
rect 117 234 120 237 
rect 117 237 120 240 
rect 117 240 120 243 
rect 117 243 120 246 
rect 117 246 120 249 
rect 117 249 120 252 
rect 117 252 120 255 
rect 117 255 120 258 
rect 117 258 120 261 
rect 117 261 120 264 
rect 117 264 120 267 
rect 117 267 120 270 
rect 117 270 120 273 
rect 117 273 120 276 
rect 117 276 120 279 
rect 117 279 120 282 
rect 117 282 120 285 
rect 117 285 120 288 
rect 117 288 120 291 
rect 117 291 120 294 
rect 117 294 120 297 
rect 117 297 120 300 
rect 117 300 120 303 
rect 117 303 120 306 
rect 117 306 120 309 
rect 117 309 120 312 
rect 117 312 120 315 
rect 117 315 120 318 
rect 117 318 120 321 
rect 117 321 120 324 
rect 117 324 120 327 
rect 117 327 120 330 
rect 117 330 120 333 
rect 117 333 120 336 
rect 117 336 120 339 
rect 117 339 120 342 
rect 117 342 120 345 
rect 117 345 120 348 
rect 117 348 120 351 
rect 117 351 120 354 
rect 117 354 120 357 
rect 117 357 120 360 
rect 117 360 120 363 
rect 117 363 120 366 
rect 117 366 120 369 
rect 117 369 120 372 
rect 117 372 120 375 
rect 117 375 120 378 
rect 117 378 120 381 
rect 117 381 120 384 
rect 117 384 120 387 
rect 117 387 120 390 
rect 117 390 120 393 
rect 117 393 120 396 
rect 117 396 120 399 
rect 117 399 120 402 
rect 117 402 120 405 
rect 117 405 120 408 
rect 117 408 120 411 
rect 117 411 120 414 
rect 117 414 120 417 
rect 117 417 120 420 
rect 117 420 120 423 
rect 117 423 120 426 
rect 117 426 120 429 
rect 117 429 120 432 
rect 117 432 120 435 
rect 117 435 120 438 
rect 117 438 120 441 
rect 117 441 120 444 
rect 117 444 120 447 
rect 117 447 120 450 
rect 117 450 120 453 
rect 117 453 120 456 
rect 117 456 120 459 
rect 117 459 120 462 
rect 117 462 120 465 
rect 117 465 120 468 
rect 117 468 120 471 
rect 117 471 120 474 
rect 117 474 120 477 
rect 117 477 120 480 
rect 117 480 120 483 
rect 117 483 120 486 
rect 117 486 120 489 
rect 117 489 120 492 
rect 117 492 120 495 
rect 117 495 120 498 
rect 117 498 120 501 
rect 117 501 120 504 
rect 117 504 120 507 
rect 117 507 120 510 
rect 120 0 123 3 
rect 120 3 123 6 
rect 120 6 123 9 
rect 120 9 123 12 
rect 120 12 123 15 
rect 120 15 123 18 
rect 120 18 123 21 
rect 120 21 123 24 
rect 120 24 123 27 
rect 120 27 123 30 
rect 120 30 123 33 
rect 120 33 123 36 
rect 120 36 123 39 
rect 120 39 123 42 
rect 120 42 123 45 
rect 120 45 123 48 
rect 120 48 123 51 
rect 120 51 123 54 
rect 120 54 123 57 
rect 120 57 123 60 
rect 120 60 123 63 
rect 120 63 123 66 
rect 120 66 123 69 
rect 120 69 123 72 
rect 120 72 123 75 
rect 120 75 123 78 
rect 120 78 123 81 
rect 120 81 123 84 
rect 120 84 123 87 
rect 120 87 123 90 
rect 120 90 123 93 
rect 120 93 123 96 
rect 120 96 123 99 
rect 120 99 123 102 
rect 120 102 123 105 
rect 120 105 123 108 
rect 120 108 123 111 
rect 120 111 123 114 
rect 120 114 123 117 
rect 120 117 123 120 
rect 120 120 123 123 
rect 120 123 123 126 
rect 120 126 123 129 
rect 120 129 123 132 
rect 120 132 123 135 
rect 120 135 123 138 
rect 120 138 123 141 
rect 120 141 123 144 
rect 120 144 123 147 
rect 120 147 123 150 
rect 120 150 123 153 
rect 120 153 123 156 
rect 120 156 123 159 
rect 120 159 123 162 
rect 120 162 123 165 
rect 120 165 123 168 
rect 120 168 123 171 
rect 120 171 123 174 
rect 120 174 123 177 
rect 120 177 123 180 
rect 120 180 123 183 
rect 120 183 123 186 
rect 120 186 123 189 
rect 120 189 123 192 
rect 120 192 123 195 
rect 120 195 123 198 
rect 120 198 123 201 
rect 120 201 123 204 
rect 120 204 123 207 
rect 120 207 123 210 
rect 120 210 123 213 
rect 120 213 123 216 
rect 120 216 123 219 
rect 120 219 123 222 
rect 120 222 123 225 
rect 120 225 123 228 
rect 120 228 123 231 
rect 120 231 123 234 
rect 120 234 123 237 
rect 120 237 123 240 
rect 120 240 123 243 
rect 120 243 123 246 
rect 120 246 123 249 
rect 120 249 123 252 
rect 120 252 123 255 
rect 120 255 123 258 
rect 120 258 123 261 
rect 120 261 123 264 
rect 120 264 123 267 
rect 120 267 123 270 
rect 120 270 123 273 
rect 120 273 123 276 
rect 120 276 123 279 
rect 120 279 123 282 
rect 120 282 123 285 
rect 120 285 123 288 
rect 120 288 123 291 
rect 120 291 123 294 
rect 120 294 123 297 
rect 120 297 123 300 
rect 120 300 123 303 
rect 120 303 123 306 
rect 120 306 123 309 
rect 120 309 123 312 
rect 120 312 123 315 
rect 120 315 123 318 
rect 120 318 123 321 
rect 120 321 123 324 
rect 120 324 123 327 
rect 120 327 123 330 
rect 120 330 123 333 
rect 120 333 123 336 
rect 120 336 123 339 
rect 120 339 123 342 
rect 120 342 123 345 
rect 120 345 123 348 
rect 120 348 123 351 
rect 120 351 123 354 
rect 120 354 123 357 
rect 120 357 123 360 
rect 120 360 123 363 
rect 120 363 123 366 
rect 120 366 123 369 
rect 120 369 123 372 
rect 120 372 123 375 
rect 120 375 123 378 
rect 120 378 123 381 
rect 120 381 123 384 
rect 120 384 123 387 
rect 120 387 123 390 
rect 120 390 123 393 
rect 120 393 123 396 
rect 120 396 123 399 
rect 120 399 123 402 
rect 120 402 123 405 
rect 120 405 123 408 
rect 120 408 123 411 
rect 120 411 123 414 
rect 120 414 123 417 
rect 120 417 123 420 
rect 120 420 123 423 
rect 120 423 123 426 
rect 120 426 123 429 
rect 120 429 123 432 
rect 120 432 123 435 
rect 120 435 123 438 
rect 120 438 123 441 
rect 120 441 123 444 
rect 120 444 123 447 
rect 120 447 123 450 
rect 120 450 123 453 
rect 120 453 123 456 
rect 120 456 123 459 
rect 120 459 123 462 
rect 120 462 123 465 
rect 120 465 123 468 
rect 120 468 123 471 
rect 120 471 123 474 
rect 120 474 123 477 
rect 120 477 123 480 
rect 120 480 123 483 
rect 120 483 123 486 
rect 120 486 123 489 
rect 120 489 123 492 
rect 120 492 123 495 
rect 120 495 123 498 
rect 120 498 123 501 
rect 120 501 123 504 
rect 120 504 123 507 
rect 120 507 123 510 
rect 123 0 126 3 
rect 123 3 126 6 
rect 123 6 126 9 
rect 123 9 126 12 
rect 123 12 126 15 
rect 123 15 126 18 
rect 123 18 126 21 
rect 123 21 126 24 
rect 123 24 126 27 
rect 123 27 126 30 
rect 123 30 126 33 
rect 123 33 126 36 
rect 123 36 126 39 
rect 123 39 126 42 
rect 123 42 126 45 
rect 123 45 126 48 
rect 123 48 126 51 
rect 123 51 126 54 
rect 123 54 126 57 
rect 123 57 126 60 
rect 123 60 126 63 
rect 123 63 126 66 
rect 123 66 126 69 
rect 123 69 126 72 
rect 123 72 126 75 
rect 123 75 126 78 
rect 123 78 126 81 
rect 123 81 126 84 
rect 123 84 126 87 
rect 123 87 126 90 
rect 123 90 126 93 
rect 123 93 126 96 
rect 123 96 126 99 
rect 123 99 126 102 
rect 123 102 126 105 
rect 123 105 126 108 
rect 123 108 126 111 
rect 123 111 126 114 
rect 123 114 126 117 
rect 123 117 126 120 
rect 123 120 126 123 
rect 123 123 126 126 
rect 123 126 126 129 
rect 123 129 126 132 
rect 123 132 126 135 
rect 123 135 126 138 
rect 123 138 126 141 
rect 123 141 126 144 
rect 123 144 126 147 
rect 123 147 126 150 
rect 123 150 126 153 
rect 123 153 126 156 
rect 123 156 126 159 
rect 123 159 126 162 
rect 123 162 126 165 
rect 123 165 126 168 
rect 123 168 126 171 
rect 123 171 126 174 
rect 123 174 126 177 
rect 123 177 126 180 
rect 123 180 126 183 
rect 123 183 126 186 
rect 123 186 126 189 
rect 123 189 126 192 
rect 123 192 126 195 
rect 123 195 126 198 
rect 123 198 126 201 
rect 123 201 126 204 
rect 123 204 126 207 
rect 123 207 126 210 
rect 123 210 126 213 
rect 123 213 126 216 
rect 123 216 126 219 
rect 123 219 126 222 
rect 123 222 126 225 
rect 123 225 126 228 
rect 123 228 126 231 
rect 123 231 126 234 
rect 123 234 126 237 
rect 123 237 126 240 
rect 123 240 126 243 
rect 123 243 126 246 
rect 123 246 126 249 
rect 123 249 126 252 
rect 123 252 126 255 
rect 123 255 126 258 
rect 123 258 126 261 
rect 123 261 126 264 
rect 123 264 126 267 
rect 123 267 126 270 
rect 123 270 126 273 
rect 123 273 126 276 
rect 123 276 126 279 
rect 123 279 126 282 
rect 123 282 126 285 
rect 123 285 126 288 
rect 123 288 126 291 
rect 123 291 126 294 
rect 123 294 126 297 
rect 123 297 126 300 
rect 123 300 126 303 
rect 123 303 126 306 
rect 123 306 126 309 
rect 123 309 126 312 
rect 123 312 126 315 
rect 123 315 126 318 
rect 123 318 126 321 
rect 123 321 126 324 
rect 123 324 126 327 
rect 123 327 126 330 
rect 123 330 126 333 
rect 123 333 126 336 
rect 123 336 126 339 
rect 123 339 126 342 
rect 123 342 126 345 
rect 123 345 126 348 
rect 123 348 126 351 
rect 123 351 126 354 
rect 123 354 126 357 
rect 123 357 126 360 
rect 123 360 126 363 
rect 123 363 126 366 
rect 123 366 126 369 
rect 123 369 126 372 
rect 123 372 126 375 
rect 123 375 126 378 
rect 123 378 126 381 
rect 123 381 126 384 
rect 123 384 126 387 
rect 123 387 126 390 
rect 123 390 126 393 
rect 123 393 126 396 
rect 123 396 126 399 
rect 123 399 126 402 
rect 123 402 126 405 
rect 123 405 126 408 
rect 123 408 126 411 
rect 123 411 126 414 
rect 123 414 126 417 
rect 123 417 126 420 
rect 123 420 126 423 
rect 123 423 126 426 
rect 123 426 126 429 
rect 123 429 126 432 
rect 123 432 126 435 
rect 123 435 126 438 
rect 123 438 126 441 
rect 123 441 126 444 
rect 123 444 126 447 
rect 123 447 126 450 
rect 123 450 126 453 
rect 123 453 126 456 
rect 123 456 126 459 
rect 123 459 126 462 
rect 123 462 126 465 
rect 123 465 126 468 
rect 123 468 126 471 
rect 123 471 126 474 
rect 123 474 126 477 
rect 123 477 126 480 
rect 123 480 126 483 
rect 123 483 126 486 
rect 123 486 126 489 
rect 123 489 126 492 
rect 123 492 126 495 
rect 123 495 126 498 
rect 123 498 126 501 
rect 123 501 126 504 
rect 123 504 126 507 
rect 123 507 126 510 
rect 126 0 129 3 
rect 126 3 129 6 
rect 126 6 129 9 
rect 126 9 129 12 
rect 126 12 129 15 
rect 126 15 129 18 
rect 126 18 129 21 
rect 126 21 129 24 
rect 126 24 129 27 
rect 126 27 129 30 
rect 126 30 129 33 
rect 126 33 129 36 
rect 126 36 129 39 
rect 126 39 129 42 
rect 126 42 129 45 
rect 126 45 129 48 
rect 126 48 129 51 
rect 126 51 129 54 
rect 126 54 129 57 
rect 126 57 129 60 
rect 126 60 129 63 
rect 126 63 129 66 
rect 126 66 129 69 
rect 126 69 129 72 
rect 126 72 129 75 
rect 126 75 129 78 
rect 126 78 129 81 
rect 126 81 129 84 
rect 126 84 129 87 
rect 126 87 129 90 
rect 126 90 129 93 
rect 126 93 129 96 
rect 126 96 129 99 
rect 126 99 129 102 
rect 126 102 129 105 
rect 126 105 129 108 
rect 126 108 129 111 
rect 126 111 129 114 
rect 126 114 129 117 
rect 126 117 129 120 
rect 126 120 129 123 
rect 126 123 129 126 
rect 126 126 129 129 
rect 126 129 129 132 
rect 126 132 129 135 
rect 126 135 129 138 
rect 126 138 129 141 
rect 126 141 129 144 
rect 126 144 129 147 
rect 126 147 129 150 
rect 126 150 129 153 
rect 126 153 129 156 
rect 126 156 129 159 
rect 126 159 129 162 
rect 126 162 129 165 
rect 126 165 129 168 
rect 126 168 129 171 
rect 126 171 129 174 
rect 126 174 129 177 
rect 126 177 129 180 
rect 126 180 129 183 
rect 126 183 129 186 
rect 126 186 129 189 
rect 126 189 129 192 
rect 126 192 129 195 
rect 126 195 129 198 
rect 126 198 129 201 
rect 126 201 129 204 
rect 126 204 129 207 
rect 126 207 129 210 
rect 126 210 129 213 
rect 126 213 129 216 
rect 126 216 129 219 
rect 126 219 129 222 
rect 126 222 129 225 
rect 126 225 129 228 
rect 126 228 129 231 
rect 126 231 129 234 
rect 126 234 129 237 
rect 126 237 129 240 
rect 126 240 129 243 
rect 126 243 129 246 
rect 126 246 129 249 
rect 126 249 129 252 
rect 126 252 129 255 
rect 126 255 129 258 
rect 126 258 129 261 
rect 126 261 129 264 
rect 126 264 129 267 
rect 126 267 129 270 
rect 126 270 129 273 
rect 126 273 129 276 
rect 126 276 129 279 
rect 126 279 129 282 
rect 126 282 129 285 
rect 126 285 129 288 
rect 126 288 129 291 
rect 126 291 129 294 
rect 126 294 129 297 
rect 126 297 129 300 
rect 126 300 129 303 
rect 126 303 129 306 
rect 126 306 129 309 
rect 126 309 129 312 
rect 126 312 129 315 
rect 126 315 129 318 
rect 126 318 129 321 
rect 126 321 129 324 
rect 126 324 129 327 
rect 126 327 129 330 
rect 126 330 129 333 
rect 126 333 129 336 
rect 126 336 129 339 
rect 126 339 129 342 
rect 126 342 129 345 
rect 126 345 129 348 
rect 126 348 129 351 
rect 126 351 129 354 
rect 126 354 129 357 
rect 126 357 129 360 
rect 126 360 129 363 
rect 126 363 129 366 
rect 126 366 129 369 
rect 126 369 129 372 
rect 126 372 129 375 
rect 126 375 129 378 
rect 126 378 129 381 
rect 126 381 129 384 
rect 126 384 129 387 
rect 126 387 129 390 
rect 126 390 129 393 
rect 126 393 129 396 
rect 126 396 129 399 
rect 126 399 129 402 
rect 126 402 129 405 
rect 126 405 129 408 
rect 126 408 129 411 
rect 126 411 129 414 
rect 126 414 129 417 
rect 126 417 129 420 
rect 126 420 129 423 
rect 126 423 129 426 
rect 126 426 129 429 
rect 126 429 129 432 
rect 126 432 129 435 
rect 126 435 129 438 
rect 126 438 129 441 
rect 126 441 129 444 
rect 126 444 129 447 
rect 126 447 129 450 
rect 126 450 129 453 
rect 126 453 129 456 
rect 126 456 129 459 
rect 126 459 129 462 
rect 126 462 129 465 
rect 126 465 129 468 
rect 126 468 129 471 
rect 126 471 129 474 
rect 126 474 129 477 
rect 126 477 129 480 
rect 126 480 129 483 
rect 126 483 129 486 
rect 126 486 129 489 
rect 126 489 129 492 
rect 126 492 129 495 
rect 126 495 129 498 
rect 126 498 129 501 
rect 126 501 129 504 
rect 126 504 129 507 
rect 126 507 129 510 
rect 129 0 132 3 
rect 129 3 132 6 
rect 129 6 132 9 
rect 129 9 132 12 
rect 129 12 132 15 
rect 129 15 132 18 
rect 129 18 132 21 
rect 129 21 132 24 
rect 129 24 132 27 
rect 129 27 132 30 
rect 129 30 132 33 
rect 129 33 132 36 
rect 129 36 132 39 
rect 129 39 132 42 
rect 129 42 132 45 
rect 129 45 132 48 
rect 129 48 132 51 
rect 129 51 132 54 
rect 129 54 132 57 
rect 129 57 132 60 
rect 129 60 132 63 
rect 129 63 132 66 
rect 129 66 132 69 
rect 129 69 132 72 
rect 129 72 132 75 
rect 129 75 132 78 
rect 129 78 132 81 
rect 129 81 132 84 
rect 129 84 132 87 
rect 129 87 132 90 
rect 129 90 132 93 
rect 129 93 132 96 
rect 129 96 132 99 
rect 129 99 132 102 
rect 129 102 132 105 
rect 129 105 132 108 
rect 129 108 132 111 
rect 129 111 132 114 
rect 129 114 132 117 
rect 129 117 132 120 
rect 129 120 132 123 
rect 129 123 132 126 
rect 129 126 132 129 
rect 129 129 132 132 
rect 129 132 132 135 
rect 129 135 132 138 
rect 129 138 132 141 
rect 129 141 132 144 
rect 129 144 132 147 
rect 129 147 132 150 
rect 129 150 132 153 
rect 129 153 132 156 
rect 129 156 132 159 
rect 129 159 132 162 
rect 129 162 132 165 
rect 129 165 132 168 
rect 129 168 132 171 
rect 129 171 132 174 
rect 129 174 132 177 
rect 129 177 132 180 
rect 129 180 132 183 
rect 129 183 132 186 
rect 129 186 132 189 
rect 129 189 132 192 
rect 129 192 132 195 
rect 129 195 132 198 
rect 129 198 132 201 
rect 129 201 132 204 
rect 129 204 132 207 
rect 129 207 132 210 
rect 129 210 132 213 
rect 129 213 132 216 
rect 129 216 132 219 
rect 129 219 132 222 
rect 129 222 132 225 
rect 129 225 132 228 
rect 129 228 132 231 
rect 129 231 132 234 
rect 129 234 132 237 
rect 129 237 132 240 
rect 129 240 132 243 
rect 129 243 132 246 
rect 129 246 132 249 
rect 129 249 132 252 
rect 129 252 132 255 
rect 129 255 132 258 
rect 129 258 132 261 
rect 129 261 132 264 
rect 129 264 132 267 
rect 129 267 132 270 
rect 129 270 132 273 
rect 129 273 132 276 
rect 129 276 132 279 
rect 129 279 132 282 
rect 129 282 132 285 
rect 129 285 132 288 
rect 129 288 132 291 
rect 129 291 132 294 
rect 129 294 132 297 
rect 129 297 132 300 
rect 129 300 132 303 
rect 129 303 132 306 
rect 129 306 132 309 
rect 129 309 132 312 
rect 129 312 132 315 
rect 129 315 132 318 
rect 129 318 132 321 
rect 129 321 132 324 
rect 129 324 132 327 
rect 129 327 132 330 
rect 129 330 132 333 
rect 129 333 132 336 
rect 129 336 132 339 
rect 129 339 132 342 
rect 129 342 132 345 
rect 129 345 132 348 
rect 129 348 132 351 
rect 129 351 132 354 
rect 129 354 132 357 
rect 129 357 132 360 
rect 129 360 132 363 
rect 129 363 132 366 
rect 129 366 132 369 
rect 129 369 132 372 
rect 129 372 132 375 
rect 129 375 132 378 
rect 129 378 132 381 
rect 129 381 132 384 
rect 129 384 132 387 
rect 129 387 132 390 
rect 129 390 132 393 
rect 129 393 132 396 
rect 129 396 132 399 
rect 129 399 132 402 
rect 129 402 132 405 
rect 129 405 132 408 
rect 129 408 132 411 
rect 129 411 132 414 
rect 129 414 132 417 
rect 129 417 132 420 
rect 129 420 132 423 
rect 129 423 132 426 
rect 129 426 132 429 
rect 129 429 132 432 
rect 129 432 132 435 
rect 129 435 132 438 
rect 129 438 132 441 
rect 129 441 132 444 
rect 129 444 132 447 
rect 129 447 132 450 
rect 129 450 132 453 
rect 129 453 132 456 
rect 129 456 132 459 
rect 129 459 132 462 
rect 129 462 132 465 
rect 129 465 132 468 
rect 129 468 132 471 
rect 129 471 132 474 
rect 129 474 132 477 
rect 129 477 132 480 
rect 129 480 132 483 
rect 129 483 132 486 
rect 129 486 132 489 
rect 129 489 132 492 
rect 129 492 132 495 
rect 129 495 132 498 
rect 129 498 132 501 
rect 129 501 132 504 
rect 129 504 132 507 
rect 129 507 132 510 
rect 132 0 135 3 
rect 132 3 135 6 
rect 132 6 135 9 
rect 132 9 135 12 
rect 132 12 135 15 
rect 132 15 135 18 
rect 132 18 135 21 
rect 132 21 135 24 
rect 132 24 135 27 
rect 132 27 135 30 
rect 132 30 135 33 
rect 132 33 135 36 
rect 132 36 135 39 
rect 132 39 135 42 
rect 132 42 135 45 
rect 132 45 135 48 
rect 132 48 135 51 
rect 132 51 135 54 
rect 132 54 135 57 
rect 132 57 135 60 
rect 132 60 135 63 
rect 132 63 135 66 
rect 132 66 135 69 
rect 132 69 135 72 
rect 132 72 135 75 
rect 132 75 135 78 
rect 132 78 135 81 
rect 132 81 135 84 
rect 132 84 135 87 
rect 132 87 135 90 
rect 132 90 135 93 
rect 132 93 135 96 
rect 132 96 135 99 
rect 132 99 135 102 
rect 132 102 135 105 
rect 132 105 135 108 
rect 132 108 135 111 
rect 132 111 135 114 
rect 132 114 135 117 
rect 132 117 135 120 
rect 132 120 135 123 
rect 132 123 135 126 
rect 132 126 135 129 
rect 132 129 135 132 
rect 132 132 135 135 
rect 132 135 135 138 
rect 132 138 135 141 
rect 132 141 135 144 
rect 132 144 135 147 
rect 132 147 135 150 
rect 132 150 135 153 
rect 132 153 135 156 
rect 132 156 135 159 
rect 132 159 135 162 
rect 132 162 135 165 
rect 132 165 135 168 
rect 132 168 135 171 
rect 132 171 135 174 
rect 132 174 135 177 
rect 132 177 135 180 
rect 132 180 135 183 
rect 132 183 135 186 
rect 132 186 135 189 
rect 132 189 135 192 
rect 132 192 135 195 
rect 132 195 135 198 
rect 132 198 135 201 
rect 132 201 135 204 
rect 132 204 135 207 
rect 132 207 135 210 
rect 132 210 135 213 
rect 132 213 135 216 
rect 132 216 135 219 
rect 132 219 135 222 
rect 132 222 135 225 
rect 132 225 135 228 
rect 132 228 135 231 
rect 132 231 135 234 
rect 132 234 135 237 
rect 132 237 135 240 
rect 132 240 135 243 
rect 132 243 135 246 
rect 132 246 135 249 
rect 132 249 135 252 
rect 132 252 135 255 
rect 132 255 135 258 
rect 132 258 135 261 
rect 132 261 135 264 
rect 132 264 135 267 
rect 132 267 135 270 
rect 132 270 135 273 
rect 132 273 135 276 
rect 132 276 135 279 
rect 132 279 135 282 
rect 132 282 135 285 
rect 132 285 135 288 
rect 132 288 135 291 
rect 132 291 135 294 
rect 132 294 135 297 
rect 132 297 135 300 
rect 132 300 135 303 
rect 132 303 135 306 
rect 132 306 135 309 
rect 132 309 135 312 
rect 132 312 135 315 
rect 132 315 135 318 
rect 132 318 135 321 
rect 132 321 135 324 
rect 132 324 135 327 
rect 132 327 135 330 
rect 132 330 135 333 
rect 132 333 135 336 
rect 132 336 135 339 
rect 132 339 135 342 
rect 132 342 135 345 
rect 132 345 135 348 
rect 132 348 135 351 
rect 132 351 135 354 
rect 132 354 135 357 
rect 132 357 135 360 
rect 132 360 135 363 
rect 132 363 135 366 
rect 132 366 135 369 
rect 132 369 135 372 
rect 132 372 135 375 
rect 132 375 135 378 
rect 132 378 135 381 
rect 132 381 135 384 
rect 132 384 135 387 
rect 132 387 135 390 
rect 132 390 135 393 
rect 132 393 135 396 
rect 132 396 135 399 
rect 132 399 135 402 
rect 132 402 135 405 
rect 132 405 135 408 
rect 132 408 135 411 
rect 132 411 135 414 
rect 132 414 135 417 
rect 132 417 135 420 
rect 132 420 135 423 
rect 132 423 135 426 
rect 132 426 135 429 
rect 132 429 135 432 
rect 132 432 135 435 
rect 132 435 135 438 
rect 132 438 135 441 
rect 132 441 135 444 
rect 132 444 135 447 
rect 132 447 135 450 
rect 132 450 135 453 
rect 132 453 135 456 
rect 132 456 135 459 
rect 132 459 135 462 
rect 132 462 135 465 
rect 132 465 135 468 
rect 132 468 135 471 
rect 132 471 135 474 
rect 132 474 135 477 
rect 132 477 135 480 
rect 132 480 135 483 
rect 132 483 135 486 
rect 132 486 135 489 
rect 132 489 135 492 
rect 132 492 135 495 
rect 132 495 135 498 
rect 132 498 135 501 
rect 132 501 135 504 
rect 132 504 135 507 
rect 132 507 135 510 
rect 135 0 138 3 
rect 135 3 138 6 
rect 135 6 138 9 
rect 135 9 138 12 
rect 135 12 138 15 
rect 135 15 138 18 
rect 135 18 138 21 
rect 135 21 138 24 
rect 135 24 138 27 
rect 135 27 138 30 
rect 135 30 138 33 
rect 135 33 138 36 
rect 135 36 138 39 
rect 135 39 138 42 
rect 135 42 138 45 
rect 135 45 138 48 
rect 135 48 138 51 
rect 135 51 138 54 
rect 135 54 138 57 
rect 135 57 138 60 
rect 135 60 138 63 
rect 135 63 138 66 
rect 135 66 138 69 
rect 135 69 138 72 
rect 135 72 138 75 
rect 135 75 138 78 
rect 135 78 138 81 
rect 135 81 138 84 
rect 135 84 138 87 
rect 135 87 138 90 
rect 135 90 138 93 
rect 135 93 138 96 
rect 135 96 138 99 
rect 135 99 138 102 
rect 135 102 138 105 
rect 135 105 138 108 
rect 135 108 138 111 
rect 135 111 138 114 
rect 135 114 138 117 
rect 135 117 138 120 
rect 135 120 138 123 
rect 135 123 138 126 
rect 135 126 138 129 
rect 135 129 138 132 
rect 135 132 138 135 
rect 135 135 138 138 
rect 135 138 138 141 
rect 135 141 138 144 
rect 135 144 138 147 
rect 135 147 138 150 
rect 135 150 138 153 
rect 135 153 138 156 
rect 135 156 138 159 
rect 135 159 138 162 
rect 135 162 138 165 
rect 135 165 138 168 
rect 135 168 138 171 
rect 135 171 138 174 
rect 135 174 138 177 
rect 135 177 138 180 
rect 135 180 138 183 
rect 135 183 138 186 
rect 135 186 138 189 
rect 135 189 138 192 
rect 135 192 138 195 
rect 135 195 138 198 
rect 135 198 138 201 
rect 135 201 138 204 
rect 135 204 138 207 
rect 135 207 138 210 
rect 135 210 138 213 
rect 135 213 138 216 
rect 135 216 138 219 
rect 135 219 138 222 
rect 135 222 138 225 
rect 135 225 138 228 
rect 135 228 138 231 
rect 135 231 138 234 
rect 135 234 138 237 
rect 135 237 138 240 
rect 135 240 138 243 
rect 135 243 138 246 
rect 135 246 138 249 
rect 135 249 138 252 
rect 135 252 138 255 
rect 135 255 138 258 
rect 135 258 138 261 
rect 135 261 138 264 
rect 135 264 138 267 
rect 135 267 138 270 
rect 135 270 138 273 
rect 135 273 138 276 
rect 135 276 138 279 
rect 135 279 138 282 
rect 135 282 138 285 
rect 135 285 138 288 
rect 135 288 138 291 
rect 135 291 138 294 
rect 135 294 138 297 
rect 135 297 138 300 
rect 135 300 138 303 
rect 135 303 138 306 
rect 135 306 138 309 
rect 135 309 138 312 
rect 135 312 138 315 
rect 135 315 138 318 
rect 135 318 138 321 
rect 135 321 138 324 
rect 135 324 138 327 
rect 135 327 138 330 
rect 135 330 138 333 
rect 135 333 138 336 
rect 135 336 138 339 
rect 135 339 138 342 
rect 135 342 138 345 
rect 135 345 138 348 
rect 135 348 138 351 
rect 135 351 138 354 
rect 135 354 138 357 
rect 135 357 138 360 
rect 135 360 138 363 
rect 135 363 138 366 
rect 135 366 138 369 
rect 135 369 138 372 
rect 135 372 138 375 
rect 135 375 138 378 
rect 135 378 138 381 
rect 135 381 138 384 
rect 135 384 138 387 
rect 135 387 138 390 
rect 135 390 138 393 
rect 135 393 138 396 
rect 135 396 138 399 
rect 135 399 138 402 
rect 135 402 138 405 
rect 135 405 138 408 
rect 135 408 138 411 
rect 135 411 138 414 
rect 135 414 138 417 
rect 135 417 138 420 
rect 135 420 138 423 
rect 135 423 138 426 
rect 135 426 138 429 
rect 135 429 138 432 
rect 135 432 138 435 
rect 135 435 138 438 
rect 135 438 138 441 
rect 135 441 138 444 
rect 135 444 138 447 
rect 135 447 138 450 
rect 135 450 138 453 
rect 135 453 138 456 
rect 135 456 138 459 
rect 135 459 138 462 
rect 135 462 138 465 
rect 135 465 138 468 
rect 135 468 138 471 
rect 135 471 138 474 
rect 135 474 138 477 
rect 135 477 138 480 
rect 135 480 138 483 
rect 135 483 138 486 
rect 135 486 138 489 
rect 135 489 138 492 
rect 135 492 138 495 
rect 135 495 138 498 
rect 135 498 138 501 
rect 135 501 138 504 
rect 135 504 138 507 
rect 135 507 138 510 
rect 138 0 141 3 
rect 138 3 141 6 
rect 138 6 141 9 
rect 138 9 141 12 
rect 138 12 141 15 
rect 138 15 141 18 
rect 138 18 141 21 
rect 138 21 141 24 
rect 138 24 141 27 
rect 138 27 141 30 
rect 138 30 141 33 
rect 138 33 141 36 
rect 138 36 141 39 
rect 138 39 141 42 
rect 138 42 141 45 
rect 138 45 141 48 
rect 138 48 141 51 
rect 138 51 141 54 
rect 138 54 141 57 
rect 138 57 141 60 
rect 138 60 141 63 
rect 138 63 141 66 
rect 138 66 141 69 
rect 138 69 141 72 
rect 138 72 141 75 
rect 138 75 141 78 
rect 138 78 141 81 
rect 138 81 141 84 
rect 138 84 141 87 
rect 138 87 141 90 
rect 138 90 141 93 
rect 138 93 141 96 
rect 138 96 141 99 
rect 138 99 141 102 
rect 138 102 141 105 
rect 138 105 141 108 
rect 138 108 141 111 
rect 138 111 141 114 
rect 138 114 141 117 
rect 138 117 141 120 
rect 138 120 141 123 
rect 138 123 141 126 
rect 138 126 141 129 
rect 138 129 141 132 
rect 138 132 141 135 
rect 138 135 141 138 
rect 138 138 141 141 
rect 138 141 141 144 
rect 138 144 141 147 
rect 138 147 141 150 
rect 138 150 141 153 
rect 138 153 141 156 
rect 138 156 141 159 
rect 138 159 141 162 
rect 138 162 141 165 
rect 138 165 141 168 
rect 138 168 141 171 
rect 138 171 141 174 
rect 138 174 141 177 
rect 138 177 141 180 
rect 138 180 141 183 
rect 138 183 141 186 
rect 138 186 141 189 
rect 138 189 141 192 
rect 138 192 141 195 
rect 138 195 141 198 
rect 138 198 141 201 
rect 138 201 141 204 
rect 138 204 141 207 
rect 138 207 141 210 
rect 138 210 141 213 
rect 138 213 141 216 
rect 138 216 141 219 
rect 138 219 141 222 
rect 138 222 141 225 
rect 138 225 141 228 
rect 138 228 141 231 
rect 138 231 141 234 
rect 138 234 141 237 
rect 138 237 141 240 
rect 138 240 141 243 
rect 138 243 141 246 
rect 138 246 141 249 
rect 138 249 141 252 
rect 138 252 141 255 
rect 138 255 141 258 
rect 138 258 141 261 
rect 138 261 141 264 
rect 138 264 141 267 
rect 138 267 141 270 
rect 138 270 141 273 
rect 138 273 141 276 
rect 138 276 141 279 
rect 138 279 141 282 
rect 138 282 141 285 
rect 138 285 141 288 
rect 138 288 141 291 
rect 138 291 141 294 
rect 138 294 141 297 
rect 138 297 141 300 
rect 138 300 141 303 
rect 138 303 141 306 
rect 138 306 141 309 
rect 138 309 141 312 
rect 138 312 141 315 
rect 138 315 141 318 
rect 138 318 141 321 
rect 138 321 141 324 
rect 138 324 141 327 
rect 138 327 141 330 
rect 138 330 141 333 
rect 138 333 141 336 
rect 138 336 141 339 
rect 138 339 141 342 
rect 138 342 141 345 
rect 138 345 141 348 
rect 138 348 141 351 
rect 138 351 141 354 
rect 138 354 141 357 
rect 138 357 141 360 
rect 138 360 141 363 
rect 138 363 141 366 
rect 138 366 141 369 
rect 138 369 141 372 
rect 138 372 141 375 
rect 138 375 141 378 
rect 138 378 141 381 
rect 138 381 141 384 
rect 138 384 141 387 
rect 138 387 141 390 
rect 138 390 141 393 
rect 138 393 141 396 
rect 138 396 141 399 
rect 138 399 141 402 
rect 138 402 141 405 
rect 138 405 141 408 
rect 138 408 141 411 
rect 138 411 141 414 
rect 138 414 141 417 
rect 138 417 141 420 
rect 138 420 141 423 
rect 138 423 141 426 
rect 138 426 141 429 
rect 138 429 141 432 
rect 138 432 141 435 
rect 138 435 141 438 
rect 138 438 141 441 
rect 138 441 141 444 
rect 138 444 141 447 
rect 138 447 141 450 
rect 138 450 141 453 
rect 138 453 141 456 
rect 138 456 141 459 
rect 138 459 141 462 
rect 138 462 141 465 
rect 138 465 141 468 
rect 138 468 141 471 
rect 138 471 141 474 
rect 138 474 141 477 
rect 138 477 141 480 
rect 138 480 141 483 
rect 138 483 141 486 
rect 138 486 141 489 
rect 138 489 141 492 
rect 138 492 141 495 
rect 138 495 141 498 
rect 138 498 141 501 
rect 138 501 141 504 
rect 138 504 141 507 
rect 138 507 141 510 
rect 141 0 144 3 
rect 141 3 144 6 
rect 141 6 144 9 
rect 141 9 144 12 
rect 141 12 144 15 
rect 141 15 144 18 
rect 141 18 144 21 
rect 141 21 144 24 
rect 141 24 144 27 
rect 141 27 144 30 
rect 141 30 144 33 
rect 141 33 144 36 
rect 141 36 144 39 
rect 141 39 144 42 
rect 141 42 144 45 
rect 141 45 144 48 
rect 141 48 144 51 
rect 141 51 144 54 
rect 141 54 144 57 
rect 141 57 144 60 
rect 141 60 144 63 
rect 141 63 144 66 
rect 141 66 144 69 
rect 141 69 144 72 
rect 141 72 144 75 
rect 141 75 144 78 
rect 141 78 144 81 
rect 141 81 144 84 
rect 141 84 144 87 
rect 141 87 144 90 
rect 141 90 144 93 
rect 141 93 144 96 
rect 141 96 144 99 
rect 141 99 144 102 
rect 141 102 144 105 
rect 141 105 144 108 
rect 141 108 144 111 
rect 141 111 144 114 
rect 141 114 144 117 
rect 141 117 144 120 
rect 141 120 144 123 
rect 141 123 144 126 
rect 141 126 144 129 
rect 141 129 144 132 
rect 141 132 144 135 
rect 141 135 144 138 
rect 141 138 144 141 
rect 141 141 144 144 
rect 141 144 144 147 
rect 141 147 144 150 
rect 141 150 144 153 
rect 141 153 144 156 
rect 141 156 144 159 
rect 141 159 144 162 
rect 141 162 144 165 
rect 141 165 144 168 
rect 141 168 144 171 
rect 141 171 144 174 
rect 141 174 144 177 
rect 141 177 144 180 
rect 141 180 144 183 
rect 141 183 144 186 
rect 141 186 144 189 
rect 141 189 144 192 
rect 141 192 144 195 
rect 141 195 144 198 
rect 141 198 144 201 
rect 141 201 144 204 
rect 141 204 144 207 
rect 141 207 144 210 
rect 141 210 144 213 
rect 141 213 144 216 
rect 141 216 144 219 
rect 141 219 144 222 
rect 141 222 144 225 
rect 141 225 144 228 
rect 141 228 144 231 
rect 141 231 144 234 
rect 141 234 144 237 
rect 141 237 144 240 
rect 141 240 144 243 
rect 141 243 144 246 
rect 141 246 144 249 
rect 141 249 144 252 
rect 141 252 144 255 
rect 141 255 144 258 
rect 141 258 144 261 
rect 141 261 144 264 
rect 141 264 144 267 
rect 141 267 144 270 
rect 141 270 144 273 
rect 141 273 144 276 
rect 141 276 144 279 
rect 141 279 144 282 
rect 141 282 144 285 
rect 141 285 144 288 
rect 141 288 144 291 
rect 141 291 144 294 
rect 141 294 144 297 
rect 141 297 144 300 
rect 141 300 144 303 
rect 141 303 144 306 
rect 141 306 144 309 
rect 141 309 144 312 
rect 141 312 144 315 
rect 141 315 144 318 
rect 141 318 144 321 
rect 141 321 144 324 
rect 141 324 144 327 
rect 141 327 144 330 
rect 141 330 144 333 
rect 141 333 144 336 
rect 141 336 144 339 
rect 141 339 144 342 
rect 141 342 144 345 
rect 141 345 144 348 
rect 141 348 144 351 
rect 141 351 144 354 
rect 141 354 144 357 
rect 141 357 144 360 
rect 141 360 144 363 
rect 141 363 144 366 
rect 141 366 144 369 
rect 141 369 144 372 
rect 141 372 144 375 
rect 141 375 144 378 
rect 141 378 144 381 
rect 141 381 144 384 
rect 141 384 144 387 
rect 141 387 144 390 
rect 141 390 144 393 
rect 141 393 144 396 
rect 141 396 144 399 
rect 141 399 144 402 
rect 141 402 144 405 
rect 141 405 144 408 
rect 141 408 144 411 
rect 141 411 144 414 
rect 141 414 144 417 
rect 141 417 144 420 
rect 141 420 144 423 
rect 141 423 144 426 
rect 141 426 144 429 
rect 141 429 144 432 
rect 141 432 144 435 
rect 141 435 144 438 
rect 141 438 144 441 
rect 141 441 144 444 
rect 141 444 144 447 
rect 141 447 144 450 
rect 141 450 144 453 
rect 141 453 144 456 
rect 141 456 144 459 
rect 141 459 144 462 
rect 141 462 144 465 
rect 141 465 144 468 
rect 141 468 144 471 
rect 141 471 144 474 
rect 141 474 144 477 
rect 141 477 144 480 
rect 141 480 144 483 
rect 141 483 144 486 
rect 141 486 144 489 
rect 141 489 144 492 
rect 141 492 144 495 
rect 141 495 144 498 
rect 141 498 144 501 
rect 141 501 144 504 
rect 141 504 144 507 
rect 141 507 144 510 
rect 144 0 147 3 
rect 144 3 147 6 
rect 144 6 147 9 
rect 144 9 147 12 
rect 144 12 147 15 
rect 144 15 147 18 
rect 144 18 147 21 
rect 144 21 147 24 
rect 144 24 147 27 
rect 144 27 147 30 
rect 144 30 147 33 
rect 144 33 147 36 
rect 144 36 147 39 
rect 144 39 147 42 
rect 144 42 147 45 
rect 144 45 147 48 
rect 144 48 147 51 
rect 144 51 147 54 
rect 144 54 147 57 
rect 144 57 147 60 
rect 144 60 147 63 
rect 144 63 147 66 
rect 144 66 147 69 
rect 144 69 147 72 
rect 144 72 147 75 
rect 144 75 147 78 
rect 144 78 147 81 
rect 144 81 147 84 
rect 144 84 147 87 
rect 144 87 147 90 
rect 144 90 147 93 
rect 144 93 147 96 
rect 144 96 147 99 
rect 144 99 147 102 
rect 144 102 147 105 
rect 144 105 147 108 
rect 144 108 147 111 
rect 144 111 147 114 
rect 144 114 147 117 
rect 144 117 147 120 
rect 144 120 147 123 
rect 144 123 147 126 
rect 144 126 147 129 
rect 144 129 147 132 
rect 144 132 147 135 
rect 144 135 147 138 
rect 144 138 147 141 
rect 144 141 147 144 
rect 144 144 147 147 
rect 144 147 147 150 
rect 144 150 147 153 
rect 144 153 147 156 
rect 144 156 147 159 
rect 144 159 147 162 
rect 144 162 147 165 
rect 144 165 147 168 
rect 144 168 147 171 
rect 144 171 147 174 
rect 144 174 147 177 
rect 144 177 147 180 
rect 144 180 147 183 
rect 144 183 147 186 
rect 144 186 147 189 
rect 144 189 147 192 
rect 144 192 147 195 
rect 144 195 147 198 
rect 144 198 147 201 
rect 144 201 147 204 
rect 144 204 147 207 
rect 144 207 147 210 
rect 144 210 147 213 
rect 144 213 147 216 
rect 144 216 147 219 
rect 144 219 147 222 
rect 144 222 147 225 
rect 144 225 147 228 
rect 144 228 147 231 
rect 144 231 147 234 
rect 144 234 147 237 
rect 144 237 147 240 
rect 144 240 147 243 
rect 144 243 147 246 
rect 144 246 147 249 
rect 144 249 147 252 
rect 144 252 147 255 
rect 144 255 147 258 
rect 144 258 147 261 
rect 144 261 147 264 
rect 144 264 147 267 
rect 144 267 147 270 
rect 144 270 147 273 
rect 144 273 147 276 
rect 144 276 147 279 
rect 144 279 147 282 
rect 144 282 147 285 
rect 144 285 147 288 
rect 144 288 147 291 
rect 144 291 147 294 
rect 144 294 147 297 
rect 144 297 147 300 
rect 144 300 147 303 
rect 144 303 147 306 
rect 144 306 147 309 
rect 144 309 147 312 
rect 144 312 147 315 
rect 144 315 147 318 
rect 144 318 147 321 
rect 144 321 147 324 
rect 144 324 147 327 
rect 144 327 147 330 
rect 144 330 147 333 
rect 144 333 147 336 
rect 144 336 147 339 
rect 144 339 147 342 
rect 144 342 147 345 
rect 144 345 147 348 
rect 144 348 147 351 
rect 144 351 147 354 
rect 144 354 147 357 
rect 144 357 147 360 
rect 144 360 147 363 
rect 144 363 147 366 
rect 144 366 147 369 
rect 144 369 147 372 
rect 144 372 147 375 
rect 144 375 147 378 
rect 144 378 147 381 
rect 144 381 147 384 
rect 144 384 147 387 
rect 144 387 147 390 
rect 144 390 147 393 
rect 144 393 147 396 
rect 144 396 147 399 
rect 144 399 147 402 
rect 144 402 147 405 
rect 144 405 147 408 
rect 144 408 147 411 
rect 144 411 147 414 
rect 144 414 147 417 
rect 144 417 147 420 
rect 144 420 147 423 
rect 144 423 147 426 
rect 144 426 147 429 
rect 144 429 147 432 
rect 144 432 147 435 
rect 144 435 147 438 
rect 144 438 147 441 
rect 144 441 147 444 
rect 144 444 147 447 
rect 144 447 147 450 
rect 144 450 147 453 
rect 144 453 147 456 
rect 144 456 147 459 
rect 144 459 147 462 
rect 144 462 147 465 
rect 144 465 147 468 
rect 144 468 147 471 
rect 144 471 147 474 
rect 144 474 147 477 
rect 144 477 147 480 
rect 144 480 147 483 
rect 144 483 147 486 
rect 144 486 147 489 
rect 144 489 147 492 
rect 144 492 147 495 
rect 144 495 147 498 
rect 144 498 147 501 
rect 144 501 147 504 
rect 144 504 147 507 
rect 144 507 147 510 
rect 147 0 150 3 
rect 147 3 150 6 
rect 147 6 150 9 
rect 147 9 150 12 
rect 147 12 150 15 
rect 147 15 150 18 
rect 147 18 150 21 
rect 147 21 150 24 
rect 147 24 150 27 
rect 147 27 150 30 
rect 147 30 150 33 
rect 147 33 150 36 
rect 147 36 150 39 
rect 147 39 150 42 
rect 147 42 150 45 
rect 147 45 150 48 
rect 147 48 150 51 
rect 147 51 150 54 
rect 147 54 150 57 
rect 147 57 150 60 
rect 147 60 150 63 
rect 147 63 150 66 
rect 147 66 150 69 
rect 147 69 150 72 
rect 147 72 150 75 
rect 147 75 150 78 
rect 147 78 150 81 
rect 147 81 150 84 
rect 147 84 150 87 
rect 147 87 150 90 
rect 147 90 150 93 
rect 147 93 150 96 
rect 147 96 150 99 
rect 147 99 150 102 
rect 147 102 150 105 
rect 147 105 150 108 
rect 147 108 150 111 
rect 147 111 150 114 
rect 147 114 150 117 
rect 147 117 150 120 
rect 147 120 150 123 
rect 147 123 150 126 
rect 147 126 150 129 
rect 147 129 150 132 
rect 147 132 150 135 
rect 147 135 150 138 
rect 147 138 150 141 
rect 147 141 150 144 
rect 147 144 150 147 
rect 147 147 150 150 
rect 147 150 150 153 
rect 147 153 150 156 
rect 147 156 150 159 
rect 147 159 150 162 
rect 147 162 150 165 
rect 147 165 150 168 
rect 147 168 150 171 
rect 147 171 150 174 
rect 147 174 150 177 
rect 147 177 150 180 
rect 147 180 150 183 
rect 147 183 150 186 
rect 147 186 150 189 
rect 147 189 150 192 
rect 147 192 150 195 
rect 147 195 150 198 
rect 147 198 150 201 
rect 147 201 150 204 
rect 147 204 150 207 
rect 147 207 150 210 
rect 147 210 150 213 
rect 147 213 150 216 
rect 147 216 150 219 
rect 147 219 150 222 
rect 147 222 150 225 
rect 147 225 150 228 
rect 147 228 150 231 
rect 147 231 150 234 
rect 147 234 150 237 
rect 147 237 150 240 
rect 147 240 150 243 
rect 147 243 150 246 
rect 147 246 150 249 
rect 147 249 150 252 
rect 147 252 150 255 
rect 147 255 150 258 
rect 147 258 150 261 
rect 147 261 150 264 
rect 147 264 150 267 
rect 147 267 150 270 
rect 147 270 150 273 
rect 147 273 150 276 
rect 147 276 150 279 
rect 147 279 150 282 
rect 147 282 150 285 
rect 147 285 150 288 
rect 147 288 150 291 
rect 147 291 150 294 
rect 147 294 150 297 
rect 147 297 150 300 
rect 147 300 150 303 
rect 147 303 150 306 
rect 147 306 150 309 
rect 147 309 150 312 
rect 147 312 150 315 
rect 147 315 150 318 
rect 147 318 150 321 
rect 147 321 150 324 
rect 147 324 150 327 
rect 147 327 150 330 
rect 147 330 150 333 
rect 147 333 150 336 
rect 147 336 150 339 
rect 147 339 150 342 
rect 147 342 150 345 
rect 147 345 150 348 
rect 147 348 150 351 
rect 147 351 150 354 
rect 147 354 150 357 
rect 147 357 150 360 
rect 147 360 150 363 
rect 147 363 150 366 
rect 147 366 150 369 
rect 147 369 150 372 
rect 147 372 150 375 
rect 147 375 150 378 
rect 147 378 150 381 
rect 147 381 150 384 
rect 147 384 150 387 
rect 147 387 150 390 
rect 147 390 150 393 
rect 147 393 150 396 
rect 147 396 150 399 
rect 147 399 150 402 
rect 147 402 150 405 
rect 147 405 150 408 
rect 147 408 150 411 
rect 147 411 150 414 
rect 147 414 150 417 
rect 147 417 150 420 
rect 147 420 150 423 
rect 147 423 150 426 
rect 147 426 150 429 
rect 147 429 150 432 
rect 147 432 150 435 
rect 147 435 150 438 
rect 147 438 150 441 
rect 147 441 150 444 
rect 147 444 150 447 
rect 147 447 150 450 
rect 147 450 150 453 
rect 147 453 150 456 
rect 147 456 150 459 
rect 147 459 150 462 
rect 147 462 150 465 
rect 147 465 150 468 
rect 147 468 150 471 
rect 147 471 150 474 
rect 147 474 150 477 
rect 147 477 150 480 
rect 147 480 150 483 
rect 147 483 150 486 
rect 147 486 150 489 
rect 147 489 150 492 
rect 147 492 150 495 
rect 147 495 150 498 
rect 147 498 150 501 
rect 147 501 150 504 
rect 147 504 150 507 
rect 147 507 150 510 
rect 150 0 153 3 
rect 150 3 153 6 
rect 150 6 153 9 
rect 150 9 153 12 
rect 150 12 153 15 
rect 150 15 153 18 
rect 150 18 153 21 
rect 150 21 153 24 
rect 150 24 153 27 
rect 150 27 153 30 
rect 150 30 153 33 
rect 150 33 153 36 
rect 150 36 153 39 
rect 150 39 153 42 
rect 150 42 153 45 
rect 150 45 153 48 
rect 150 48 153 51 
rect 150 51 153 54 
rect 150 54 153 57 
rect 150 57 153 60 
rect 150 60 153 63 
rect 150 63 153 66 
rect 150 66 153 69 
rect 150 69 153 72 
rect 150 72 153 75 
rect 150 75 153 78 
rect 150 78 153 81 
rect 150 81 153 84 
rect 150 84 153 87 
rect 150 87 153 90 
rect 150 90 153 93 
rect 150 93 153 96 
rect 150 96 153 99 
rect 150 99 153 102 
rect 150 102 153 105 
rect 150 105 153 108 
rect 150 108 153 111 
rect 150 111 153 114 
rect 150 114 153 117 
rect 150 117 153 120 
rect 150 120 153 123 
rect 150 123 153 126 
rect 150 126 153 129 
rect 150 129 153 132 
rect 150 132 153 135 
rect 150 135 153 138 
rect 150 138 153 141 
rect 150 141 153 144 
rect 150 144 153 147 
rect 150 147 153 150 
rect 150 150 153 153 
rect 150 153 153 156 
rect 150 156 153 159 
rect 150 159 153 162 
rect 150 162 153 165 
rect 150 165 153 168 
rect 150 168 153 171 
rect 150 171 153 174 
rect 150 174 153 177 
rect 150 177 153 180 
rect 150 180 153 183 
rect 150 183 153 186 
rect 150 186 153 189 
rect 150 189 153 192 
rect 150 192 153 195 
rect 150 195 153 198 
rect 150 198 153 201 
rect 150 201 153 204 
rect 150 204 153 207 
rect 150 207 153 210 
rect 150 210 153 213 
rect 150 213 153 216 
rect 150 216 153 219 
rect 150 219 153 222 
rect 150 222 153 225 
rect 150 225 153 228 
rect 150 228 153 231 
rect 150 231 153 234 
rect 150 234 153 237 
rect 150 237 153 240 
rect 150 240 153 243 
rect 150 243 153 246 
rect 150 246 153 249 
rect 150 249 153 252 
rect 150 252 153 255 
rect 150 255 153 258 
rect 150 258 153 261 
rect 150 261 153 264 
rect 150 264 153 267 
rect 150 267 153 270 
rect 150 270 153 273 
rect 150 273 153 276 
rect 150 276 153 279 
rect 150 279 153 282 
rect 150 282 153 285 
rect 150 285 153 288 
rect 150 288 153 291 
rect 150 291 153 294 
rect 150 294 153 297 
rect 150 297 153 300 
rect 150 300 153 303 
rect 150 303 153 306 
rect 150 306 153 309 
rect 150 309 153 312 
rect 150 312 153 315 
rect 150 315 153 318 
rect 150 318 153 321 
rect 150 321 153 324 
rect 150 324 153 327 
rect 150 327 153 330 
rect 150 330 153 333 
rect 150 333 153 336 
rect 150 336 153 339 
rect 150 339 153 342 
rect 150 342 153 345 
rect 150 345 153 348 
rect 150 348 153 351 
rect 150 351 153 354 
rect 150 354 153 357 
rect 150 357 153 360 
rect 150 360 153 363 
rect 150 363 153 366 
rect 150 366 153 369 
rect 150 369 153 372 
rect 150 372 153 375 
rect 150 375 153 378 
rect 150 378 153 381 
rect 150 381 153 384 
rect 150 384 153 387 
rect 150 387 153 390 
rect 150 390 153 393 
rect 150 393 153 396 
rect 150 396 153 399 
rect 150 399 153 402 
rect 150 402 153 405 
rect 150 405 153 408 
rect 150 408 153 411 
rect 150 411 153 414 
rect 150 414 153 417 
rect 150 417 153 420 
rect 150 420 153 423 
rect 150 423 153 426 
rect 150 426 153 429 
rect 150 429 153 432 
rect 150 432 153 435 
rect 150 435 153 438 
rect 150 438 153 441 
rect 150 441 153 444 
rect 150 444 153 447 
rect 150 447 153 450 
rect 150 450 153 453 
rect 150 453 153 456 
rect 150 456 153 459 
rect 150 459 153 462 
rect 150 462 153 465 
rect 150 465 153 468 
rect 150 468 153 471 
rect 150 471 153 474 
rect 150 474 153 477 
rect 150 477 153 480 
rect 150 480 153 483 
rect 150 483 153 486 
rect 150 486 153 489 
rect 150 489 153 492 
rect 150 492 153 495 
rect 150 495 153 498 
rect 150 498 153 501 
rect 150 501 153 504 
rect 150 504 153 507 
rect 150 507 153 510 
rect 153 0 156 3 
rect 153 3 156 6 
rect 153 6 156 9 
rect 153 9 156 12 
rect 153 12 156 15 
rect 153 15 156 18 
rect 153 18 156 21 
rect 153 21 156 24 
rect 153 24 156 27 
rect 153 27 156 30 
rect 153 30 156 33 
rect 153 33 156 36 
rect 153 36 156 39 
rect 153 39 156 42 
rect 153 42 156 45 
rect 153 45 156 48 
rect 153 48 156 51 
rect 153 51 156 54 
rect 153 54 156 57 
rect 153 57 156 60 
rect 153 60 156 63 
rect 153 63 156 66 
rect 153 66 156 69 
rect 153 69 156 72 
rect 153 72 156 75 
rect 153 75 156 78 
rect 153 78 156 81 
rect 153 81 156 84 
rect 153 84 156 87 
rect 153 87 156 90 
rect 153 90 156 93 
rect 153 93 156 96 
rect 153 96 156 99 
rect 153 99 156 102 
rect 153 102 156 105 
rect 153 105 156 108 
rect 153 108 156 111 
rect 153 111 156 114 
rect 153 114 156 117 
rect 153 117 156 120 
rect 153 120 156 123 
rect 153 123 156 126 
rect 153 126 156 129 
rect 153 129 156 132 
rect 153 132 156 135 
rect 153 135 156 138 
rect 153 138 156 141 
rect 153 141 156 144 
rect 153 144 156 147 
rect 153 147 156 150 
rect 153 150 156 153 
rect 153 153 156 156 
rect 153 156 156 159 
rect 153 159 156 162 
rect 153 162 156 165 
rect 153 165 156 168 
rect 153 168 156 171 
rect 153 171 156 174 
rect 153 174 156 177 
rect 153 177 156 180 
rect 153 180 156 183 
rect 153 183 156 186 
rect 153 186 156 189 
rect 153 189 156 192 
rect 153 192 156 195 
rect 153 195 156 198 
rect 153 198 156 201 
rect 153 201 156 204 
rect 153 204 156 207 
rect 153 207 156 210 
rect 153 210 156 213 
rect 153 213 156 216 
rect 153 216 156 219 
rect 153 219 156 222 
rect 153 222 156 225 
rect 153 225 156 228 
rect 153 228 156 231 
rect 153 231 156 234 
rect 153 234 156 237 
rect 153 237 156 240 
rect 153 240 156 243 
rect 153 243 156 246 
rect 153 246 156 249 
rect 153 249 156 252 
rect 153 252 156 255 
rect 153 255 156 258 
rect 153 258 156 261 
rect 153 261 156 264 
rect 153 264 156 267 
rect 153 267 156 270 
rect 153 270 156 273 
rect 153 273 156 276 
rect 153 276 156 279 
rect 153 279 156 282 
rect 153 282 156 285 
rect 153 285 156 288 
rect 153 288 156 291 
rect 153 291 156 294 
rect 153 294 156 297 
rect 153 297 156 300 
rect 153 300 156 303 
rect 153 303 156 306 
rect 153 306 156 309 
rect 153 309 156 312 
rect 153 312 156 315 
rect 153 315 156 318 
rect 153 318 156 321 
rect 153 321 156 324 
rect 153 324 156 327 
rect 153 327 156 330 
rect 153 330 156 333 
rect 153 333 156 336 
rect 153 336 156 339 
rect 153 339 156 342 
rect 153 342 156 345 
rect 153 345 156 348 
rect 153 348 156 351 
rect 153 351 156 354 
rect 153 354 156 357 
rect 153 357 156 360 
rect 153 360 156 363 
rect 153 363 156 366 
rect 153 366 156 369 
rect 153 369 156 372 
rect 153 372 156 375 
rect 153 375 156 378 
rect 153 378 156 381 
rect 153 381 156 384 
rect 153 384 156 387 
rect 153 387 156 390 
rect 153 390 156 393 
rect 153 393 156 396 
rect 153 396 156 399 
rect 153 399 156 402 
rect 153 402 156 405 
rect 153 405 156 408 
rect 153 408 156 411 
rect 153 411 156 414 
rect 153 414 156 417 
rect 153 417 156 420 
rect 153 420 156 423 
rect 153 423 156 426 
rect 153 426 156 429 
rect 153 429 156 432 
rect 153 432 156 435 
rect 153 435 156 438 
rect 153 438 156 441 
rect 153 441 156 444 
rect 153 444 156 447 
rect 153 447 156 450 
rect 153 450 156 453 
rect 153 453 156 456 
rect 153 456 156 459 
rect 153 459 156 462 
rect 153 462 156 465 
rect 153 465 156 468 
rect 153 468 156 471 
rect 153 471 156 474 
rect 153 474 156 477 
rect 153 477 156 480 
rect 153 480 156 483 
rect 153 483 156 486 
rect 153 486 156 489 
rect 153 489 156 492 
rect 153 492 156 495 
rect 153 495 156 498 
rect 153 498 156 501 
rect 153 501 156 504 
rect 153 504 156 507 
rect 153 507 156 510 
rect 156 0 159 3 
rect 156 3 159 6 
rect 156 6 159 9 
rect 156 9 159 12 
rect 156 12 159 15 
rect 156 15 159 18 
rect 156 18 159 21 
rect 156 21 159 24 
rect 156 24 159 27 
rect 156 27 159 30 
rect 156 30 159 33 
rect 156 33 159 36 
rect 156 36 159 39 
rect 156 39 159 42 
rect 156 42 159 45 
rect 156 45 159 48 
rect 156 48 159 51 
rect 156 51 159 54 
rect 156 54 159 57 
rect 156 57 159 60 
rect 156 60 159 63 
rect 156 63 159 66 
rect 156 66 159 69 
rect 156 69 159 72 
rect 156 72 159 75 
rect 156 75 159 78 
rect 156 78 159 81 
rect 156 81 159 84 
rect 156 84 159 87 
rect 156 87 159 90 
rect 156 90 159 93 
rect 156 93 159 96 
rect 156 96 159 99 
rect 156 99 159 102 
rect 156 102 159 105 
rect 156 105 159 108 
rect 156 108 159 111 
rect 156 111 159 114 
rect 156 114 159 117 
rect 156 117 159 120 
rect 156 120 159 123 
rect 156 123 159 126 
rect 156 126 159 129 
rect 156 129 159 132 
rect 156 132 159 135 
rect 156 135 159 138 
rect 156 138 159 141 
rect 156 141 159 144 
rect 156 144 159 147 
rect 156 147 159 150 
rect 156 150 159 153 
rect 156 153 159 156 
rect 156 156 159 159 
rect 156 159 159 162 
rect 156 162 159 165 
rect 156 165 159 168 
rect 156 168 159 171 
rect 156 171 159 174 
rect 156 174 159 177 
rect 156 177 159 180 
rect 156 180 159 183 
rect 156 183 159 186 
rect 156 186 159 189 
rect 156 189 159 192 
rect 156 192 159 195 
rect 156 195 159 198 
rect 156 198 159 201 
rect 156 201 159 204 
rect 156 204 159 207 
rect 156 207 159 210 
rect 156 210 159 213 
rect 156 213 159 216 
rect 156 216 159 219 
rect 156 219 159 222 
rect 156 222 159 225 
rect 156 225 159 228 
rect 156 228 159 231 
rect 156 231 159 234 
rect 156 234 159 237 
rect 156 237 159 240 
rect 156 240 159 243 
rect 156 243 159 246 
rect 156 246 159 249 
rect 156 249 159 252 
rect 156 252 159 255 
rect 156 255 159 258 
rect 156 258 159 261 
rect 156 261 159 264 
rect 156 264 159 267 
rect 156 267 159 270 
rect 156 270 159 273 
rect 156 273 159 276 
rect 156 276 159 279 
rect 156 279 159 282 
rect 156 282 159 285 
rect 156 285 159 288 
rect 156 288 159 291 
rect 156 291 159 294 
rect 156 294 159 297 
rect 156 297 159 300 
rect 156 300 159 303 
rect 156 303 159 306 
rect 156 306 159 309 
rect 156 309 159 312 
rect 156 312 159 315 
rect 156 315 159 318 
rect 156 318 159 321 
rect 156 321 159 324 
rect 156 324 159 327 
rect 156 327 159 330 
rect 156 330 159 333 
rect 156 333 159 336 
rect 156 336 159 339 
rect 156 339 159 342 
rect 156 342 159 345 
rect 156 345 159 348 
rect 156 348 159 351 
rect 156 351 159 354 
rect 156 354 159 357 
rect 156 357 159 360 
rect 156 360 159 363 
rect 156 363 159 366 
rect 156 366 159 369 
rect 156 369 159 372 
rect 156 372 159 375 
rect 156 375 159 378 
rect 156 378 159 381 
rect 156 381 159 384 
rect 156 384 159 387 
rect 156 387 159 390 
rect 156 390 159 393 
rect 156 393 159 396 
rect 156 396 159 399 
rect 156 399 159 402 
rect 156 402 159 405 
rect 156 405 159 408 
rect 156 408 159 411 
rect 156 411 159 414 
rect 156 414 159 417 
rect 156 417 159 420 
rect 156 420 159 423 
rect 156 423 159 426 
rect 156 426 159 429 
rect 156 429 159 432 
rect 156 432 159 435 
rect 156 435 159 438 
rect 156 438 159 441 
rect 156 441 159 444 
rect 156 444 159 447 
rect 156 447 159 450 
rect 156 450 159 453 
rect 156 453 159 456 
rect 156 456 159 459 
rect 156 459 159 462 
rect 156 462 159 465 
rect 156 465 159 468 
rect 156 468 159 471 
rect 156 471 159 474 
rect 156 474 159 477 
rect 156 477 159 480 
rect 156 480 159 483 
rect 156 483 159 486 
rect 156 486 159 489 
rect 156 489 159 492 
rect 156 492 159 495 
rect 156 495 159 498 
rect 156 498 159 501 
rect 156 501 159 504 
rect 156 504 159 507 
rect 156 507 159 510 
rect 159 0 162 3 
rect 159 3 162 6 
rect 159 6 162 9 
rect 159 9 162 12 
rect 159 12 162 15 
rect 159 15 162 18 
rect 159 18 162 21 
rect 159 21 162 24 
rect 159 24 162 27 
rect 159 27 162 30 
rect 159 30 162 33 
rect 159 33 162 36 
rect 159 36 162 39 
rect 159 39 162 42 
rect 159 42 162 45 
rect 159 45 162 48 
rect 159 48 162 51 
rect 159 51 162 54 
rect 159 54 162 57 
rect 159 57 162 60 
rect 159 60 162 63 
rect 159 63 162 66 
rect 159 66 162 69 
rect 159 69 162 72 
rect 159 72 162 75 
rect 159 75 162 78 
rect 159 78 162 81 
rect 159 81 162 84 
rect 159 84 162 87 
rect 159 87 162 90 
rect 159 90 162 93 
rect 159 93 162 96 
rect 159 96 162 99 
rect 159 99 162 102 
rect 159 102 162 105 
rect 159 105 162 108 
rect 159 108 162 111 
rect 159 111 162 114 
rect 159 114 162 117 
rect 159 117 162 120 
rect 159 120 162 123 
rect 159 123 162 126 
rect 159 126 162 129 
rect 159 129 162 132 
rect 159 132 162 135 
rect 159 135 162 138 
rect 159 138 162 141 
rect 159 141 162 144 
rect 159 144 162 147 
rect 159 147 162 150 
rect 159 150 162 153 
rect 159 153 162 156 
rect 159 156 162 159 
rect 159 159 162 162 
rect 159 162 162 165 
rect 159 165 162 168 
rect 159 168 162 171 
rect 159 171 162 174 
rect 159 174 162 177 
rect 159 177 162 180 
rect 159 180 162 183 
rect 159 183 162 186 
rect 159 186 162 189 
rect 159 189 162 192 
rect 159 192 162 195 
rect 159 195 162 198 
rect 159 198 162 201 
rect 159 201 162 204 
rect 159 204 162 207 
rect 159 207 162 210 
rect 159 210 162 213 
rect 159 213 162 216 
rect 159 216 162 219 
rect 159 219 162 222 
rect 159 222 162 225 
rect 159 225 162 228 
rect 159 228 162 231 
rect 159 231 162 234 
rect 159 234 162 237 
rect 159 237 162 240 
rect 159 240 162 243 
rect 159 243 162 246 
rect 159 246 162 249 
rect 159 249 162 252 
rect 159 252 162 255 
rect 159 255 162 258 
rect 159 258 162 261 
rect 159 261 162 264 
rect 159 264 162 267 
rect 159 267 162 270 
rect 159 270 162 273 
rect 159 273 162 276 
rect 159 276 162 279 
rect 159 279 162 282 
rect 159 282 162 285 
rect 159 285 162 288 
rect 159 288 162 291 
rect 159 291 162 294 
rect 159 294 162 297 
rect 159 297 162 300 
rect 159 300 162 303 
rect 159 303 162 306 
rect 159 306 162 309 
rect 159 309 162 312 
rect 159 312 162 315 
rect 159 315 162 318 
rect 159 318 162 321 
rect 159 321 162 324 
rect 159 324 162 327 
rect 159 327 162 330 
rect 159 330 162 333 
rect 159 333 162 336 
rect 159 336 162 339 
rect 159 339 162 342 
rect 159 342 162 345 
rect 159 345 162 348 
rect 159 348 162 351 
rect 159 351 162 354 
rect 159 354 162 357 
rect 159 357 162 360 
rect 159 360 162 363 
rect 159 363 162 366 
rect 159 366 162 369 
rect 159 369 162 372 
rect 159 372 162 375 
rect 159 375 162 378 
rect 159 378 162 381 
rect 159 381 162 384 
rect 159 384 162 387 
rect 159 387 162 390 
rect 159 390 162 393 
rect 159 393 162 396 
rect 159 396 162 399 
rect 159 399 162 402 
rect 159 402 162 405 
rect 159 405 162 408 
rect 159 408 162 411 
rect 159 411 162 414 
rect 159 414 162 417 
rect 159 417 162 420 
rect 159 420 162 423 
rect 159 423 162 426 
rect 159 426 162 429 
rect 159 429 162 432 
rect 159 432 162 435 
rect 159 435 162 438 
rect 159 438 162 441 
rect 159 441 162 444 
rect 159 444 162 447 
rect 159 447 162 450 
rect 159 450 162 453 
rect 159 453 162 456 
rect 159 456 162 459 
rect 159 459 162 462 
rect 159 462 162 465 
rect 159 465 162 468 
rect 159 468 162 471 
rect 159 471 162 474 
rect 159 474 162 477 
rect 159 477 162 480 
rect 159 480 162 483 
rect 159 483 162 486 
rect 159 486 162 489 
rect 159 489 162 492 
rect 159 492 162 495 
rect 159 495 162 498 
rect 159 498 162 501 
rect 159 501 162 504 
rect 159 504 162 507 
rect 159 507 162 510 
rect 162 0 165 3 
rect 162 3 165 6 
rect 162 6 165 9 
rect 162 9 165 12 
rect 162 12 165 15 
rect 162 15 165 18 
rect 162 18 165 21 
rect 162 21 165 24 
rect 162 24 165 27 
rect 162 27 165 30 
rect 162 30 165 33 
rect 162 33 165 36 
rect 162 36 165 39 
rect 162 39 165 42 
rect 162 42 165 45 
rect 162 45 165 48 
rect 162 48 165 51 
rect 162 51 165 54 
rect 162 54 165 57 
rect 162 57 165 60 
rect 162 60 165 63 
rect 162 63 165 66 
rect 162 66 165 69 
rect 162 69 165 72 
rect 162 72 165 75 
rect 162 75 165 78 
rect 162 78 165 81 
rect 162 81 165 84 
rect 162 84 165 87 
rect 162 87 165 90 
rect 162 90 165 93 
rect 162 93 165 96 
rect 162 96 165 99 
rect 162 99 165 102 
rect 162 102 165 105 
rect 162 105 165 108 
rect 162 108 165 111 
rect 162 111 165 114 
rect 162 114 165 117 
rect 162 117 165 120 
rect 162 120 165 123 
rect 162 123 165 126 
rect 162 126 165 129 
rect 162 129 165 132 
rect 162 132 165 135 
rect 162 135 165 138 
rect 162 138 165 141 
rect 162 141 165 144 
rect 162 144 165 147 
rect 162 147 165 150 
rect 162 150 165 153 
rect 162 153 165 156 
rect 162 156 165 159 
rect 162 159 165 162 
rect 162 162 165 165 
rect 162 165 165 168 
rect 162 168 165 171 
rect 162 171 165 174 
rect 162 174 165 177 
rect 162 177 165 180 
rect 162 180 165 183 
rect 162 183 165 186 
rect 162 186 165 189 
rect 162 189 165 192 
rect 162 192 165 195 
rect 162 195 165 198 
rect 162 198 165 201 
rect 162 201 165 204 
rect 162 204 165 207 
rect 162 207 165 210 
rect 162 210 165 213 
rect 162 213 165 216 
rect 162 216 165 219 
rect 162 219 165 222 
rect 162 222 165 225 
rect 162 225 165 228 
rect 162 228 165 231 
rect 162 231 165 234 
rect 162 234 165 237 
rect 162 237 165 240 
rect 162 240 165 243 
rect 162 243 165 246 
rect 162 246 165 249 
rect 162 249 165 252 
rect 162 252 165 255 
rect 162 255 165 258 
rect 162 258 165 261 
rect 162 261 165 264 
rect 162 264 165 267 
rect 162 267 165 270 
rect 162 270 165 273 
rect 162 273 165 276 
rect 162 276 165 279 
rect 162 279 165 282 
rect 162 282 165 285 
rect 162 285 165 288 
rect 162 288 165 291 
rect 162 291 165 294 
rect 162 294 165 297 
rect 162 297 165 300 
rect 162 300 165 303 
rect 162 303 165 306 
rect 162 306 165 309 
rect 162 309 165 312 
rect 162 312 165 315 
rect 162 315 165 318 
rect 162 318 165 321 
rect 162 321 165 324 
rect 162 324 165 327 
rect 162 327 165 330 
rect 162 330 165 333 
rect 162 333 165 336 
rect 162 336 165 339 
rect 162 339 165 342 
rect 162 342 165 345 
rect 162 345 165 348 
rect 162 348 165 351 
rect 162 351 165 354 
rect 162 354 165 357 
rect 162 357 165 360 
rect 162 360 165 363 
rect 162 363 165 366 
rect 162 366 165 369 
rect 162 369 165 372 
rect 162 372 165 375 
rect 162 375 165 378 
rect 162 378 165 381 
rect 162 381 165 384 
rect 162 384 165 387 
rect 162 387 165 390 
rect 162 390 165 393 
rect 162 393 165 396 
rect 162 396 165 399 
rect 162 399 165 402 
rect 162 402 165 405 
rect 162 405 165 408 
rect 162 408 165 411 
rect 162 411 165 414 
rect 162 414 165 417 
rect 162 417 165 420 
rect 162 420 165 423 
rect 162 423 165 426 
rect 162 426 165 429 
rect 162 429 165 432 
rect 162 432 165 435 
rect 162 435 165 438 
rect 162 438 165 441 
rect 162 441 165 444 
rect 162 444 165 447 
rect 162 447 165 450 
rect 162 450 165 453 
rect 162 453 165 456 
rect 162 456 165 459 
rect 162 459 165 462 
rect 162 462 165 465 
rect 162 465 165 468 
rect 162 468 165 471 
rect 162 471 165 474 
rect 162 474 165 477 
rect 162 477 165 480 
rect 162 480 165 483 
rect 162 483 165 486 
rect 162 486 165 489 
rect 162 489 165 492 
rect 162 492 165 495 
rect 162 495 165 498 
rect 162 498 165 501 
rect 162 501 165 504 
rect 162 504 165 507 
rect 162 507 165 510 
rect 165 0 168 3 
rect 165 3 168 6 
rect 165 6 168 9 
rect 165 9 168 12 
rect 165 12 168 15 
rect 165 15 168 18 
rect 165 18 168 21 
rect 165 21 168 24 
rect 165 24 168 27 
rect 165 27 168 30 
rect 165 30 168 33 
rect 165 33 168 36 
rect 165 36 168 39 
rect 165 39 168 42 
rect 165 42 168 45 
rect 165 45 168 48 
rect 165 48 168 51 
rect 165 51 168 54 
rect 165 54 168 57 
rect 165 57 168 60 
rect 165 60 168 63 
rect 165 63 168 66 
rect 165 66 168 69 
rect 165 69 168 72 
rect 165 72 168 75 
rect 165 75 168 78 
rect 165 78 168 81 
rect 165 81 168 84 
rect 165 84 168 87 
rect 165 87 168 90 
rect 165 90 168 93 
rect 165 93 168 96 
rect 165 96 168 99 
rect 165 99 168 102 
rect 165 102 168 105 
rect 165 105 168 108 
rect 165 108 168 111 
rect 165 111 168 114 
rect 165 114 168 117 
rect 165 117 168 120 
rect 165 120 168 123 
rect 165 123 168 126 
rect 165 126 168 129 
rect 165 129 168 132 
rect 165 132 168 135 
rect 165 135 168 138 
rect 165 138 168 141 
rect 165 141 168 144 
rect 165 144 168 147 
rect 165 147 168 150 
rect 165 150 168 153 
rect 165 153 168 156 
rect 165 156 168 159 
rect 165 159 168 162 
rect 165 162 168 165 
rect 165 165 168 168 
rect 165 168 168 171 
rect 165 171 168 174 
rect 165 174 168 177 
rect 165 177 168 180 
rect 165 180 168 183 
rect 165 183 168 186 
rect 165 186 168 189 
rect 165 189 168 192 
rect 165 192 168 195 
rect 165 195 168 198 
rect 165 198 168 201 
rect 165 201 168 204 
rect 165 204 168 207 
rect 165 207 168 210 
rect 165 210 168 213 
rect 165 213 168 216 
rect 165 216 168 219 
rect 165 219 168 222 
rect 165 222 168 225 
rect 165 225 168 228 
rect 165 228 168 231 
rect 165 231 168 234 
rect 165 234 168 237 
rect 165 237 168 240 
rect 165 240 168 243 
rect 165 243 168 246 
rect 165 246 168 249 
rect 165 249 168 252 
rect 165 252 168 255 
rect 165 255 168 258 
rect 165 258 168 261 
rect 165 261 168 264 
rect 165 264 168 267 
rect 165 267 168 270 
rect 165 270 168 273 
rect 165 273 168 276 
rect 165 276 168 279 
rect 165 279 168 282 
rect 165 282 168 285 
rect 165 285 168 288 
rect 165 288 168 291 
rect 165 291 168 294 
rect 165 294 168 297 
rect 165 297 168 300 
rect 165 300 168 303 
rect 165 303 168 306 
rect 165 306 168 309 
rect 165 309 168 312 
rect 165 312 168 315 
rect 165 315 168 318 
rect 165 318 168 321 
rect 165 321 168 324 
rect 165 324 168 327 
rect 165 327 168 330 
rect 165 330 168 333 
rect 165 333 168 336 
rect 165 336 168 339 
rect 165 339 168 342 
rect 165 342 168 345 
rect 165 345 168 348 
rect 165 348 168 351 
rect 165 351 168 354 
rect 165 354 168 357 
rect 165 357 168 360 
rect 165 360 168 363 
rect 165 363 168 366 
rect 165 366 168 369 
rect 165 369 168 372 
rect 165 372 168 375 
rect 165 375 168 378 
rect 165 378 168 381 
rect 165 381 168 384 
rect 165 384 168 387 
rect 165 387 168 390 
rect 165 390 168 393 
rect 165 393 168 396 
rect 165 396 168 399 
rect 165 399 168 402 
rect 165 402 168 405 
rect 165 405 168 408 
rect 165 408 168 411 
rect 165 411 168 414 
rect 165 414 168 417 
rect 165 417 168 420 
rect 165 420 168 423 
rect 165 423 168 426 
rect 165 426 168 429 
rect 165 429 168 432 
rect 165 432 168 435 
rect 165 435 168 438 
rect 165 438 168 441 
rect 165 441 168 444 
rect 165 444 168 447 
rect 165 447 168 450 
rect 165 450 168 453 
rect 165 453 168 456 
rect 165 456 168 459 
rect 165 459 168 462 
rect 165 462 168 465 
rect 165 465 168 468 
rect 165 468 168 471 
rect 165 471 168 474 
rect 165 474 168 477 
rect 165 477 168 480 
rect 165 480 168 483 
rect 165 483 168 486 
rect 165 486 168 489 
rect 165 489 168 492 
rect 165 492 168 495 
rect 165 495 168 498 
rect 165 498 168 501 
rect 165 501 168 504 
rect 165 504 168 507 
rect 165 507 168 510 
rect 168 0 171 3 
rect 168 3 171 6 
rect 168 6 171 9 
rect 168 9 171 12 
rect 168 12 171 15 
rect 168 15 171 18 
rect 168 18 171 21 
rect 168 21 171 24 
rect 168 24 171 27 
rect 168 27 171 30 
rect 168 30 171 33 
rect 168 33 171 36 
rect 168 36 171 39 
rect 168 39 171 42 
rect 168 42 171 45 
rect 168 45 171 48 
rect 168 48 171 51 
rect 168 51 171 54 
rect 168 54 171 57 
rect 168 57 171 60 
rect 168 60 171 63 
rect 168 63 171 66 
rect 168 66 171 69 
rect 168 69 171 72 
rect 168 72 171 75 
rect 168 75 171 78 
rect 168 78 171 81 
rect 168 81 171 84 
rect 168 84 171 87 
rect 168 87 171 90 
rect 168 90 171 93 
rect 168 93 171 96 
rect 168 96 171 99 
rect 168 99 171 102 
rect 168 102 171 105 
rect 168 105 171 108 
rect 168 108 171 111 
rect 168 111 171 114 
rect 168 114 171 117 
rect 168 117 171 120 
rect 168 120 171 123 
rect 168 123 171 126 
rect 168 126 171 129 
rect 168 129 171 132 
rect 168 132 171 135 
rect 168 135 171 138 
rect 168 138 171 141 
rect 168 141 171 144 
rect 168 144 171 147 
rect 168 147 171 150 
rect 168 150 171 153 
rect 168 153 171 156 
rect 168 156 171 159 
rect 168 159 171 162 
rect 168 162 171 165 
rect 168 165 171 168 
rect 168 168 171 171 
rect 168 171 171 174 
rect 168 174 171 177 
rect 168 177 171 180 
rect 168 180 171 183 
rect 168 183 171 186 
rect 168 186 171 189 
rect 168 189 171 192 
rect 168 192 171 195 
rect 168 195 171 198 
rect 168 198 171 201 
rect 168 201 171 204 
rect 168 204 171 207 
rect 168 207 171 210 
rect 168 210 171 213 
rect 168 213 171 216 
rect 168 216 171 219 
rect 168 219 171 222 
rect 168 222 171 225 
rect 168 225 171 228 
rect 168 228 171 231 
rect 168 231 171 234 
rect 168 234 171 237 
rect 168 237 171 240 
rect 168 240 171 243 
rect 168 243 171 246 
rect 168 246 171 249 
rect 168 249 171 252 
rect 168 252 171 255 
rect 168 255 171 258 
rect 168 258 171 261 
rect 168 261 171 264 
rect 168 264 171 267 
rect 168 267 171 270 
rect 168 270 171 273 
rect 168 273 171 276 
rect 168 276 171 279 
rect 168 279 171 282 
rect 168 282 171 285 
rect 168 285 171 288 
rect 168 288 171 291 
rect 168 291 171 294 
rect 168 294 171 297 
rect 168 297 171 300 
rect 168 300 171 303 
rect 168 303 171 306 
rect 168 306 171 309 
rect 168 309 171 312 
rect 168 312 171 315 
rect 168 315 171 318 
rect 168 318 171 321 
rect 168 321 171 324 
rect 168 324 171 327 
rect 168 327 171 330 
rect 168 330 171 333 
rect 168 333 171 336 
rect 168 336 171 339 
rect 168 339 171 342 
rect 168 342 171 345 
rect 168 345 171 348 
rect 168 348 171 351 
rect 168 351 171 354 
rect 168 354 171 357 
rect 168 357 171 360 
rect 168 360 171 363 
rect 168 363 171 366 
rect 168 366 171 369 
rect 168 369 171 372 
rect 168 372 171 375 
rect 168 375 171 378 
rect 168 378 171 381 
rect 168 381 171 384 
rect 168 384 171 387 
rect 168 387 171 390 
rect 168 390 171 393 
rect 168 393 171 396 
rect 168 396 171 399 
rect 168 399 171 402 
rect 168 402 171 405 
rect 168 405 171 408 
rect 168 408 171 411 
rect 168 411 171 414 
rect 168 414 171 417 
rect 168 417 171 420 
rect 168 420 171 423 
rect 168 423 171 426 
rect 168 426 171 429 
rect 168 429 171 432 
rect 168 432 171 435 
rect 168 435 171 438 
rect 168 438 171 441 
rect 168 441 171 444 
rect 168 444 171 447 
rect 168 447 171 450 
rect 168 450 171 453 
rect 168 453 171 456 
rect 168 456 171 459 
rect 168 459 171 462 
rect 168 462 171 465 
rect 168 465 171 468 
rect 168 468 171 471 
rect 168 471 171 474 
rect 168 474 171 477 
rect 168 477 171 480 
rect 168 480 171 483 
rect 168 483 171 486 
rect 168 486 171 489 
rect 168 489 171 492 
rect 168 492 171 495 
rect 168 495 171 498 
rect 168 498 171 501 
rect 168 501 171 504 
rect 168 504 171 507 
rect 168 507 171 510 
rect 171 0 174 3 
rect 171 3 174 6 
rect 171 6 174 9 
rect 171 9 174 12 
rect 171 12 174 15 
rect 171 15 174 18 
rect 171 18 174 21 
rect 171 21 174 24 
rect 171 24 174 27 
rect 171 27 174 30 
rect 171 30 174 33 
rect 171 33 174 36 
rect 171 36 174 39 
rect 171 39 174 42 
rect 171 42 174 45 
rect 171 45 174 48 
rect 171 48 174 51 
rect 171 51 174 54 
rect 171 54 174 57 
rect 171 57 174 60 
rect 171 60 174 63 
rect 171 63 174 66 
rect 171 66 174 69 
rect 171 69 174 72 
rect 171 72 174 75 
rect 171 75 174 78 
rect 171 78 174 81 
rect 171 81 174 84 
rect 171 84 174 87 
rect 171 87 174 90 
rect 171 90 174 93 
rect 171 93 174 96 
rect 171 96 174 99 
rect 171 99 174 102 
rect 171 102 174 105 
rect 171 105 174 108 
rect 171 108 174 111 
rect 171 111 174 114 
rect 171 114 174 117 
rect 171 117 174 120 
rect 171 120 174 123 
rect 171 123 174 126 
rect 171 126 174 129 
rect 171 129 174 132 
rect 171 132 174 135 
rect 171 135 174 138 
rect 171 138 174 141 
rect 171 141 174 144 
rect 171 144 174 147 
rect 171 147 174 150 
rect 171 150 174 153 
rect 171 153 174 156 
rect 171 156 174 159 
rect 171 159 174 162 
rect 171 162 174 165 
rect 171 165 174 168 
rect 171 168 174 171 
rect 171 171 174 174 
rect 171 174 174 177 
rect 171 177 174 180 
rect 171 180 174 183 
rect 171 183 174 186 
rect 171 186 174 189 
rect 171 189 174 192 
rect 171 192 174 195 
rect 171 195 174 198 
rect 171 198 174 201 
rect 171 201 174 204 
rect 171 204 174 207 
rect 171 207 174 210 
rect 171 210 174 213 
rect 171 213 174 216 
rect 171 216 174 219 
rect 171 219 174 222 
rect 171 222 174 225 
rect 171 225 174 228 
rect 171 228 174 231 
rect 171 231 174 234 
rect 171 234 174 237 
rect 171 237 174 240 
rect 171 240 174 243 
rect 171 243 174 246 
rect 171 246 174 249 
rect 171 249 174 252 
rect 171 252 174 255 
rect 171 255 174 258 
rect 171 258 174 261 
rect 171 261 174 264 
rect 171 264 174 267 
rect 171 267 174 270 
rect 171 270 174 273 
rect 171 273 174 276 
rect 171 276 174 279 
rect 171 279 174 282 
rect 171 282 174 285 
rect 171 285 174 288 
rect 171 288 174 291 
rect 171 291 174 294 
rect 171 294 174 297 
rect 171 297 174 300 
rect 171 300 174 303 
rect 171 303 174 306 
rect 171 306 174 309 
rect 171 309 174 312 
rect 171 312 174 315 
rect 171 315 174 318 
rect 171 318 174 321 
rect 171 321 174 324 
rect 171 324 174 327 
rect 171 327 174 330 
rect 171 330 174 333 
rect 171 333 174 336 
rect 171 336 174 339 
rect 171 339 174 342 
rect 171 342 174 345 
rect 171 345 174 348 
rect 171 348 174 351 
rect 171 351 174 354 
rect 171 354 174 357 
rect 171 357 174 360 
rect 171 360 174 363 
rect 171 363 174 366 
rect 171 366 174 369 
rect 171 369 174 372 
rect 171 372 174 375 
rect 171 375 174 378 
rect 171 378 174 381 
rect 171 381 174 384 
rect 171 384 174 387 
rect 171 387 174 390 
rect 171 390 174 393 
rect 171 393 174 396 
rect 171 396 174 399 
rect 171 399 174 402 
rect 171 402 174 405 
rect 171 405 174 408 
rect 171 408 174 411 
rect 171 411 174 414 
rect 171 414 174 417 
rect 171 417 174 420 
rect 171 420 174 423 
rect 171 423 174 426 
rect 171 426 174 429 
rect 171 429 174 432 
rect 171 432 174 435 
rect 171 435 174 438 
rect 171 438 174 441 
rect 171 441 174 444 
rect 171 444 174 447 
rect 171 447 174 450 
rect 171 450 174 453 
rect 171 453 174 456 
rect 171 456 174 459 
rect 171 459 174 462 
rect 171 462 174 465 
rect 171 465 174 468 
rect 171 468 174 471 
rect 171 471 174 474 
rect 171 474 174 477 
rect 171 477 174 480 
rect 171 480 174 483 
rect 171 483 174 486 
rect 171 486 174 489 
rect 171 489 174 492 
rect 171 492 174 495 
rect 171 495 174 498 
rect 171 498 174 501 
rect 171 501 174 504 
rect 171 504 174 507 
rect 171 507 174 510 
rect 174 0 177 3 
rect 174 3 177 6 
rect 174 6 177 9 
rect 174 9 177 12 
rect 174 12 177 15 
rect 174 15 177 18 
rect 174 18 177 21 
rect 174 21 177 24 
rect 174 24 177 27 
rect 174 27 177 30 
rect 174 30 177 33 
rect 174 33 177 36 
rect 174 36 177 39 
rect 174 39 177 42 
rect 174 42 177 45 
rect 174 45 177 48 
rect 174 48 177 51 
rect 174 51 177 54 
rect 174 54 177 57 
rect 174 57 177 60 
rect 174 60 177 63 
rect 174 63 177 66 
rect 174 66 177 69 
rect 174 69 177 72 
rect 174 72 177 75 
rect 174 75 177 78 
rect 174 78 177 81 
rect 174 81 177 84 
rect 174 84 177 87 
rect 174 87 177 90 
rect 174 90 177 93 
rect 174 93 177 96 
rect 174 96 177 99 
rect 174 99 177 102 
rect 174 102 177 105 
rect 174 105 177 108 
rect 174 108 177 111 
rect 174 111 177 114 
rect 174 114 177 117 
rect 174 117 177 120 
rect 174 120 177 123 
rect 174 123 177 126 
rect 174 126 177 129 
rect 174 129 177 132 
rect 174 132 177 135 
rect 174 135 177 138 
rect 174 138 177 141 
rect 174 141 177 144 
rect 174 144 177 147 
rect 174 147 177 150 
rect 174 150 177 153 
rect 174 153 177 156 
rect 174 156 177 159 
rect 174 159 177 162 
rect 174 162 177 165 
rect 174 165 177 168 
rect 174 168 177 171 
rect 174 171 177 174 
rect 174 174 177 177 
rect 174 177 177 180 
rect 174 180 177 183 
rect 174 183 177 186 
rect 174 186 177 189 
rect 174 189 177 192 
rect 174 192 177 195 
rect 174 195 177 198 
rect 174 198 177 201 
rect 174 201 177 204 
rect 174 204 177 207 
rect 174 207 177 210 
rect 174 210 177 213 
rect 174 213 177 216 
rect 174 216 177 219 
rect 174 219 177 222 
rect 174 222 177 225 
rect 174 225 177 228 
rect 174 228 177 231 
rect 174 231 177 234 
rect 174 234 177 237 
rect 174 237 177 240 
rect 174 240 177 243 
rect 174 243 177 246 
rect 174 246 177 249 
rect 174 249 177 252 
rect 174 252 177 255 
rect 174 255 177 258 
rect 174 258 177 261 
rect 174 261 177 264 
rect 174 264 177 267 
rect 174 267 177 270 
rect 174 270 177 273 
rect 174 273 177 276 
rect 174 276 177 279 
rect 174 279 177 282 
rect 174 282 177 285 
rect 174 285 177 288 
rect 174 288 177 291 
rect 174 291 177 294 
rect 174 294 177 297 
rect 174 297 177 300 
rect 174 300 177 303 
rect 174 303 177 306 
rect 174 306 177 309 
rect 174 309 177 312 
rect 174 312 177 315 
rect 174 315 177 318 
rect 174 318 177 321 
rect 174 321 177 324 
rect 174 324 177 327 
rect 174 327 177 330 
rect 174 330 177 333 
rect 174 333 177 336 
rect 174 336 177 339 
rect 174 339 177 342 
rect 174 342 177 345 
rect 174 345 177 348 
rect 174 348 177 351 
rect 174 351 177 354 
rect 174 354 177 357 
rect 174 357 177 360 
rect 174 360 177 363 
rect 174 363 177 366 
rect 174 366 177 369 
rect 174 369 177 372 
rect 174 372 177 375 
rect 174 375 177 378 
rect 174 378 177 381 
rect 174 381 177 384 
rect 174 384 177 387 
rect 174 387 177 390 
rect 174 390 177 393 
rect 174 393 177 396 
rect 174 396 177 399 
rect 174 399 177 402 
rect 174 402 177 405 
rect 174 405 177 408 
rect 174 408 177 411 
rect 174 411 177 414 
rect 174 414 177 417 
rect 174 417 177 420 
rect 174 420 177 423 
rect 174 423 177 426 
rect 174 426 177 429 
rect 174 429 177 432 
rect 174 432 177 435 
rect 174 435 177 438 
rect 174 438 177 441 
rect 174 441 177 444 
rect 174 444 177 447 
rect 174 447 177 450 
rect 174 450 177 453 
rect 174 453 177 456 
rect 174 456 177 459 
rect 174 459 177 462 
rect 174 462 177 465 
rect 174 465 177 468 
rect 174 468 177 471 
rect 174 471 177 474 
rect 174 474 177 477 
rect 174 477 177 480 
rect 174 480 177 483 
rect 174 483 177 486 
rect 174 486 177 489 
rect 174 489 177 492 
rect 174 492 177 495 
rect 174 495 177 498 
rect 174 498 177 501 
rect 174 501 177 504 
rect 174 504 177 507 
rect 174 507 177 510 
rect 177 0 180 3 
rect 177 3 180 6 
rect 177 6 180 9 
rect 177 9 180 12 
rect 177 12 180 15 
rect 177 15 180 18 
rect 177 18 180 21 
rect 177 21 180 24 
rect 177 24 180 27 
rect 177 27 180 30 
rect 177 30 180 33 
rect 177 33 180 36 
rect 177 36 180 39 
rect 177 39 180 42 
rect 177 42 180 45 
rect 177 45 180 48 
rect 177 48 180 51 
rect 177 51 180 54 
rect 177 54 180 57 
rect 177 57 180 60 
rect 177 60 180 63 
rect 177 63 180 66 
rect 177 66 180 69 
rect 177 69 180 72 
rect 177 72 180 75 
rect 177 75 180 78 
rect 177 78 180 81 
rect 177 81 180 84 
rect 177 84 180 87 
rect 177 87 180 90 
rect 177 90 180 93 
rect 177 93 180 96 
rect 177 96 180 99 
rect 177 99 180 102 
rect 177 102 180 105 
rect 177 105 180 108 
rect 177 108 180 111 
rect 177 111 180 114 
rect 177 114 180 117 
rect 177 117 180 120 
rect 177 120 180 123 
rect 177 123 180 126 
rect 177 126 180 129 
rect 177 129 180 132 
rect 177 132 180 135 
rect 177 135 180 138 
rect 177 138 180 141 
rect 177 141 180 144 
rect 177 144 180 147 
rect 177 147 180 150 
rect 177 150 180 153 
rect 177 153 180 156 
rect 177 156 180 159 
rect 177 159 180 162 
rect 177 162 180 165 
rect 177 165 180 168 
rect 177 168 180 171 
rect 177 171 180 174 
rect 177 174 180 177 
rect 177 177 180 180 
rect 177 180 180 183 
rect 177 183 180 186 
rect 177 186 180 189 
rect 177 189 180 192 
rect 177 192 180 195 
rect 177 195 180 198 
rect 177 198 180 201 
rect 177 201 180 204 
rect 177 204 180 207 
rect 177 207 180 210 
rect 177 210 180 213 
rect 177 213 180 216 
rect 177 216 180 219 
rect 177 219 180 222 
rect 177 222 180 225 
rect 177 225 180 228 
rect 177 228 180 231 
rect 177 231 180 234 
rect 177 234 180 237 
rect 177 237 180 240 
rect 177 240 180 243 
rect 177 243 180 246 
rect 177 246 180 249 
rect 177 249 180 252 
rect 177 252 180 255 
rect 177 255 180 258 
rect 177 258 180 261 
rect 177 261 180 264 
rect 177 264 180 267 
rect 177 267 180 270 
rect 177 270 180 273 
rect 177 273 180 276 
rect 177 276 180 279 
rect 177 279 180 282 
rect 177 282 180 285 
rect 177 285 180 288 
rect 177 288 180 291 
rect 177 291 180 294 
rect 177 294 180 297 
rect 177 297 180 300 
rect 177 300 180 303 
rect 177 303 180 306 
rect 177 306 180 309 
rect 177 309 180 312 
rect 177 312 180 315 
rect 177 315 180 318 
rect 177 318 180 321 
rect 177 321 180 324 
rect 177 324 180 327 
rect 177 327 180 330 
rect 177 330 180 333 
rect 177 333 180 336 
rect 177 336 180 339 
rect 177 339 180 342 
rect 177 342 180 345 
rect 177 345 180 348 
rect 177 348 180 351 
rect 177 351 180 354 
rect 177 354 180 357 
rect 177 357 180 360 
rect 177 360 180 363 
rect 177 363 180 366 
rect 177 366 180 369 
rect 177 369 180 372 
rect 177 372 180 375 
rect 177 375 180 378 
rect 177 378 180 381 
rect 177 381 180 384 
rect 177 384 180 387 
rect 177 387 180 390 
rect 177 390 180 393 
rect 177 393 180 396 
rect 177 396 180 399 
rect 177 399 180 402 
rect 177 402 180 405 
rect 177 405 180 408 
rect 177 408 180 411 
rect 177 411 180 414 
rect 177 414 180 417 
rect 177 417 180 420 
rect 177 420 180 423 
rect 177 423 180 426 
rect 177 426 180 429 
rect 177 429 180 432 
rect 177 432 180 435 
rect 177 435 180 438 
rect 177 438 180 441 
rect 177 441 180 444 
rect 177 444 180 447 
rect 177 447 180 450 
rect 177 450 180 453 
rect 177 453 180 456 
rect 177 456 180 459 
rect 177 459 180 462 
rect 177 462 180 465 
rect 177 465 180 468 
rect 177 468 180 471 
rect 177 471 180 474 
rect 177 474 180 477 
rect 177 477 180 480 
rect 177 480 180 483 
rect 177 483 180 486 
rect 177 486 180 489 
rect 177 489 180 492 
rect 177 492 180 495 
rect 177 495 180 498 
rect 177 498 180 501 
rect 177 501 180 504 
rect 177 504 180 507 
rect 177 507 180 510 
rect 180 0 183 3 
rect 180 3 183 6 
rect 180 6 183 9 
rect 180 9 183 12 
rect 180 12 183 15 
rect 180 15 183 18 
rect 180 18 183 21 
rect 180 21 183 24 
rect 180 24 183 27 
rect 180 27 183 30 
rect 180 30 183 33 
rect 180 33 183 36 
rect 180 36 183 39 
rect 180 39 183 42 
rect 180 42 183 45 
rect 180 45 183 48 
rect 180 48 183 51 
rect 180 51 183 54 
rect 180 54 183 57 
rect 180 57 183 60 
rect 180 60 183 63 
rect 180 63 183 66 
rect 180 66 183 69 
rect 180 69 183 72 
rect 180 72 183 75 
rect 180 75 183 78 
rect 180 78 183 81 
rect 180 81 183 84 
rect 180 84 183 87 
rect 180 87 183 90 
rect 180 90 183 93 
rect 180 93 183 96 
rect 180 96 183 99 
rect 180 99 183 102 
rect 180 102 183 105 
rect 180 105 183 108 
rect 180 108 183 111 
rect 180 111 183 114 
rect 180 114 183 117 
rect 180 117 183 120 
rect 180 120 183 123 
rect 180 123 183 126 
rect 180 126 183 129 
rect 180 129 183 132 
rect 180 132 183 135 
rect 180 135 183 138 
rect 180 138 183 141 
rect 180 141 183 144 
rect 180 144 183 147 
rect 180 147 183 150 
rect 180 150 183 153 
rect 180 153 183 156 
rect 180 156 183 159 
rect 180 159 183 162 
rect 180 162 183 165 
rect 180 165 183 168 
rect 180 168 183 171 
rect 180 171 183 174 
rect 180 174 183 177 
rect 180 177 183 180 
rect 180 180 183 183 
rect 180 183 183 186 
rect 180 186 183 189 
rect 180 189 183 192 
rect 180 192 183 195 
rect 180 195 183 198 
rect 180 198 183 201 
rect 180 201 183 204 
rect 180 204 183 207 
rect 180 207 183 210 
rect 180 210 183 213 
rect 180 213 183 216 
rect 180 216 183 219 
rect 180 219 183 222 
rect 180 222 183 225 
rect 180 225 183 228 
rect 180 228 183 231 
rect 180 231 183 234 
rect 180 234 183 237 
rect 180 237 183 240 
rect 180 240 183 243 
rect 180 243 183 246 
rect 180 246 183 249 
rect 180 249 183 252 
rect 180 252 183 255 
rect 180 255 183 258 
rect 180 258 183 261 
rect 180 261 183 264 
rect 180 264 183 267 
rect 180 267 183 270 
rect 180 270 183 273 
rect 180 273 183 276 
rect 180 276 183 279 
rect 180 279 183 282 
rect 180 282 183 285 
rect 180 285 183 288 
rect 180 288 183 291 
rect 180 291 183 294 
rect 180 294 183 297 
rect 180 297 183 300 
rect 180 300 183 303 
rect 180 303 183 306 
rect 180 306 183 309 
rect 180 309 183 312 
rect 180 312 183 315 
rect 180 315 183 318 
rect 180 318 183 321 
rect 180 321 183 324 
rect 180 324 183 327 
rect 180 327 183 330 
rect 180 330 183 333 
rect 180 333 183 336 
rect 180 336 183 339 
rect 180 339 183 342 
rect 180 342 183 345 
rect 180 345 183 348 
rect 180 348 183 351 
rect 180 351 183 354 
rect 180 354 183 357 
rect 180 357 183 360 
rect 180 360 183 363 
rect 180 363 183 366 
rect 180 366 183 369 
rect 180 369 183 372 
rect 180 372 183 375 
rect 180 375 183 378 
rect 180 378 183 381 
rect 180 381 183 384 
rect 180 384 183 387 
rect 180 387 183 390 
rect 180 390 183 393 
rect 180 393 183 396 
rect 180 396 183 399 
rect 180 399 183 402 
rect 180 402 183 405 
rect 180 405 183 408 
rect 180 408 183 411 
rect 180 411 183 414 
rect 180 414 183 417 
rect 180 417 183 420 
rect 180 420 183 423 
rect 180 423 183 426 
rect 180 426 183 429 
rect 180 429 183 432 
rect 180 432 183 435 
rect 180 435 183 438 
rect 180 438 183 441 
rect 180 441 183 444 
rect 180 444 183 447 
rect 180 447 183 450 
rect 180 450 183 453 
rect 180 453 183 456 
rect 180 456 183 459 
rect 180 459 183 462 
rect 180 462 183 465 
rect 180 465 183 468 
rect 180 468 183 471 
rect 180 471 183 474 
rect 180 474 183 477 
rect 180 477 183 480 
rect 180 480 183 483 
rect 180 483 183 486 
rect 180 486 183 489 
rect 180 489 183 492 
rect 180 492 183 495 
rect 180 495 183 498 
rect 180 498 183 501 
rect 180 501 183 504 
rect 180 504 183 507 
rect 180 507 183 510 
rect 183 0 186 3 
rect 183 3 186 6 
rect 183 6 186 9 
rect 183 9 186 12 
rect 183 12 186 15 
rect 183 15 186 18 
rect 183 18 186 21 
rect 183 21 186 24 
rect 183 24 186 27 
rect 183 27 186 30 
rect 183 30 186 33 
rect 183 33 186 36 
rect 183 36 186 39 
rect 183 39 186 42 
rect 183 42 186 45 
rect 183 45 186 48 
rect 183 48 186 51 
rect 183 51 186 54 
rect 183 54 186 57 
rect 183 57 186 60 
rect 183 60 186 63 
rect 183 63 186 66 
rect 183 66 186 69 
rect 183 69 186 72 
rect 183 72 186 75 
rect 183 75 186 78 
rect 183 78 186 81 
rect 183 81 186 84 
rect 183 84 186 87 
rect 183 87 186 90 
rect 183 90 186 93 
rect 183 93 186 96 
rect 183 96 186 99 
rect 183 99 186 102 
rect 183 102 186 105 
rect 183 105 186 108 
rect 183 108 186 111 
rect 183 111 186 114 
rect 183 114 186 117 
rect 183 117 186 120 
rect 183 120 186 123 
rect 183 123 186 126 
rect 183 126 186 129 
rect 183 129 186 132 
rect 183 132 186 135 
rect 183 135 186 138 
rect 183 138 186 141 
rect 183 141 186 144 
rect 183 144 186 147 
rect 183 147 186 150 
rect 183 150 186 153 
rect 183 153 186 156 
rect 183 156 186 159 
rect 183 159 186 162 
rect 183 162 186 165 
rect 183 165 186 168 
rect 183 168 186 171 
rect 183 171 186 174 
rect 183 174 186 177 
rect 183 177 186 180 
rect 183 180 186 183 
rect 183 183 186 186 
rect 183 186 186 189 
rect 183 189 186 192 
rect 183 192 186 195 
rect 183 195 186 198 
rect 183 198 186 201 
rect 183 201 186 204 
rect 183 204 186 207 
rect 183 207 186 210 
rect 183 210 186 213 
rect 183 213 186 216 
rect 183 216 186 219 
rect 183 219 186 222 
rect 183 222 186 225 
rect 183 225 186 228 
rect 183 228 186 231 
rect 183 231 186 234 
rect 183 234 186 237 
rect 183 237 186 240 
rect 183 240 186 243 
rect 183 243 186 246 
rect 183 246 186 249 
rect 183 249 186 252 
rect 183 252 186 255 
rect 183 255 186 258 
rect 183 258 186 261 
rect 183 261 186 264 
rect 183 264 186 267 
rect 183 267 186 270 
rect 183 270 186 273 
rect 183 273 186 276 
rect 183 276 186 279 
rect 183 279 186 282 
rect 183 282 186 285 
rect 183 285 186 288 
rect 183 288 186 291 
rect 183 291 186 294 
rect 183 294 186 297 
rect 183 297 186 300 
rect 183 300 186 303 
rect 183 303 186 306 
rect 183 306 186 309 
rect 183 309 186 312 
rect 183 312 186 315 
rect 183 315 186 318 
rect 183 318 186 321 
rect 183 321 186 324 
rect 183 324 186 327 
rect 183 327 186 330 
rect 183 330 186 333 
rect 183 333 186 336 
rect 183 336 186 339 
rect 183 339 186 342 
rect 183 342 186 345 
rect 183 345 186 348 
rect 183 348 186 351 
rect 183 351 186 354 
rect 183 354 186 357 
rect 183 357 186 360 
rect 183 360 186 363 
rect 183 363 186 366 
rect 183 366 186 369 
rect 183 369 186 372 
rect 183 372 186 375 
rect 183 375 186 378 
rect 183 378 186 381 
rect 183 381 186 384 
rect 183 384 186 387 
rect 183 387 186 390 
rect 183 390 186 393 
rect 183 393 186 396 
rect 183 396 186 399 
rect 183 399 186 402 
rect 183 402 186 405 
rect 183 405 186 408 
rect 183 408 186 411 
rect 183 411 186 414 
rect 183 414 186 417 
rect 183 417 186 420 
rect 183 420 186 423 
rect 183 423 186 426 
rect 183 426 186 429 
rect 183 429 186 432 
rect 183 432 186 435 
rect 183 435 186 438 
rect 183 438 186 441 
rect 183 441 186 444 
rect 183 444 186 447 
rect 183 447 186 450 
rect 183 450 186 453 
rect 183 453 186 456 
rect 183 456 186 459 
rect 183 459 186 462 
rect 183 462 186 465 
rect 183 465 186 468 
rect 183 468 186 471 
rect 183 471 186 474 
rect 183 474 186 477 
rect 183 477 186 480 
rect 183 480 186 483 
rect 183 483 186 486 
rect 183 486 186 489 
rect 183 489 186 492 
rect 183 492 186 495 
rect 183 495 186 498 
rect 183 498 186 501 
rect 183 501 186 504 
rect 183 504 186 507 
rect 183 507 186 510 
rect 186 0 189 3 
rect 186 3 189 6 
rect 186 6 189 9 
rect 186 9 189 12 
rect 186 12 189 15 
rect 186 15 189 18 
rect 186 18 189 21 
rect 186 21 189 24 
rect 186 24 189 27 
rect 186 27 189 30 
rect 186 30 189 33 
rect 186 33 189 36 
rect 186 36 189 39 
rect 186 39 189 42 
rect 186 42 189 45 
rect 186 45 189 48 
rect 186 48 189 51 
rect 186 51 189 54 
rect 186 54 189 57 
rect 186 57 189 60 
rect 186 60 189 63 
rect 186 63 189 66 
rect 186 66 189 69 
rect 186 69 189 72 
rect 186 72 189 75 
rect 186 75 189 78 
rect 186 78 189 81 
rect 186 81 189 84 
rect 186 84 189 87 
rect 186 87 189 90 
rect 186 90 189 93 
rect 186 93 189 96 
rect 186 96 189 99 
rect 186 99 189 102 
rect 186 102 189 105 
rect 186 105 189 108 
rect 186 108 189 111 
rect 186 111 189 114 
rect 186 114 189 117 
rect 186 117 189 120 
rect 186 120 189 123 
rect 186 123 189 126 
rect 186 126 189 129 
rect 186 129 189 132 
rect 186 132 189 135 
rect 186 135 189 138 
rect 186 138 189 141 
rect 186 141 189 144 
rect 186 144 189 147 
rect 186 147 189 150 
rect 186 150 189 153 
rect 186 153 189 156 
rect 186 156 189 159 
rect 186 159 189 162 
rect 186 162 189 165 
rect 186 165 189 168 
rect 186 168 189 171 
rect 186 171 189 174 
rect 186 174 189 177 
rect 186 177 189 180 
rect 186 180 189 183 
rect 186 183 189 186 
rect 186 186 189 189 
rect 186 189 189 192 
rect 186 192 189 195 
rect 186 195 189 198 
rect 186 198 189 201 
rect 186 201 189 204 
rect 186 204 189 207 
rect 186 207 189 210 
rect 186 210 189 213 
rect 186 213 189 216 
rect 186 216 189 219 
rect 186 219 189 222 
rect 186 222 189 225 
rect 186 225 189 228 
rect 186 228 189 231 
rect 186 231 189 234 
rect 186 234 189 237 
rect 186 237 189 240 
rect 186 240 189 243 
rect 186 243 189 246 
rect 186 246 189 249 
rect 186 249 189 252 
rect 186 252 189 255 
rect 186 255 189 258 
rect 186 258 189 261 
rect 186 261 189 264 
rect 186 264 189 267 
rect 186 267 189 270 
rect 186 270 189 273 
rect 186 273 189 276 
rect 186 276 189 279 
rect 186 279 189 282 
rect 186 282 189 285 
rect 186 285 189 288 
rect 186 288 189 291 
rect 186 291 189 294 
rect 186 294 189 297 
rect 186 297 189 300 
rect 186 300 189 303 
rect 186 303 189 306 
rect 186 306 189 309 
rect 186 309 189 312 
rect 186 312 189 315 
rect 186 315 189 318 
rect 186 318 189 321 
rect 186 321 189 324 
rect 186 324 189 327 
rect 186 327 189 330 
rect 186 330 189 333 
rect 186 333 189 336 
rect 186 336 189 339 
rect 186 339 189 342 
rect 186 342 189 345 
rect 186 345 189 348 
rect 186 348 189 351 
rect 186 351 189 354 
rect 186 354 189 357 
rect 186 357 189 360 
rect 186 360 189 363 
rect 186 363 189 366 
rect 186 366 189 369 
rect 186 369 189 372 
rect 186 372 189 375 
rect 186 375 189 378 
rect 186 378 189 381 
rect 186 381 189 384 
rect 186 384 189 387 
rect 186 387 189 390 
rect 186 390 189 393 
rect 186 393 189 396 
rect 186 396 189 399 
rect 186 399 189 402 
rect 186 402 189 405 
rect 186 405 189 408 
rect 186 408 189 411 
rect 186 411 189 414 
rect 186 414 189 417 
rect 186 417 189 420 
rect 186 420 189 423 
rect 186 423 189 426 
rect 186 426 189 429 
rect 186 429 189 432 
rect 186 432 189 435 
rect 186 435 189 438 
rect 186 438 189 441 
rect 186 441 189 444 
rect 186 444 189 447 
rect 186 447 189 450 
rect 186 450 189 453 
rect 186 453 189 456 
rect 186 456 189 459 
rect 186 459 189 462 
rect 186 462 189 465 
rect 186 465 189 468 
rect 186 468 189 471 
rect 186 471 189 474 
rect 186 474 189 477 
rect 186 477 189 480 
rect 186 480 189 483 
rect 186 483 189 486 
rect 186 486 189 489 
rect 186 489 189 492 
rect 186 492 189 495 
rect 186 495 189 498 
rect 186 498 189 501 
rect 186 501 189 504 
rect 186 504 189 507 
rect 186 507 189 510 
rect 189 0 192 3 
rect 189 3 192 6 
rect 189 6 192 9 
rect 189 9 192 12 
rect 189 12 192 15 
rect 189 15 192 18 
rect 189 18 192 21 
rect 189 21 192 24 
rect 189 24 192 27 
rect 189 27 192 30 
rect 189 30 192 33 
rect 189 33 192 36 
rect 189 36 192 39 
rect 189 39 192 42 
rect 189 42 192 45 
rect 189 45 192 48 
rect 189 48 192 51 
rect 189 51 192 54 
rect 189 54 192 57 
rect 189 57 192 60 
rect 189 60 192 63 
rect 189 63 192 66 
rect 189 66 192 69 
rect 189 69 192 72 
rect 189 72 192 75 
rect 189 75 192 78 
rect 189 78 192 81 
rect 189 81 192 84 
rect 189 84 192 87 
rect 189 87 192 90 
rect 189 90 192 93 
rect 189 93 192 96 
rect 189 96 192 99 
rect 189 99 192 102 
rect 189 102 192 105 
rect 189 105 192 108 
rect 189 108 192 111 
rect 189 111 192 114 
rect 189 114 192 117 
rect 189 117 192 120 
rect 189 120 192 123 
rect 189 123 192 126 
rect 189 126 192 129 
rect 189 129 192 132 
rect 189 132 192 135 
rect 189 135 192 138 
rect 189 138 192 141 
rect 189 141 192 144 
rect 189 144 192 147 
rect 189 147 192 150 
rect 189 150 192 153 
rect 189 153 192 156 
rect 189 156 192 159 
rect 189 159 192 162 
rect 189 162 192 165 
rect 189 165 192 168 
rect 189 168 192 171 
rect 189 171 192 174 
rect 189 174 192 177 
rect 189 177 192 180 
rect 189 180 192 183 
rect 189 183 192 186 
rect 189 186 192 189 
rect 189 189 192 192 
rect 189 192 192 195 
rect 189 195 192 198 
rect 189 198 192 201 
rect 189 201 192 204 
rect 189 204 192 207 
rect 189 207 192 210 
rect 189 210 192 213 
rect 189 213 192 216 
rect 189 216 192 219 
rect 189 219 192 222 
rect 189 222 192 225 
rect 189 225 192 228 
rect 189 228 192 231 
rect 189 231 192 234 
rect 189 234 192 237 
rect 189 237 192 240 
rect 189 240 192 243 
rect 189 243 192 246 
rect 189 246 192 249 
rect 189 249 192 252 
rect 189 252 192 255 
rect 189 255 192 258 
rect 189 258 192 261 
rect 189 261 192 264 
rect 189 264 192 267 
rect 189 267 192 270 
rect 189 270 192 273 
rect 189 273 192 276 
rect 189 276 192 279 
rect 189 279 192 282 
rect 189 282 192 285 
rect 189 285 192 288 
rect 189 288 192 291 
rect 189 291 192 294 
rect 189 294 192 297 
rect 189 297 192 300 
rect 189 300 192 303 
rect 189 303 192 306 
rect 189 306 192 309 
rect 189 309 192 312 
rect 189 312 192 315 
rect 189 315 192 318 
rect 189 318 192 321 
rect 189 321 192 324 
rect 189 324 192 327 
rect 189 327 192 330 
rect 189 330 192 333 
rect 189 333 192 336 
rect 189 336 192 339 
rect 189 339 192 342 
rect 189 342 192 345 
rect 189 345 192 348 
rect 189 348 192 351 
rect 189 351 192 354 
rect 189 354 192 357 
rect 189 357 192 360 
rect 189 360 192 363 
rect 189 363 192 366 
rect 189 366 192 369 
rect 189 369 192 372 
rect 189 372 192 375 
rect 189 375 192 378 
rect 189 378 192 381 
rect 189 381 192 384 
rect 189 384 192 387 
rect 189 387 192 390 
rect 189 390 192 393 
rect 189 393 192 396 
rect 189 396 192 399 
rect 189 399 192 402 
rect 189 402 192 405 
rect 189 405 192 408 
rect 189 408 192 411 
rect 189 411 192 414 
rect 189 414 192 417 
rect 189 417 192 420 
rect 189 420 192 423 
rect 189 423 192 426 
rect 189 426 192 429 
rect 189 429 192 432 
rect 189 432 192 435 
rect 189 435 192 438 
rect 189 438 192 441 
rect 189 441 192 444 
rect 189 444 192 447 
rect 189 447 192 450 
rect 189 450 192 453 
rect 189 453 192 456 
rect 189 456 192 459 
rect 189 459 192 462 
rect 189 462 192 465 
rect 189 465 192 468 
rect 189 468 192 471 
rect 189 471 192 474 
rect 189 474 192 477 
rect 189 477 192 480 
rect 189 480 192 483 
rect 189 483 192 486 
rect 189 486 192 489 
rect 189 489 192 492 
rect 189 492 192 495 
rect 189 495 192 498 
rect 189 498 192 501 
rect 189 501 192 504 
rect 189 504 192 507 
rect 189 507 192 510 
rect 192 0 195 3 
rect 192 3 195 6 
rect 192 6 195 9 
rect 192 9 195 12 
rect 192 12 195 15 
rect 192 15 195 18 
rect 192 18 195 21 
rect 192 21 195 24 
rect 192 24 195 27 
rect 192 27 195 30 
rect 192 30 195 33 
rect 192 33 195 36 
rect 192 36 195 39 
rect 192 39 195 42 
rect 192 42 195 45 
rect 192 45 195 48 
rect 192 48 195 51 
rect 192 51 195 54 
rect 192 54 195 57 
rect 192 57 195 60 
rect 192 60 195 63 
rect 192 63 195 66 
rect 192 66 195 69 
rect 192 69 195 72 
rect 192 72 195 75 
rect 192 75 195 78 
rect 192 78 195 81 
rect 192 81 195 84 
rect 192 84 195 87 
rect 192 87 195 90 
rect 192 90 195 93 
rect 192 93 195 96 
rect 192 96 195 99 
rect 192 99 195 102 
rect 192 102 195 105 
rect 192 105 195 108 
rect 192 108 195 111 
rect 192 111 195 114 
rect 192 114 195 117 
rect 192 117 195 120 
rect 192 120 195 123 
rect 192 123 195 126 
rect 192 126 195 129 
rect 192 129 195 132 
rect 192 132 195 135 
rect 192 135 195 138 
rect 192 138 195 141 
rect 192 141 195 144 
rect 192 144 195 147 
rect 192 147 195 150 
rect 192 150 195 153 
rect 192 153 195 156 
rect 192 156 195 159 
rect 192 159 195 162 
rect 192 162 195 165 
rect 192 165 195 168 
rect 192 168 195 171 
rect 192 171 195 174 
rect 192 174 195 177 
rect 192 177 195 180 
rect 192 180 195 183 
rect 192 183 195 186 
rect 192 186 195 189 
rect 192 189 195 192 
rect 192 192 195 195 
rect 192 195 195 198 
rect 192 198 195 201 
rect 192 201 195 204 
rect 192 204 195 207 
rect 192 207 195 210 
rect 192 210 195 213 
rect 192 213 195 216 
rect 192 216 195 219 
rect 192 219 195 222 
rect 192 222 195 225 
rect 192 225 195 228 
rect 192 228 195 231 
rect 192 231 195 234 
rect 192 234 195 237 
rect 192 237 195 240 
rect 192 240 195 243 
rect 192 243 195 246 
rect 192 246 195 249 
rect 192 249 195 252 
rect 192 252 195 255 
rect 192 255 195 258 
rect 192 258 195 261 
rect 192 261 195 264 
rect 192 264 195 267 
rect 192 267 195 270 
rect 192 270 195 273 
rect 192 273 195 276 
rect 192 276 195 279 
rect 192 279 195 282 
rect 192 282 195 285 
rect 192 285 195 288 
rect 192 288 195 291 
rect 192 291 195 294 
rect 192 294 195 297 
rect 192 297 195 300 
rect 192 300 195 303 
rect 192 303 195 306 
rect 192 306 195 309 
rect 192 309 195 312 
rect 192 312 195 315 
rect 192 315 195 318 
rect 192 318 195 321 
rect 192 321 195 324 
rect 192 324 195 327 
rect 192 327 195 330 
rect 192 330 195 333 
rect 192 333 195 336 
rect 192 336 195 339 
rect 192 339 195 342 
rect 192 342 195 345 
rect 192 345 195 348 
rect 192 348 195 351 
rect 192 351 195 354 
rect 192 354 195 357 
rect 192 357 195 360 
rect 192 360 195 363 
rect 192 363 195 366 
rect 192 366 195 369 
rect 192 369 195 372 
rect 192 372 195 375 
rect 192 375 195 378 
rect 192 378 195 381 
rect 192 381 195 384 
rect 192 384 195 387 
rect 192 387 195 390 
rect 192 390 195 393 
rect 192 393 195 396 
rect 192 396 195 399 
rect 192 399 195 402 
rect 192 402 195 405 
rect 192 405 195 408 
rect 192 408 195 411 
rect 192 411 195 414 
rect 192 414 195 417 
rect 192 417 195 420 
rect 192 420 195 423 
rect 192 423 195 426 
rect 192 426 195 429 
rect 192 429 195 432 
rect 192 432 195 435 
rect 192 435 195 438 
rect 192 438 195 441 
rect 192 441 195 444 
rect 192 444 195 447 
rect 192 447 195 450 
rect 192 450 195 453 
rect 192 453 195 456 
rect 192 456 195 459 
rect 192 459 195 462 
rect 192 462 195 465 
rect 192 465 195 468 
rect 192 468 195 471 
rect 192 471 195 474 
rect 192 474 195 477 
rect 192 477 195 480 
rect 192 480 195 483 
rect 192 483 195 486 
rect 192 486 195 489 
rect 192 489 195 492 
rect 192 492 195 495 
rect 192 495 195 498 
rect 192 498 195 501 
rect 192 501 195 504 
rect 192 504 195 507 
rect 192 507 195 510 
rect 195 0 198 3 
rect 195 3 198 6 
rect 195 6 198 9 
rect 195 9 198 12 
rect 195 12 198 15 
rect 195 15 198 18 
rect 195 18 198 21 
rect 195 21 198 24 
rect 195 24 198 27 
rect 195 27 198 30 
rect 195 30 198 33 
rect 195 33 198 36 
rect 195 36 198 39 
rect 195 39 198 42 
rect 195 42 198 45 
rect 195 45 198 48 
rect 195 48 198 51 
rect 195 51 198 54 
rect 195 54 198 57 
rect 195 57 198 60 
rect 195 60 198 63 
rect 195 63 198 66 
rect 195 66 198 69 
rect 195 69 198 72 
rect 195 72 198 75 
rect 195 75 198 78 
rect 195 78 198 81 
rect 195 81 198 84 
rect 195 84 198 87 
rect 195 87 198 90 
rect 195 90 198 93 
rect 195 93 198 96 
rect 195 96 198 99 
rect 195 99 198 102 
rect 195 102 198 105 
rect 195 105 198 108 
rect 195 108 198 111 
rect 195 111 198 114 
rect 195 114 198 117 
rect 195 117 198 120 
rect 195 120 198 123 
rect 195 123 198 126 
rect 195 126 198 129 
rect 195 129 198 132 
rect 195 132 198 135 
rect 195 135 198 138 
rect 195 138 198 141 
rect 195 141 198 144 
rect 195 144 198 147 
rect 195 147 198 150 
rect 195 150 198 153 
rect 195 153 198 156 
rect 195 156 198 159 
rect 195 159 198 162 
rect 195 162 198 165 
rect 195 165 198 168 
rect 195 168 198 171 
rect 195 171 198 174 
rect 195 174 198 177 
rect 195 177 198 180 
rect 195 180 198 183 
rect 195 183 198 186 
rect 195 186 198 189 
rect 195 189 198 192 
rect 195 192 198 195 
rect 195 195 198 198 
rect 195 198 198 201 
rect 195 201 198 204 
rect 195 204 198 207 
rect 195 207 198 210 
rect 195 210 198 213 
rect 195 213 198 216 
rect 195 216 198 219 
rect 195 219 198 222 
rect 195 222 198 225 
rect 195 225 198 228 
rect 195 228 198 231 
rect 195 231 198 234 
rect 195 234 198 237 
rect 195 237 198 240 
rect 195 240 198 243 
rect 195 243 198 246 
rect 195 246 198 249 
rect 195 249 198 252 
rect 195 252 198 255 
rect 195 255 198 258 
rect 195 258 198 261 
rect 195 261 198 264 
rect 195 264 198 267 
rect 195 267 198 270 
rect 195 270 198 273 
rect 195 273 198 276 
rect 195 276 198 279 
rect 195 279 198 282 
rect 195 282 198 285 
rect 195 285 198 288 
rect 195 288 198 291 
rect 195 291 198 294 
rect 195 294 198 297 
rect 195 297 198 300 
rect 195 300 198 303 
rect 195 303 198 306 
rect 195 306 198 309 
rect 195 309 198 312 
rect 195 312 198 315 
rect 195 315 198 318 
rect 195 318 198 321 
rect 195 321 198 324 
rect 195 324 198 327 
rect 195 327 198 330 
rect 195 330 198 333 
rect 195 333 198 336 
rect 195 336 198 339 
rect 195 339 198 342 
rect 195 342 198 345 
rect 195 345 198 348 
rect 195 348 198 351 
rect 195 351 198 354 
rect 195 354 198 357 
rect 195 357 198 360 
rect 195 360 198 363 
rect 195 363 198 366 
rect 195 366 198 369 
rect 195 369 198 372 
rect 195 372 198 375 
rect 195 375 198 378 
rect 195 378 198 381 
rect 195 381 198 384 
rect 195 384 198 387 
rect 195 387 198 390 
rect 195 390 198 393 
rect 195 393 198 396 
rect 195 396 198 399 
rect 195 399 198 402 
rect 195 402 198 405 
rect 195 405 198 408 
rect 195 408 198 411 
rect 195 411 198 414 
rect 195 414 198 417 
rect 195 417 198 420 
rect 195 420 198 423 
rect 195 423 198 426 
rect 195 426 198 429 
rect 195 429 198 432 
rect 195 432 198 435 
rect 195 435 198 438 
rect 195 438 198 441 
rect 195 441 198 444 
rect 195 444 198 447 
rect 195 447 198 450 
rect 195 450 198 453 
rect 195 453 198 456 
rect 195 456 198 459 
rect 195 459 198 462 
rect 195 462 198 465 
rect 195 465 198 468 
rect 195 468 198 471 
rect 195 471 198 474 
rect 195 474 198 477 
rect 195 477 198 480 
rect 195 480 198 483 
rect 195 483 198 486 
rect 195 486 198 489 
rect 195 489 198 492 
rect 195 492 198 495 
rect 195 495 198 498 
rect 195 498 198 501 
rect 195 501 198 504 
rect 195 504 198 507 
rect 195 507 198 510 
rect 198 0 201 3 
rect 198 3 201 6 
rect 198 6 201 9 
rect 198 9 201 12 
rect 198 12 201 15 
rect 198 15 201 18 
rect 198 18 201 21 
rect 198 21 201 24 
rect 198 24 201 27 
rect 198 27 201 30 
rect 198 30 201 33 
rect 198 33 201 36 
rect 198 36 201 39 
rect 198 39 201 42 
rect 198 42 201 45 
rect 198 45 201 48 
rect 198 48 201 51 
rect 198 51 201 54 
rect 198 54 201 57 
rect 198 57 201 60 
rect 198 60 201 63 
rect 198 63 201 66 
rect 198 66 201 69 
rect 198 69 201 72 
rect 198 72 201 75 
rect 198 75 201 78 
rect 198 78 201 81 
rect 198 81 201 84 
rect 198 84 201 87 
rect 198 87 201 90 
rect 198 90 201 93 
rect 198 93 201 96 
rect 198 96 201 99 
rect 198 99 201 102 
rect 198 102 201 105 
rect 198 105 201 108 
rect 198 108 201 111 
rect 198 111 201 114 
rect 198 114 201 117 
rect 198 117 201 120 
rect 198 120 201 123 
rect 198 123 201 126 
rect 198 126 201 129 
rect 198 129 201 132 
rect 198 132 201 135 
rect 198 135 201 138 
rect 198 138 201 141 
rect 198 141 201 144 
rect 198 144 201 147 
rect 198 147 201 150 
rect 198 150 201 153 
rect 198 153 201 156 
rect 198 156 201 159 
rect 198 159 201 162 
rect 198 162 201 165 
rect 198 165 201 168 
rect 198 168 201 171 
rect 198 171 201 174 
rect 198 174 201 177 
rect 198 177 201 180 
rect 198 180 201 183 
rect 198 183 201 186 
rect 198 186 201 189 
rect 198 189 201 192 
rect 198 192 201 195 
rect 198 195 201 198 
rect 198 198 201 201 
rect 198 201 201 204 
rect 198 204 201 207 
rect 198 207 201 210 
rect 198 210 201 213 
rect 198 213 201 216 
rect 198 216 201 219 
rect 198 219 201 222 
rect 198 222 201 225 
rect 198 225 201 228 
rect 198 228 201 231 
rect 198 231 201 234 
rect 198 234 201 237 
rect 198 237 201 240 
rect 198 240 201 243 
rect 198 243 201 246 
rect 198 246 201 249 
rect 198 249 201 252 
rect 198 252 201 255 
rect 198 255 201 258 
rect 198 258 201 261 
rect 198 261 201 264 
rect 198 264 201 267 
rect 198 267 201 270 
rect 198 270 201 273 
rect 198 273 201 276 
rect 198 276 201 279 
rect 198 279 201 282 
rect 198 282 201 285 
rect 198 285 201 288 
rect 198 288 201 291 
rect 198 291 201 294 
rect 198 294 201 297 
rect 198 297 201 300 
rect 198 300 201 303 
rect 198 303 201 306 
rect 198 306 201 309 
rect 198 309 201 312 
rect 198 312 201 315 
rect 198 315 201 318 
rect 198 318 201 321 
rect 198 321 201 324 
rect 198 324 201 327 
rect 198 327 201 330 
rect 198 330 201 333 
rect 198 333 201 336 
rect 198 336 201 339 
rect 198 339 201 342 
rect 198 342 201 345 
rect 198 345 201 348 
rect 198 348 201 351 
rect 198 351 201 354 
rect 198 354 201 357 
rect 198 357 201 360 
rect 198 360 201 363 
rect 198 363 201 366 
rect 198 366 201 369 
rect 198 369 201 372 
rect 198 372 201 375 
rect 198 375 201 378 
rect 198 378 201 381 
rect 198 381 201 384 
rect 198 384 201 387 
rect 198 387 201 390 
rect 198 390 201 393 
rect 198 393 201 396 
rect 198 396 201 399 
rect 198 399 201 402 
rect 198 402 201 405 
rect 198 405 201 408 
rect 198 408 201 411 
rect 198 411 201 414 
rect 198 414 201 417 
rect 198 417 201 420 
rect 198 420 201 423 
rect 198 423 201 426 
rect 198 426 201 429 
rect 198 429 201 432 
rect 198 432 201 435 
rect 198 435 201 438 
rect 198 438 201 441 
rect 198 441 201 444 
rect 198 444 201 447 
rect 198 447 201 450 
rect 198 450 201 453 
rect 198 453 201 456 
rect 198 456 201 459 
rect 198 459 201 462 
rect 198 462 201 465 
rect 198 465 201 468 
rect 198 468 201 471 
rect 198 471 201 474 
rect 198 474 201 477 
rect 198 477 201 480 
rect 198 480 201 483 
rect 198 483 201 486 
rect 198 486 201 489 
rect 198 489 201 492 
rect 198 492 201 495 
rect 198 495 201 498 
rect 198 498 201 501 
rect 198 501 201 504 
rect 198 504 201 507 
rect 198 507 201 510 
rect 201 0 204 3 
rect 201 3 204 6 
rect 201 6 204 9 
rect 201 9 204 12 
rect 201 12 204 15 
rect 201 15 204 18 
rect 201 18 204 21 
rect 201 21 204 24 
rect 201 24 204 27 
rect 201 27 204 30 
rect 201 30 204 33 
rect 201 33 204 36 
rect 201 36 204 39 
rect 201 39 204 42 
rect 201 42 204 45 
rect 201 45 204 48 
rect 201 48 204 51 
rect 201 51 204 54 
rect 201 54 204 57 
rect 201 57 204 60 
rect 201 60 204 63 
rect 201 63 204 66 
rect 201 66 204 69 
rect 201 69 204 72 
rect 201 72 204 75 
rect 201 75 204 78 
rect 201 78 204 81 
rect 201 81 204 84 
rect 201 84 204 87 
rect 201 87 204 90 
rect 201 90 204 93 
rect 201 93 204 96 
rect 201 96 204 99 
rect 201 99 204 102 
rect 201 102 204 105 
rect 201 105 204 108 
rect 201 108 204 111 
rect 201 111 204 114 
rect 201 114 204 117 
rect 201 117 204 120 
rect 201 120 204 123 
rect 201 123 204 126 
rect 201 126 204 129 
rect 201 129 204 132 
rect 201 132 204 135 
rect 201 135 204 138 
rect 201 138 204 141 
rect 201 141 204 144 
rect 201 144 204 147 
rect 201 147 204 150 
rect 201 150 204 153 
rect 201 153 204 156 
rect 201 156 204 159 
rect 201 159 204 162 
rect 201 162 204 165 
rect 201 165 204 168 
rect 201 168 204 171 
rect 201 171 204 174 
rect 201 174 204 177 
rect 201 177 204 180 
rect 201 180 204 183 
rect 201 183 204 186 
rect 201 186 204 189 
rect 201 189 204 192 
rect 201 192 204 195 
rect 201 195 204 198 
rect 201 198 204 201 
rect 201 201 204 204 
rect 201 204 204 207 
rect 201 207 204 210 
rect 201 210 204 213 
rect 201 213 204 216 
rect 201 216 204 219 
rect 201 219 204 222 
rect 201 222 204 225 
rect 201 225 204 228 
rect 201 228 204 231 
rect 201 231 204 234 
rect 201 234 204 237 
rect 201 237 204 240 
rect 201 240 204 243 
rect 201 243 204 246 
rect 201 246 204 249 
rect 201 249 204 252 
rect 201 252 204 255 
rect 201 255 204 258 
rect 201 258 204 261 
rect 201 261 204 264 
rect 201 264 204 267 
rect 201 267 204 270 
rect 201 270 204 273 
rect 201 273 204 276 
rect 201 276 204 279 
rect 201 279 204 282 
rect 201 282 204 285 
rect 201 285 204 288 
rect 201 288 204 291 
rect 201 291 204 294 
rect 201 294 204 297 
rect 201 297 204 300 
rect 201 300 204 303 
rect 201 303 204 306 
rect 201 306 204 309 
rect 201 309 204 312 
rect 201 312 204 315 
rect 201 315 204 318 
rect 201 318 204 321 
rect 201 321 204 324 
rect 201 324 204 327 
rect 201 327 204 330 
rect 201 330 204 333 
rect 201 333 204 336 
rect 201 336 204 339 
rect 201 339 204 342 
rect 201 342 204 345 
rect 201 345 204 348 
rect 201 348 204 351 
rect 201 351 204 354 
rect 201 354 204 357 
rect 201 357 204 360 
rect 201 360 204 363 
rect 201 363 204 366 
rect 201 366 204 369 
rect 201 369 204 372 
rect 201 372 204 375 
rect 201 375 204 378 
rect 201 378 204 381 
rect 201 381 204 384 
rect 201 384 204 387 
rect 201 387 204 390 
rect 201 390 204 393 
rect 201 393 204 396 
rect 201 396 204 399 
rect 201 399 204 402 
rect 201 402 204 405 
rect 201 405 204 408 
rect 201 408 204 411 
rect 201 411 204 414 
rect 201 414 204 417 
rect 201 417 204 420 
rect 201 420 204 423 
rect 201 423 204 426 
rect 201 426 204 429 
rect 201 429 204 432 
rect 201 432 204 435 
rect 201 435 204 438 
rect 201 438 204 441 
rect 201 441 204 444 
rect 201 444 204 447 
rect 201 447 204 450 
rect 201 450 204 453 
rect 201 453 204 456 
rect 201 456 204 459 
rect 201 459 204 462 
rect 201 462 204 465 
rect 201 465 204 468 
rect 201 468 204 471 
rect 201 471 204 474 
rect 201 474 204 477 
rect 201 477 204 480 
rect 201 480 204 483 
rect 201 483 204 486 
rect 201 486 204 489 
rect 201 489 204 492 
rect 201 492 204 495 
rect 201 495 204 498 
rect 201 498 204 501 
rect 201 501 204 504 
rect 201 504 204 507 
rect 201 507 204 510 
rect 204 0 207 3 
rect 204 3 207 6 
rect 204 6 207 9 
rect 204 9 207 12 
rect 204 12 207 15 
rect 204 15 207 18 
rect 204 18 207 21 
rect 204 21 207 24 
rect 204 24 207 27 
rect 204 27 207 30 
rect 204 30 207 33 
rect 204 33 207 36 
rect 204 36 207 39 
rect 204 39 207 42 
rect 204 42 207 45 
rect 204 45 207 48 
rect 204 48 207 51 
rect 204 51 207 54 
rect 204 54 207 57 
rect 204 57 207 60 
rect 204 60 207 63 
rect 204 63 207 66 
rect 204 66 207 69 
rect 204 69 207 72 
rect 204 72 207 75 
rect 204 75 207 78 
rect 204 78 207 81 
rect 204 81 207 84 
rect 204 84 207 87 
rect 204 87 207 90 
rect 204 90 207 93 
rect 204 93 207 96 
rect 204 96 207 99 
rect 204 99 207 102 
rect 204 102 207 105 
rect 204 105 207 108 
rect 204 108 207 111 
rect 204 111 207 114 
rect 204 114 207 117 
rect 204 117 207 120 
rect 204 120 207 123 
rect 204 123 207 126 
rect 204 126 207 129 
rect 204 129 207 132 
rect 204 132 207 135 
rect 204 135 207 138 
rect 204 138 207 141 
rect 204 141 207 144 
rect 204 144 207 147 
rect 204 147 207 150 
rect 204 150 207 153 
rect 204 153 207 156 
rect 204 156 207 159 
rect 204 159 207 162 
rect 204 162 207 165 
rect 204 165 207 168 
rect 204 168 207 171 
rect 204 171 207 174 
rect 204 174 207 177 
rect 204 177 207 180 
rect 204 180 207 183 
rect 204 183 207 186 
rect 204 186 207 189 
rect 204 189 207 192 
rect 204 192 207 195 
rect 204 195 207 198 
rect 204 198 207 201 
rect 204 201 207 204 
rect 204 204 207 207 
rect 204 207 207 210 
rect 204 210 207 213 
rect 204 213 207 216 
rect 204 216 207 219 
rect 204 219 207 222 
rect 204 222 207 225 
rect 204 225 207 228 
rect 204 228 207 231 
rect 204 231 207 234 
rect 204 234 207 237 
rect 204 237 207 240 
rect 204 240 207 243 
rect 204 243 207 246 
rect 204 246 207 249 
rect 204 249 207 252 
rect 204 252 207 255 
rect 204 255 207 258 
rect 204 258 207 261 
rect 204 261 207 264 
rect 204 264 207 267 
rect 204 267 207 270 
rect 204 270 207 273 
rect 204 273 207 276 
rect 204 276 207 279 
rect 204 279 207 282 
rect 204 282 207 285 
rect 204 285 207 288 
rect 204 288 207 291 
rect 204 291 207 294 
rect 204 294 207 297 
rect 204 297 207 300 
rect 204 300 207 303 
rect 204 303 207 306 
rect 204 306 207 309 
rect 204 309 207 312 
rect 204 312 207 315 
rect 204 315 207 318 
rect 204 318 207 321 
rect 204 321 207 324 
rect 204 324 207 327 
rect 204 327 207 330 
rect 204 330 207 333 
rect 204 333 207 336 
rect 204 336 207 339 
rect 204 339 207 342 
rect 204 342 207 345 
rect 204 345 207 348 
rect 204 348 207 351 
rect 204 351 207 354 
rect 204 354 207 357 
rect 204 357 207 360 
rect 204 360 207 363 
rect 204 363 207 366 
rect 204 366 207 369 
rect 204 369 207 372 
rect 204 372 207 375 
rect 204 375 207 378 
rect 204 378 207 381 
rect 204 381 207 384 
rect 204 384 207 387 
rect 204 387 207 390 
rect 204 390 207 393 
rect 204 393 207 396 
rect 204 396 207 399 
rect 204 399 207 402 
rect 204 402 207 405 
rect 204 405 207 408 
rect 204 408 207 411 
rect 204 411 207 414 
rect 204 414 207 417 
rect 204 417 207 420 
rect 204 420 207 423 
rect 204 423 207 426 
rect 204 426 207 429 
rect 204 429 207 432 
rect 204 432 207 435 
rect 204 435 207 438 
rect 204 438 207 441 
rect 204 441 207 444 
rect 204 444 207 447 
rect 204 447 207 450 
rect 204 450 207 453 
rect 204 453 207 456 
rect 204 456 207 459 
rect 204 459 207 462 
rect 204 462 207 465 
rect 204 465 207 468 
rect 204 468 207 471 
rect 204 471 207 474 
rect 204 474 207 477 
rect 204 477 207 480 
rect 204 480 207 483 
rect 204 483 207 486 
rect 204 486 207 489 
rect 204 489 207 492 
rect 204 492 207 495 
rect 204 495 207 498 
rect 204 498 207 501 
rect 204 501 207 504 
rect 204 504 207 507 
rect 204 507 207 510 
rect 207 0 210 3 
rect 207 3 210 6 
rect 207 6 210 9 
rect 207 9 210 12 
rect 207 12 210 15 
rect 207 15 210 18 
rect 207 18 210 21 
rect 207 21 210 24 
rect 207 24 210 27 
rect 207 27 210 30 
rect 207 30 210 33 
rect 207 33 210 36 
rect 207 36 210 39 
rect 207 39 210 42 
rect 207 42 210 45 
rect 207 45 210 48 
rect 207 48 210 51 
rect 207 51 210 54 
rect 207 54 210 57 
rect 207 57 210 60 
rect 207 60 210 63 
rect 207 63 210 66 
rect 207 66 210 69 
rect 207 69 210 72 
rect 207 72 210 75 
rect 207 75 210 78 
rect 207 78 210 81 
rect 207 81 210 84 
rect 207 84 210 87 
rect 207 87 210 90 
rect 207 90 210 93 
rect 207 93 210 96 
rect 207 96 210 99 
rect 207 99 210 102 
rect 207 102 210 105 
rect 207 105 210 108 
rect 207 108 210 111 
rect 207 111 210 114 
rect 207 114 210 117 
rect 207 117 210 120 
rect 207 120 210 123 
rect 207 123 210 126 
rect 207 126 210 129 
rect 207 129 210 132 
rect 207 132 210 135 
rect 207 135 210 138 
rect 207 138 210 141 
rect 207 141 210 144 
rect 207 144 210 147 
rect 207 147 210 150 
rect 207 150 210 153 
rect 207 153 210 156 
rect 207 156 210 159 
rect 207 159 210 162 
rect 207 162 210 165 
rect 207 165 210 168 
rect 207 168 210 171 
rect 207 171 210 174 
rect 207 174 210 177 
rect 207 177 210 180 
rect 207 180 210 183 
rect 207 183 210 186 
rect 207 186 210 189 
rect 207 189 210 192 
rect 207 192 210 195 
rect 207 195 210 198 
rect 207 198 210 201 
rect 207 201 210 204 
rect 207 204 210 207 
rect 207 207 210 210 
rect 207 210 210 213 
rect 207 213 210 216 
rect 207 216 210 219 
rect 207 219 210 222 
rect 207 222 210 225 
rect 207 225 210 228 
rect 207 228 210 231 
rect 207 231 210 234 
rect 207 234 210 237 
rect 207 237 210 240 
rect 207 240 210 243 
rect 207 243 210 246 
rect 207 246 210 249 
rect 207 249 210 252 
rect 207 252 210 255 
rect 207 255 210 258 
rect 207 258 210 261 
rect 207 261 210 264 
rect 207 264 210 267 
rect 207 267 210 270 
rect 207 270 210 273 
rect 207 273 210 276 
rect 207 276 210 279 
rect 207 279 210 282 
rect 207 282 210 285 
rect 207 285 210 288 
rect 207 288 210 291 
rect 207 291 210 294 
rect 207 294 210 297 
rect 207 297 210 300 
rect 207 300 210 303 
rect 207 303 210 306 
rect 207 306 210 309 
rect 207 309 210 312 
rect 207 312 210 315 
rect 207 315 210 318 
rect 207 318 210 321 
rect 207 321 210 324 
rect 207 324 210 327 
rect 207 327 210 330 
rect 207 330 210 333 
rect 207 333 210 336 
rect 207 336 210 339 
rect 207 339 210 342 
rect 207 342 210 345 
rect 207 345 210 348 
rect 207 348 210 351 
rect 207 351 210 354 
rect 207 354 210 357 
rect 207 357 210 360 
rect 207 360 210 363 
rect 207 363 210 366 
rect 207 366 210 369 
rect 207 369 210 372 
rect 207 372 210 375 
rect 207 375 210 378 
rect 207 378 210 381 
rect 207 381 210 384 
rect 207 384 210 387 
rect 207 387 210 390 
rect 207 390 210 393 
rect 207 393 210 396 
rect 207 396 210 399 
rect 207 399 210 402 
rect 207 402 210 405 
rect 207 405 210 408 
rect 207 408 210 411 
rect 207 411 210 414 
rect 207 414 210 417 
rect 207 417 210 420 
rect 207 420 210 423 
rect 207 423 210 426 
rect 207 426 210 429 
rect 207 429 210 432 
rect 207 432 210 435 
rect 207 435 210 438 
rect 207 438 210 441 
rect 207 441 210 444 
rect 207 444 210 447 
rect 207 447 210 450 
rect 207 450 210 453 
rect 207 453 210 456 
rect 207 456 210 459 
rect 207 459 210 462 
rect 207 462 210 465 
rect 207 465 210 468 
rect 207 468 210 471 
rect 207 471 210 474 
rect 207 474 210 477 
rect 207 477 210 480 
rect 207 480 210 483 
rect 207 483 210 486 
rect 207 486 210 489 
rect 207 489 210 492 
rect 207 492 210 495 
rect 207 495 210 498 
rect 207 498 210 501 
rect 207 501 210 504 
rect 207 504 210 507 
rect 207 507 210 510 
rect 210 0 213 3 
rect 210 3 213 6 
rect 210 6 213 9 
rect 210 9 213 12 
rect 210 12 213 15 
rect 210 15 213 18 
rect 210 18 213 21 
rect 210 21 213 24 
rect 210 24 213 27 
rect 210 27 213 30 
rect 210 30 213 33 
rect 210 33 213 36 
rect 210 36 213 39 
rect 210 39 213 42 
rect 210 42 213 45 
rect 210 45 213 48 
rect 210 48 213 51 
rect 210 51 213 54 
rect 210 54 213 57 
rect 210 57 213 60 
rect 210 60 213 63 
rect 210 63 213 66 
rect 210 66 213 69 
rect 210 69 213 72 
rect 210 72 213 75 
rect 210 75 213 78 
rect 210 78 213 81 
rect 210 81 213 84 
rect 210 84 213 87 
rect 210 87 213 90 
rect 210 90 213 93 
rect 210 93 213 96 
rect 210 96 213 99 
rect 210 99 213 102 
rect 210 102 213 105 
rect 210 105 213 108 
rect 210 108 213 111 
rect 210 111 213 114 
rect 210 114 213 117 
rect 210 117 213 120 
rect 210 120 213 123 
rect 210 123 213 126 
rect 210 126 213 129 
rect 210 129 213 132 
rect 210 132 213 135 
rect 210 135 213 138 
rect 210 138 213 141 
rect 210 141 213 144 
rect 210 144 213 147 
rect 210 147 213 150 
rect 210 150 213 153 
rect 210 153 213 156 
rect 210 156 213 159 
rect 210 159 213 162 
rect 210 162 213 165 
rect 210 165 213 168 
rect 210 168 213 171 
rect 210 171 213 174 
rect 210 174 213 177 
rect 210 177 213 180 
rect 210 180 213 183 
rect 210 183 213 186 
rect 210 186 213 189 
rect 210 189 213 192 
rect 210 192 213 195 
rect 210 195 213 198 
rect 210 198 213 201 
rect 210 201 213 204 
rect 210 204 213 207 
rect 210 207 213 210 
rect 210 210 213 213 
rect 210 213 213 216 
rect 210 216 213 219 
rect 210 219 213 222 
rect 210 222 213 225 
rect 210 225 213 228 
rect 210 228 213 231 
rect 210 231 213 234 
rect 210 234 213 237 
rect 210 237 213 240 
rect 210 240 213 243 
rect 210 243 213 246 
rect 210 246 213 249 
rect 210 249 213 252 
rect 210 252 213 255 
rect 210 255 213 258 
rect 210 258 213 261 
rect 210 261 213 264 
rect 210 264 213 267 
rect 210 267 213 270 
rect 210 270 213 273 
rect 210 273 213 276 
rect 210 276 213 279 
rect 210 279 213 282 
rect 210 282 213 285 
rect 210 285 213 288 
rect 210 288 213 291 
rect 210 291 213 294 
rect 210 294 213 297 
rect 210 297 213 300 
rect 210 300 213 303 
rect 210 303 213 306 
rect 210 306 213 309 
rect 210 309 213 312 
rect 210 312 213 315 
rect 210 315 213 318 
rect 210 318 213 321 
rect 210 321 213 324 
rect 210 324 213 327 
rect 210 327 213 330 
rect 210 330 213 333 
rect 210 333 213 336 
rect 210 336 213 339 
rect 210 339 213 342 
rect 210 342 213 345 
rect 210 345 213 348 
rect 210 348 213 351 
rect 210 351 213 354 
rect 210 354 213 357 
rect 210 357 213 360 
rect 210 360 213 363 
rect 210 363 213 366 
rect 210 366 213 369 
rect 210 369 213 372 
rect 210 372 213 375 
rect 210 375 213 378 
rect 210 378 213 381 
rect 210 381 213 384 
rect 210 384 213 387 
rect 210 387 213 390 
rect 210 390 213 393 
rect 210 393 213 396 
rect 210 396 213 399 
rect 210 399 213 402 
rect 210 402 213 405 
rect 210 405 213 408 
rect 210 408 213 411 
rect 210 411 213 414 
rect 210 414 213 417 
rect 210 417 213 420 
rect 210 420 213 423 
rect 210 423 213 426 
rect 210 426 213 429 
rect 210 429 213 432 
rect 210 432 213 435 
rect 210 435 213 438 
rect 210 438 213 441 
rect 210 441 213 444 
rect 210 444 213 447 
rect 210 447 213 450 
rect 210 450 213 453 
rect 210 453 213 456 
rect 210 456 213 459 
rect 210 459 213 462 
rect 210 462 213 465 
rect 210 465 213 468 
rect 210 468 213 471 
rect 210 471 213 474 
rect 210 474 213 477 
rect 210 477 213 480 
rect 210 480 213 483 
rect 210 483 213 486 
rect 210 486 213 489 
rect 210 489 213 492 
rect 210 492 213 495 
rect 210 495 213 498 
rect 210 498 213 501 
rect 210 501 213 504 
rect 210 504 213 507 
rect 210 507 213 510 
rect 213 0 216 3 
rect 213 3 216 6 
rect 213 6 216 9 
rect 213 9 216 12 
rect 213 12 216 15 
rect 213 15 216 18 
rect 213 18 216 21 
rect 213 21 216 24 
rect 213 24 216 27 
rect 213 27 216 30 
rect 213 30 216 33 
rect 213 33 216 36 
rect 213 36 216 39 
rect 213 39 216 42 
rect 213 42 216 45 
rect 213 45 216 48 
rect 213 48 216 51 
rect 213 51 216 54 
rect 213 54 216 57 
rect 213 57 216 60 
rect 213 60 216 63 
rect 213 63 216 66 
rect 213 66 216 69 
rect 213 69 216 72 
rect 213 72 216 75 
rect 213 75 216 78 
rect 213 78 216 81 
rect 213 81 216 84 
rect 213 84 216 87 
rect 213 87 216 90 
rect 213 90 216 93 
rect 213 93 216 96 
rect 213 96 216 99 
rect 213 99 216 102 
rect 213 102 216 105 
rect 213 105 216 108 
rect 213 108 216 111 
rect 213 111 216 114 
rect 213 114 216 117 
rect 213 117 216 120 
rect 213 120 216 123 
rect 213 123 216 126 
rect 213 126 216 129 
rect 213 129 216 132 
rect 213 132 216 135 
rect 213 135 216 138 
rect 213 138 216 141 
rect 213 141 216 144 
rect 213 144 216 147 
rect 213 147 216 150 
rect 213 150 216 153 
rect 213 153 216 156 
rect 213 156 216 159 
rect 213 159 216 162 
rect 213 162 216 165 
rect 213 165 216 168 
rect 213 168 216 171 
rect 213 171 216 174 
rect 213 174 216 177 
rect 213 177 216 180 
rect 213 180 216 183 
rect 213 183 216 186 
rect 213 186 216 189 
rect 213 189 216 192 
rect 213 192 216 195 
rect 213 195 216 198 
rect 213 198 216 201 
rect 213 201 216 204 
rect 213 204 216 207 
rect 213 207 216 210 
rect 213 210 216 213 
rect 213 213 216 216 
rect 213 216 216 219 
rect 213 219 216 222 
rect 213 222 216 225 
rect 213 225 216 228 
rect 213 228 216 231 
rect 213 231 216 234 
rect 213 234 216 237 
rect 213 237 216 240 
rect 213 240 216 243 
rect 213 243 216 246 
rect 213 246 216 249 
rect 213 249 216 252 
rect 213 252 216 255 
rect 213 255 216 258 
rect 213 258 216 261 
rect 213 261 216 264 
rect 213 264 216 267 
rect 213 267 216 270 
rect 213 270 216 273 
rect 213 273 216 276 
rect 213 276 216 279 
rect 213 279 216 282 
rect 213 282 216 285 
rect 213 285 216 288 
rect 213 288 216 291 
rect 213 291 216 294 
rect 213 294 216 297 
rect 213 297 216 300 
rect 213 300 216 303 
rect 213 303 216 306 
rect 213 306 216 309 
rect 213 309 216 312 
rect 213 312 216 315 
rect 213 315 216 318 
rect 213 318 216 321 
rect 213 321 216 324 
rect 213 324 216 327 
rect 213 327 216 330 
rect 213 330 216 333 
rect 213 333 216 336 
rect 213 336 216 339 
rect 213 339 216 342 
rect 213 342 216 345 
rect 213 345 216 348 
rect 213 348 216 351 
rect 213 351 216 354 
rect 213 354 216 357 
rect 213 357 216 360 
rect 213 360 216 363 
rect 213 363 216 366 
rect 213 366 216 369 
rect 213 369 216 372 
rect 213 372 216 375 
rect 213 375 216 378 
rect 213 378 216 381 
rect 213 381 216 384 
rect 213 384 216 387 
rect 213 387 216 390 
rect 213 390 216 393 
rect 213 393 216 396 
rect 213 396 216 399 
rect 213 399 216 402 
rect 213 402 216 405 
rect 213 405 216 408 
rect 213 408 216 411 
rect 213 411 216 414 
rect 213 414 216 417 
rect 213 417 216 420 
rect 213 420 216 423 
rect 213 423 216 426 
rect 213 426 216 429 
rect 213 429 216 432 
rect 213 432 216 435 
rect 213 435 216 438 
rect 213 438 216 441 
rect 213 441 216 444 
rect 213 444 216 447 
rect 213 447 216 450 
rect 213 450 216 453 
rect 213 453 216 456 
rect 213 456 216 459 
rect 213 459 216 462 
rect 213 462 216 465 
rect 213 465 216 468 
rect 213 468 216 471 
rect 213 471 216 474 
rect 213 474 216 477 
rect 213 477 216 480 
rect 213 480 216 483 
rect 213 483 216 486 
rect 213 486 216 489 
rect 213 489 216 492 
rect 213 492 216 495 
rect 213 495 216 498 
rect 213 498 216 501 
rect 213 501 216 504 
rect 213 504 216 507 
rect 213 507 216 510 
rect 216 0 219 3 
rect 216 3 219 6 
rect 216 6 219 9 
rect 216 9 219 12 
rect 216 12 219 15 
rect 216 15 219 18 
rect 216 18 219 21 
rect 216 21 219 24 
rect 216 24 219 27 
rect 216 27 219 30 
rect 216 30 219 33 
rect 216 33 219 36 
rect 216 36 219 39 
rect 216 39 219 42 
rect 216 42 219 45 
rect 216 45 219 48 
rect 216 48 219 51 
rect 216 51 219 54 
rect 216 54 219 57 
rect 216 57 219 60 
rect 216 60 219 63 
rect 216 63 219 66 
rect 216 66 219 69 
rect 216 69 219 72 
rect 216 72 219 75 
rect 216 75 219 78 
rect 216 78 219 81 
rect 216 81 219 84 
rect 216 84 219 87 
rect 216 87 219 90 
rect 216 90 219 93 
rect 216 93 219 96 
rect 216 96 219 99 
rect 216 99 219 102 
rect 216 102 219 105 
rect 216 105 219 108 
rect 216 108 219 111 
rect 216 111 219 114 
rect 216 114 219 117 
rect 216 117 219 120 
rect 216 120 219 123 
rect 216 123 219 126 
rect 216 126 219 129 
rect 216 129 219 132 
rect 216 132 219 135 
rect 216 135 219 138 
rect 216 138 219 141 
rect 216 141 219 144 
rect 216 144 219 147 
rect 216 147 219 150 
rect 216 150 219 153 
rect 216 153 219 156 
rect 216 156 219 159 
rect 216 159 219 162 
rect 216 162 219 165 
rect 216 165 219 168 
rect 216 168 219 171 
rect 216 171 219 174 
rect 216 174 219 177 
rect 216 177 219 180 
rect 216 180 219 183 
rect 216 183 219 186 
rect 216 186 219 189 
rect 216 189 219 192 
rect 216 192 219 195 
rect 216 195 219 198 
rect 216 198 219 201 
rect 216 201 219 204 
rect 216 204 219 207 
rect 216 207 219 210 
rect 216 210 219 213 
rect 216 213 219 216 
rect 216 216 219 219 
rect 216 219 219 222 
rect 216 222 219 225 
rect 216 225 219 228 
rect 216 228 219 231 
rect 216 231 219 234 
rect 216 234 219 237 
rect 216 237 219 240 
rect 216 240 219 243 
rect 216 243 219 246 
rect 216 246 219 249 
rect 216 249 219 252 
rect 216 252 219 255 
rect 216 255 219 258 
rect 216 258 219 261 
rect 216 261 219 264 
rect 216 264 219 267 
rect 216 267 219 270 
rect 216 270 219 273 
rect 216 273 219 276 
rect 216 276 219 279 
rect 216 279 219 282 
rect 216 282 219 285 
rect 216 285 219 288 
rect 216 288 219 291 
rect 216 291 219 294 
rect 216 294 219 297 
rect 216 297 219 300 
rect 216 300 219 303 
rect 216 303 219 306 
rect 216 306 219 309 
rect 216 309 219 312 
rect 216 312 219 315 
rect 216 315 219 318 
rect 216 318 219 321 
rect 216 321 219 324 
rect 216 324 219 327 
rect 216 327 219 330 
rect 216 330 219 333 
rect 216 333 219 336 
rect 216 336 219 339 
rect 216 339 219 342 
rect 216 342 219 345 
rect 216 345 219 348 
rect 216 348 219 351 
rect 216 351 219 354 
rect 216 354 219 357 
rect 216 357 219 360 
rect 216 360 219 363 
rect 216 363 219 366 
rect 216 366 219 369 
rect 216 369 219 372 
rect 216 372 219 375 
rect 216 375 219 378 
rect 216 378 219 381 
rect 216 381 219 384 
rect 216 384 219 387 
rect 216 387 219 390 
rect 216 390 219 393 
rect 216 393 219 396 
rect 216 396 219 399 
rect 216 399 219 402 
rect 216 402 219 405 
rect 216 405 219 408 
rect 216 408 219 411 
rect 216 411 219 414 
rect 216 414 219 417 
rect 216 417 219 420 
rect 216 420 219 423 
rect 216 423 219 426 
rect 216 426 219 429 
rect 216 429 219 432 
rect 216 432 219 435 
rect 216 435 219 438 
rect 216 438 219 441 
rect 216 441 219 444 
rect 216 444 219 447 
rect 216 447 219 450 
rect 216 450 219 453 
rect 216 453 219 456 
rect 216 456 219 459 
rect 216 459 219 462 
rect 216 462 219 465 
rect 216 465 219 468 
rect 216 468 219 471 
rect 216 471 219 474 
rect 216 474 219 477 
rect 216 477 219 480 
rect 216 480 219 483 
rect 216 483 219 486 
rect 216 486 219 489 
rect 216 489 219 492 
rect 216 492 219 495 
rect 216 495 219 498 
rect 216 498 219 501 
rect 216 501 219 504 
rect 216 504 219 507 
rect 216 507 219 510 
rect 219 0 222 3 
rect 219 3 222 6 
rect 219 6 222 9 
rect 219 9 222 12 
rect 219 12 222 15 
rect 219 15 222 18 
rect 219 18 222 21 
rect 219 21 222 24 
rect 219 24 222 27 
rect 219 27 222 30 
rect 219 30 222 33 
rect 219 33 222 36 
rect 219 36 222 39 
rect 219 39 222 42 
rect 219 42 222 45 
rect 219 45 222 48 
rect 219 48 222 51 
rect 219 51 222 54 
rect 219 54 222 57 
rect 219 57 222 60 
rect 219 60 222 63 
rect 219 63 222 66 
rect 219 66 222 69 
rect 219 69 222 72 
rect 219 72 222 75 
rect 219 75 222 78 
rect 219 78 222 81 
rect 219 81 222 84 
rect 219 84 222 87 
rect 219 87 222 90 
rect 219 90 222 93 
rect 219 93 222 96 
rect 219 96 222 99 
rect 219 99 222 102 
rect 219 102 222 105 
rect 219 105 222 108 
rect 219 108 222 111 
rect 219 111 222 114 
rect 219 114 222 117 
rect 219 117 222 120 
rect 219 120 222 123 
rect 219 123 222 126 
rect 219 126 222 129 
rect 219 129 222 132 
rect 219 132 222 135 
rect 219 135 222 138 
rect 219 138 222 141 
rect 219 141 222 144 
rect 219 144 222 147 
rect 219 147 222 150 
rect 219 150 222 153 
rect 219 153 222 156 
rect 219 156 222 159 
rect 219 159 222 162 
rect 219 162 222 165 
rect 219 165 222 168 
rect 219 168 222 171 
rect 219 171 222 174 
rect 219 174 222 177 
rect 219 177 222 180 
rect 219 180 222 183 
rect 219 183 222 186 
rect 219 186 222 189 
rect 219 189 222 192 
rect 219 192 222 195 
rect 219 195 222 198 
rect 219 198 222 201 
rect 219 201 222 204 
rect 219 204 222 207 
rect 219 207 222 210 
rect 219 210 222 213 
rect 219 213 222 216 
rect 219 216 222 219 
rect 219 219 222 222 
rect 219 222 222 225 
rect 219 225 222 228 
rect 219 228 222 231 
rect 219 231 222 234 
rect 219 234 222 237 
rect 219 237 222 240 
rect 219 240 222 243 
rect 219 243 222 246 
rect 219 246 222 249 
rect 219 249 222 252 
rect 219 252 222 255 
rect 219 255 222 258 
rect 219 258 222 261 
rect 219 261 222 264 
rect 219 264 222 267 
rect 219 267 222 270 
rect 219 270 222 273 
rect 219 273 222 276 
rect 219 276 222 279 
rect 219 279 222 282 
rect 219 282 222 285 
rect 219 285 222 288 
rect 219 288 222 291 
rect 219 291 222 294 
rect 219 294 222 297 
rect 219 297 222 300 
rect 219 300 222 303 
rect 219 303 222 306 
rect 219 306 222 309 
rect 219 309 222 312 
rect 219 312 222 315 
rect 219 315 222 318 
rect 219 318 222 321 
rect 219 321 222 324 
rect 219 324 222 327 
rect 219 327 222 330 
rect 219 330 222 333 
rect 219 333 222 336 
rect 219 336 222 339 
rect 219 339 222 342 
rect 219 342 222 345 
rect 219 345 222 348 
rect 219 348 222 351 
rect 219 351 222 354 
rect 219 354 222 357 
rect 219 357 222 360 
rect 219 360 222 363 
rect 219 363 222 366 
rect 219 366 222 369 
rect 219 369 222 372 
rect 219 372 222 375 
rect 219 375 222 378 
rect 219 378 222 381 
rect 219 381 222 384 
rect 219 384 222 387 
rect 219 387 222 390 
rect 219 390 222 393 
rect 219 393 222 396 
rect 219 396 222 399 
rect 219 399 222 402 
rect 219 402 222 405 
rect 219 405 222 408 
rect 219 408 222 411 
rect 219 411 222 414 
rect 219 414 222 417 
rect 219 417 222 420 
rect 219 420 222 423 
rect 219 423 222 426 
rect 219 426 222 429 
rect 219 429 222 432 
rect 219 432 222 435 
rect 219 435 222 438 
rect 219 438 222 441 
rect 219 441 222 444 
rect 219 444 222 447 
rect 219 447 222 450 
rect 219 450 222 453 
rect 219 453 222 456 
rect 219 456 222 459 
rect 219 459 222 462 
rect 219 462 222 465 
rect 219 465 222 468 
rect 219 468 222 471 
rect 219 471 222 474 
rect 219 474 222 477 
rect 219 477 222 480 
rect 219 480 222 483 
rect 219 483 222 486 
rect 219 486 222 489 
rect 219 489 222 492 
rect 219 492 222 495 
rect 219 495 222 498 
rect 219 498 222 501 
rect 219 501 222 504 
rect 219 504 222 507 
rect 219 507 222 510 
rect 222 0 225 3 
rect 222 3 225 6 
rect 222 6 225 9 
rect 222 9 225 12 
rect 222 12 225 15 
rect 222 15 225 18 
rect 222 18 225 21 
rect 222 21 225 24 
rect 222 24 225 27 
rect 222 27 225 30 
rect 222 30 225 33 
rect 222 33 225 36 
rect 222 36 225 39 
rect 222 39 225 42 
rect 222 42 225 45 
rect 222 45 225 48 
rect 222 48 225 51 
rect 222 51 225 54 
rect 222 54 225 57 
rect 222 57 225 60 
rect 222 60 225 63 
rect 222 63 225 66 
rect 222 66 225 69 
rect 222 69 225 72 
rect 222 72 225 75 
rect 222 75 225 78 
rect 222 78 225 81 
rect 222 81 225 84 
rect 222 84 225 87 
rect 222 87 225 90 
rect 222 90 225 93 
rect 222 93 225 96 
rect 222 96 225 99 
rect 222 99 225 102 
rect 222 102 225 105 
rect 222 105 225 108 
rect 222 108 225 111 
rect 222 111 225 114 
rect 222 114 225 117 
rect 222 117 225 120 
rect 222 120 225 123 
rect 222 123 225 126 
rect 222 126 225 129 
rect 222 129 225 132 
rect 222 132 225 135 
rect 222 135 225 138 
rect 222 138 225 141 
rect 222 141 225 144 
rect 222 144 225 147 
rect 222 147 225 150 
rect 222 150 225 153 
rect 222 153 225 156 
rect 222 156 225 159 
rect 222 159 225 162 
rect 222 162 225 165 
rect 222 165 225 168 
rect 222 168 225 171 
rect 222 171 225 174 
rect 222 174 225 177 
rect 222 177 225 180 
rect 222 180 225 183 
rect 222 183 225 186 
rect 222 186 225 189 
rect 222 189 225 192 
rect 222 192 225 195 
rect 222 195 225 198 
rect 222 198 225 201 
rect 222 201 225 204 
rect 222 204 225 207 
rect 222 207 225 210 
rect 222 210 225 213 
rect 222 213 225 216 
rect 222 216 225 219 
rect 222 219 225 222 
rect 222 222 225 225 
rect 222 225 225 228 
rect 222 228 225 231 
rect 222 231 225 234 
rect 222 234 225 237 
rect 222 237 225 240 
rect 222 240 225 243 
rect 222 243 225 246 
rect 222 246 225 249 
rect 222 249 225 252 
rect 222 252 225 255 
rect 222 255 225 258 
rect 222 258 225 261 
rect 222 261 225 264 
rect 222 264 225 267 
rect 222 267 225 270 
rect 222 270 225 273 
rect 222 273 225 276 
rect 222 276 225 279 
rect 222 279 225 282 
rect 222 282 225 285 
rect 222 285 225 288 
rect 222 288 225 291 
rect 222 291 225 294 
rect 222 294 225 297 
rect 222 297 225 300 
rect 222 300 225 303 
rect 222 303 225 306 
rect 222 306 225 309 
rect 222 309 225 312 
rect 222 312 225 315 
rect 222 315 225 318 
rect 222 318 225 321 
rect 222 321 225 324 
rect 222 324 225 327 
rect 222 327 225 330 
rect 222 330 225 333 
rect 222 333 225 336 
rect 222 336 225 339 
rect 222 339 225 342 
rect 222 342 225 345 
rect 222 345 225 348 
rect 222 348 225 351 
rect 222 351 225 354 
rect 222 354 225 357 
rect 222 357 225 360 
rect 222 360 225 363 
rect 222 363 225 366 
rect 222 366 225 369 
rect 222 369 225 372 
rect 222 372 225 375 
rect 222 375 225 378 
rect 222 378 225 381 
rect 222 381 225 384 
rect 222 384 225 387 
rect 222 387 225 390 
rect 222 390 225 393 
rect 222 393 225 396 
rect 222 396 225 399 
rect 222 399 225 402 
rect 222 402 225 405 
rect 222 405 225 408 
rect 222 408 225 411 
rect 222 411 225 414 
rect 222 414 225 417 
rect 222 417 225 420 
rect 222 420 225 423 
rect 222 423 225 426 
rect 222 426 225 429 
rect 222 429 225 432 
rect 222 432 225 435 
rect 222 435 225 438 
rect 222 438 225 441 
rect 222 441 225 444 
rect 222 444 225 447 
rect 222 447 225 450 
rect 222 450 225 453 
rect 222 453 225 456 
rect 222 456 225 459 
rect 222 459 225 462 
rect 222 462 225 465 
rect 222 465 225 468 
rect 222 468 225 471 
rect 222 471 225 474 
rect 222 474 225 477 
rect 222 477 225 480 
rect 222 480 225 483 
rect 222 483 225 486 
rect 222 486 225 489 
rect 222 489 225 492 
rect 222 492 225 495 
rect 222 495 225 498 
rect 222 498 225 501 
rect 222 501 225 504 
rect 222 504 225 507 
rect 222 507 225 510 
rect 225 0 228 3 
rect 225 3 228 6 
rect 225 6 228 9 
rect 225 9 228 12 
rect 225 12 228 15 
rect 225 15 228 18 
rect 225 18 228 21 
rect 225 21 228 24 
rect 225 24 228 27 
rect 225 27 228 30 
rect 225 30 228 33 
rect 225 33 228 36 
rect 225 36 228 39 
rect 225 39 228 42 
rect 225 42 228 45 
rect 225 45 228 48 
rect 225 48 228 51 
rect 225 51 228 54 
rect 225 54 228 57 
rect 225 57 228 60 
rect 225 60 228 63 
rect 225 63 228 66 
rect 225 66 228 69 
rect 225 69 228 72 
rect 225 72 228 75 
rect 225 75 228 78 
rect 225 78 228 81 
rect 225 81 228 84 
rect 225 84 228 87 
rect 225 87 228 90 
rect 225 90 228 93 
rect 225 93 228 96 
rect 225 96 228 99 
rect 225 99 228 102 
rect 225 102 228 105 
rect 225 105 228 108 
rect 225 108 228 111 
rect 225 111 228 114 
rect 225 114 228 117 
rect 225 117 228 120 
rect 225 120 228 123 
rect 225 123 228 126 
rect 225 126 228 129 
rect 225 129 228 132 
rect 225 132 228 135 
rect 225 135 228 138 
rect 225 138 228 141 
rect 225 141 228 144 
rect 225 144 228 147 
rect 225 147 228 150 
rect 225 150 228 153 
rect 225 153 228 156 
rect 225 156 228 159 
rect 225 159 228 162 
rect 225 162 228 165 
rect 225 165 228 168 
rect 225 168 228 171 
rect 225 171 228 174 
rect 225 174 228 177 
rect 225 177 228 180 
rect 225 180 228 183 
rect 225 183 228 186 
rect 225 186 228 189 
rect 225 189 228 192 
rect 225 192 228 195 
rect 225 195 228 198 
rect 225 198 228 201 
rect 225 201 228 204 
rect 225 204 228 207 
rect 225 207 228 210 
rect 225 210 228 213 
rect 225 213 228 216 
rect 225 216 228 219 
rect 225 219 228 222 
rect 225 222 228 225 
rect 225 225 228 228 
rect 225 228 228 231 
rect 225 231 228 234 
rect 225 234 228 237 
rect 225 237 228 240 
rect 225 240 228 243 
rect 225 243 228 246 
rect 225 246 228 249 
rect 225 249 228 252 
rect 225 252 228 255 
rect 225 255 228 258 
rect 225 258 228 261 
rect 225 261 228 264 
rect 225 264 228 267 
rect 225 267 228 270 
rect 225 270 228 273 
rect 225 273 228 276 
rect 225 276 228 279 
rect 225 279 228 282 
rect 225 282 228 285 
rect 225 285 228 288 
rect 225 288 228 291 
rect 225 291 228 294 
rect 225 294 228 297 
rect 225 297 228 300 
rect 225 300 228 303 
rect 225 303 228 306 
rect 225 306 228 309 
rect 225 309 228 312 
rect 225 312 228 315 
rect 225 315 228 318 
rect 225 318 228 321 
rect 225 321 228 324 
rect 225 324 228 327 
rect 225 327 228 330 
rect 225 330 228 333 
rect 225 333 228 336 
rect 225 336 228 339 
rect 225 339 228 342 
rect 225 342 228 345 
rect 225 345 228 348 
rect 225 348 228 351 
rect 225 351 228 354 
rect 225 354 228 357 
rect 225 357 228 360 
rect 225 360 228 363 
rect 225 363 228 366 
rect 225 366 228 369 
rect 225 369 228 372 
rect 225 372 228 375 
rect 225 375 228 378 
rect 225 378 228 381 
rect 225 381 228 384 
rect 225 384 228 387 
rect 225 387 228 390 
rect 225 390 228 393 
rect 225 393 228 396 
rect 225 396 228 399 
rect 225 399 228 402 
rect 225 402 228 405 
rect 225 405 228 408 
rect 225 408 228 411 
rect 225 411 228 414 
rect 225 414 228 417 
rect 225 417 228 420 
rect 225 420 228 423 
rect 225 423 228 426 
rect 225 426 228 429 
rect 225 429 228 432 
rect 225 432 228 435 
rect 225 435 228 438 
rect 225 438 228 441 
rect 225 441 228 444 
rect 225 444 228 447 
rect 225 447 228 450 
rect 225 450 228 453 
rect 225 453 228 456 
rect 225 456 228 459 
rect 225 459 228 462 
rect 225 462 228 465 
rect 225 465 228 468 
rect 225 468 228 471 
rect 225 471 228 474 
rect 225 474 228 477 
rect 225 477 228 480 
rect 225 480 228 483 
rect 225 483 228 486 
rect 225 486 228 489 
rect 225 489 228 492 
rect 225 492 228 495 
rect 225 495 228 498 
rect 225 498 228 501 
rect 225 501 228 504 
rect 225 504 228 507 
rect 225 507 228 510 
rect 228 0 231 3 
rect 228 3 231 6 
rect 228 6 231 9 
rect 228 9 231 12 
rect 228 12 231 15 
rect 228 15 231 18 
rect 228 18 231 21 
rect 228 21 231 24 
rect 228 24 231 27 
rect 228 27 231 30 
rect 228 30 231 33 
rect 228 33 231 36 
rect 228 36 231 39 
rect 228 39 231 42 
rect 228 42 231 45 
rect 228 45 231 48 
rect 228 48 231 51 
rect 228 51 231 54 
rect 228 54 231 57 
rect 228 57 231 60 
rect 228 60 231 63 
rect 228 63 231 66 
rect 228 66 231 69 
rect 228 69 231 72 
rect 228 72 231 75 
rect 228 75 231 78 
rect 228 78 231 81 
rect 228 81 231 84 
rect 228 84 231 87 
rect 228 87 231 90 
rect 228 90 231 93 
rect 228 93 231 96 
rect 228 96 231 99 
rect 228 99 231 102 
rect 228 102 231 105 
rect 228 105 231 108 
rect 228 108 231 111 
rect 228 111 231 114 
rect 228 114 231 117 
rect 228 117 231 120 
rect 228 120 231 123 
rect 228 123 231 126 
rect 228 126 231 129 
rect 228 129 231 132 
rect 228 132 231 135 
rect 228 135 231 138 
rect 228 138 231 141 
rect 228 141 231 144 
rect 228 144 231 147 
rect 228 147 231 150 
rect 228 150 231 153 
rect 228 153 231 156 
rect 228 156 231 159 
rect 228 159 231 162 
rect 228 162 231 165 
rect 228 165 231 168 
rect 228 168 231 171 
rect 228 171 231 174 
rect 228 174 231 177 
rect 228 177 231 180 
rect 228 180 231 183 
rect 228 183 231 186 
rect 228 186 231 189 
rect 228 189 231 192 
rect 228 192 231 195 
rect 228 195 231 198 
rect 228 198 231 201 
rect 228 201 231 204 
rect 228 204 231 207 
rect 228 207 231 210 
rect 228 210 231 213 
rect 228 213 231 216 
rect 228 216 231 219 
rect 228 219 231 222 
rect 228 222 231 225 
rect 228 225 231 228 
rect 228 228 231 231 
rect 228 231 231 234 
rect 228 234 231 237 
rect 228 237 231 240 
rect 228 240 231 243 
rect 228 243 231 246 
rect 228 246 231 249 
rect 228 249 231 252 
rect 228 252 231 255 
rect 228 255 231 258 
rect 228 258 231 261 
rect 228 261 231 264 
rect 228 264 231 267 
rect 228 267 231 270 
rect 228 270 231 273 
rect 228 273 231 276 
rect 228 276 231 279 
rect 228 279 231 282 
rect 228 282 231 285 
rect 228 285 231 288 
rect 228 288 231 291 
rect 228 291 231 294 
rect 228 294 231 297 
rect 228 297 231 300 
rect 228 300 231 303 
rect 228 303 231 306 
rect 228 306 231 309 
rect 228 309 231 312 
rect 228 312 231 315 
rect 228 315 231 318 
rect 228 318 231 321 
rect 228 321 231 324 
rect 228 324 231 327 
rect 228 327 231 330 
rect 228 330 231 333 
rect 228 333 231 336 
rect 228 336 231 339 
rect 228 339 231 342 
rect 228 342 231 345 
rect 228 345 231 348 
rect 228 348 231 351 
rect 228 351 231 354 
rect 228 354 231 357 
rect 228 357 231 360 
rect 228 360 231 363 
rect 228 363 231 366 
rect 228 366 231 369 
rect 228 369 231 372 
rect 228 372 231 375 
rect 228 375 231 378 
rect 228 378 231 381 
rect 228 381 231 384 
rect 228 384 231 387 
rect 228 387 231 390 
rect 228 390 231 393 
rect 228 393 231 396 
rect 228 396 231 399 
rect 228 399 231 402 
rect 228 402 231 405 
rect 228 405 231 408 
rect 228 408 231 411 
rect 228 411 231 414 
rect 228 414 231 417 
rect 228 417 231 420 
rect 228 420 231 423 
rect 228 423 231 426 
rect 228 426 231 429 
rect 228 429 231 432 
rect 228 432 231 435 
rect 228 435 231 438 
rect 228 438 231 441 
rect 228 441 231 444 
rect 228 444 231 447 
rect 228 447 231 450 
rect 228 450 231 453 
rect 228 453 231 456 
rect 228 456 231 459 
rect 228 459 231 462 
rect 228 462 231 465 
rect 228 465 231 468 
rect 228 468 231 471 
rect 228 471 231 474 
rect 228 474 231 477 
rect 228 477 231 480 
rect 228 480 231 483 
rect 228 483 231 486 
rect 228 486 231 489 
rect 228 489 231 492 
rect 228 492 231 495 
rect 228 495 231 498 
rect 228 498 231 501 
rect 228 501 231 504 
rect 228 504 231 507 
rect 228 507 231 510 
rect 231 0 234 3 
rect 231 3 234 6 
rect 231 6 234 9 
rect 231 9 234 12 
rect 231 12 234 15 
rect 231 15 234 18 
rect 231 18 234 21 
rect 231 21 234 24 
rect 231 24 234 27 
rect 231 27 234 30 
rect 231 30 234 33 
rect 231 33 234 36 
rect 231 36 234 39 
rect 231 39 234 42 
rect 231 42 234 45 
rect 231 45 234 48 
rect 231 48 234 51 
rect 231 51 234 54 
rect 231 54 234 57 
rect 231 57 234 60 
rect 231 60 234 63 
rect 231 63 234 66 
rect 231 66 234 69 
rect 231 69 234 72 
rect 231 72 234 75 
rect 231 75 234 78 
rect 231 78 234 81 
rect 231 81 234 84 
rect 231 84 234 87 
rect 231 87 234 90 
rect 231 90 234 93 
rect 231 93 234 96 
rect 231 96 234 99 
rect 231 99 234 102 
rect 231 102 234 105 
rect 231 105 234 108 
rect 231 108 234 111 
rect 231 111 234 114 
rect 231 114 234 117 
rect 231 117 234 120 
rect 231 120 234 123 
rect 231 123 234 126 
rect 231 126 234 129 
rect 231 129 234 132 
rect 231 132 234 135 
rect 231 135 234 138 
rect 231 138 234 141 
rect 231 141 234 144 
rect 231 144 234 147 
rect 231 147 234 150 
rect 231 150 234 153 
rect 231 153 234 156 
rect 231 156 234 159 
rect 231 159 234 162 
rect 231 162 234 165 
rect 231 165 234 168 
rect 231 168 234 171 
rect 231 171 234 174 
rect 231 174 234 177 
rect 231 177 234 180 
rect 231 180 234 183 
rect 231 183 234 186 
rect 231 186 234 189 
rect 231 189 234 192 
rect 231 192 234 195 
rect 231 195 234 198 
rect 231 198 234 201 
rect 231 201 234 204 
rect 231 204 234 207 
rect 231 207 234 210 
rect 231 210 234 213 
rect 231 213 234 216 
rect 231 216 234 219 
rect 231 219 234 222 
rect 231 222 234 225 
rect 231 225 234 228 
rect 231 228 234 231 
rect 231 231 234 234 
rect 231 234 234 237 
rect 231 237 234 240 
rect 231 240 234 243 
rect 231 243 234 246 
rect 231 246 234 249 
rect 231 249 234 252 
rect 231 252 234 255 
rect 231 255 234 258 
rect 231 258 234 261 
rect 231 261 234 264 
rect 231 264 234 267 
rect 231 267 234 270 
rect 231 270 234 273 
rect 231 273 234 276 
rect 231 276 234 279 
rect 231 279 234 282 
rect 231 282 234 285 
rect 231 285 234 288 
rect 231 288 234 291 
rect 231 291 234 294 
rect 231 294 234 297 
rect 231 297 234 300 
rect 231 300 234 303 
rect 231 303 234 306 
rect 231 306 234 309 
rect 231 309 234 312 
rect 231 312 234 315 
rect 231 315 234 318 
rect 231 318 234 321 
rect 231 321 234 324 
rect 231 324 234 327 
rect 231 327 234 330 
rect 231 330 234 333 
rect 231 333 234 336 
rect 231 336 234 339 
rect 231 339 234 342 
rect 231 342 234 345 
rect 231 345 234 348 
rect 231 348 234 351 
rect 231 351 234 354 
rect 231 354 234 357 
rect 231 357 234 360 
rect 231 360 234 363 
rect 231 363 234 366 
rect 231 366 234 369 
rect 231 369 234 372 
rect 231 372 234 375 
rect 231 375 234 378 
rect 231 378 234 381 
rect 231 381 234 384 
rect 231 384 234 387 
rect 231 387 234 390 
rect 231 390 234 393 
rect 231 393 234 396 
rect 231 396 234 399 
rect 231 399 234 402 
rect 231 402 234 405 
rect 231 405 234 408 
rect 231 408 234 411 
rect 231 411 234 414 
rect 231 414 234 417 
rect 231 417 234 420 
rect 231 420 234 423 
rect 231 423 234 426 
rect 231 426 234 429 
rect 231 429 234 432 
rect 231 432 234 435 
rect 231 435 234 438 
rect 231 438 234 441 
rect 231 441 234 444 
rect 231 444 234 447 
rect 231 447 234 450 
rect 231 450 234 453 
rect 231 453 234 456 
rect 231 456 234 459 
rect 231 459 234 462 
rect 231 462 234 465 
rect 231 465 234 468 
rect 231 468 234 471 
rect 231 471 234 474 
rect 231 474 234 477 
rect 231 477 234 480 
rect 231 480 234 483 
rect 231 483 234 486 
rect 231 486 234 489 
rect 231 489 234 492 
rect 231 492 234 495 
rect 231 495 234 498 
rect 231 498 234 501 
rect 231 501 234 504 
rect 231 504 234 507 
rect 231 507 234 510 
rect 234 0 237 3 
rect 234 3 237 6 
rect 234 6 237 9 
rect 234 9 237 12 
rect 234 12 237 15 
rect 234 15 237 18 
rect 234 18 237 21 
rect 234 21 237 24 
rect 234 24 237 27 
rect 234 27 237 30 
rect 234 30 237 33 
rect 234 33 237 36 
rect 234 36 237 39 
rect 234 39 237 42 
rect 234 42 237 45 
rect 234 45 237 48 
rect 234 48 237 51 
rect 234 51 237 54 
rect 234 54 237 57 
rect 234 57 237 60 
rect 234 60 237 63 
rect 234 63 237 66 
rect 234 66 237 69 
rect 234 69 237 72 
rect 234 72 237 75 
rect 234 75 237 78 
rect 234 78 237 81 
rect 234 81 237 84 
rect 234 84 237 87 
rect 234 87 237 90 
rect 234 90 237 93 
rect 234 93 237 96 
rect 234 96 237 99 
rect 234 99 237 102 
rect 234 102 237 105 
rect 234 105 237 108 
rect 234 108 237 111 
rect 234 111 237 114 
rect 234 114 237 117 
rect 234 117 237 120 
rect 234 120 237 123 
rect 234 123 237 126 
rect 234 126 237 129 
rect 234 129 237 132 
rect 234 132 237 135 
rect 234 135 237 138 
rect 234 138 237 141 
rect 234 141 237 144 
rect 234 144 237 147 
rect 234 147 237 150 
rect 234 150 237 153 
rect 234 153 237 156 
rect 234 156 237 159 
rect 234 159 237 162 
rect 234 162 237 165 
rect 234 165 237 168 
rect 234 168 237 171 
rect 234 171 237 174 
rect 234 174 237 177 
rect 234 177 237 180 
rect 234 180 237 183 
rect 234 183 237 186 
rect 234 186 237 189 
rect 234 189 237 192 
rect 234 192 237 195 
rect 234 195 237 198 
rect 234 198 237 201 
rect 234 201 237 204 
rect 234 204 237 207 
rect 234 207 237 210 
rect 234 210 237 213 
rect 234 213 237 216 
rect 234 216 237 219 
rect 234 219 237 222 
rect 234 222 237 225 
rect 234 225 237 228 
rect 234 228 237 231 
rect 234 231 237 234 
rect 234 234 237 237 
rect 234 237 237 240 
rect 234 240 237 243 
rect 234 243 237 246 
rect 234 246 237 249 
rect 234 249 237 252 
rect 234 252 237 255 
rect 234 255 237 258 
rect 234 258 237 261 
rect 234 261 237 264 
rect 234 264 237 267 
rect 234 267 237 270 
rect 234 270 237 273 
rect 234 273 237 276 
rect 234 276 237 279 
rect 234 279 237 282 
rect 234 282 237 285 
rect 234 285 237 288 
rect 234 288 237 291 
rect 234 291 237 294 
rect 234 294 237 297 
rect 234 297 237 300 
rect 234 300 237 303 
rect 234 303 237 306 
rect 234 306 237 309 
rect 234 309 237 312 
rect 234 312 237 315 
rect 234 315 237 318 
rect 234 318 237 321 
rect 234 321 237 324 
rect 234 324 237 327 
rect 234 327 237 330 
rect 234 330 237 333 
rect 234 333 237 336 
rect 234 336 237 339 
rect 234 339 237 342 
rect 234 342 237 345 
rect 234 345 237 348 
rect 234 348 237 351 
rect 234 351 237 354 
rect 234 354 237 357 
rect 234 357 237 360 
rect 234 360 237 363 
rect 234 363 237 366 
rect 234 366 237 369 
rect 234 369 237 372 
rect 234 372 237 375 
rect 234 375 237 378 
rect 234 378 237 381 
rect 234 381 237 384 
rect 234 384 237 387 
rect 234 387 237 390 
rect 234 390 237 393 
rect 234 393 237 396 
rect 234 396 237 399 
rect 234 399 237 402 
rect 234 402 237 405 
rect 234 405 237 408 
rect 234 408 237 411 
rect 234 411 237 414 
rect 234 414 237 417 
rect 234 417 237 420 
rect 234 420 237 423 
rect 234 423 237 426 
rect 234 426 237 429 
rect 234 429 237 432 
rect 234 432 237 435 
rect 234 435 237 438 
rect 234 438 237 441 
rect 234 441 237 444 
rect 234 444 237 447 
rect 234 447 237 450 
rect 234 450 237 453 
rect 234 453 237 456 
rect 234 456 237 459 
rect 234 459 237 462 
rect 234 462 237 465 
rect 234 465 237 468 
rect 234 468 237 471 
rect 234 471 237 474 
rect 234 474 237 477 
rect 234 477 237 480 
rect 234 480 237 483 
rect 234 483 237 486 
rect 234 486 237 489 
rect 234 489 237 492 
rect 234 492 237 495 
rect 234 495 237 498 
rect 234 498 237 501 
rect 234 501 237 504 
rect 234 504 237 507 
rect 234 507 237 510 
rect 237 0 240 3 
rect 237 3 240 6 
rect 237 6 240 9 
rect 237 9 240 12 
rect 237 12 240 15 
rect 237 15 240 18 
rect 237 18 240 21 
rect 237 21 240 24 
rect 237 24 240 27 
rect 237 27 240 30 
rect 237 30 240 33 
rect 237 33 240 36 
rect 237 36 240 39 
rect 237 39 240 42 
rect 237 42 240 45 
rect 237 45 240 48 
rect 237 48 240 51 
rect 237 51 240 54 
rect 237 54 240 57 
rect 237 57 240 60 
rect 237 60 240 63 
rect 237 63 240 66 
rect 237 66 240 69 
rect 237 69 240 72 
rect 237 72 240 75 
rect 237 75 240 78 
rect 237 78 240 81 
rect 237 81 240 84 
rect 237 84 240 87 
rect 237 87 240 90 
rect 237 90 240 93 
rect 237 93 240 96 
rect 237 96 240 99 
rect 237 99 240 102 
rect 237 102 240 105 
rect 237 105 240 108 
rect 237 108 240 111 
rect 237 111 240 114 
rect 237 114 240 117 
rect 237 117 240 120 
rect 237 120 240 123 
rect 237 123 240 126 
rect 237 126 240 129 
rect 237 129 240 132 
rect 237 132 240 135 
rect 237 135 240 138 
rect 237 138 240 141 
rect 237 141 240 144 
rect 237 144 240 147 
rect 237 147 240 150 
rect 237 150 240 153 
rect 237 153 240 156 
rect 237 156 240 159 
rect 237 159 240 162 
rect 237 162 240 165 
rect 237 165 240 168 
rect 237 168 240 171 
rect 237 171 240 174 
rect 237 174 240 177 
rect 237 177 240 180 
rect 237 180 240 183 
rect 237 183 240 186 
rect 237 186 240 189 
rect 237 189 240 192 
rect 237 192 240 195 
rect 237 195 240 198 
rect 237 198 240 201 
rect 237 201 240 204 
rect 237 204 240 207 
rect 237 207 240 210 
rect 237 210 240 213 
rect 237 213 240 216 
rect 237 216 240 219 
rect 237 219 240 222 
rect 237 222 240 225 
rect 237 225 240 228 
rect 237 228 240 231 
rect 237 231 240 234 
rect 237 234 240 237 
rect 237 237 240 240 
rect 237 240 240 243 
rect 237 243 240 246 
rect 237 246 240 249 
rect 237 249 240 252 
rect 237 252 240 255 
rect 237 255 240 258 
rect 237 258 240 261 
rect 237 261 240 264 
rect 237 264 240 267 
rect 237 267 240 270 
rect 237 270 240 273 
rect 237 273 240 276 
rect 237 276 240 279 
rect 237 279 240 282 
rect 237 282 240 285 
rect 237 285 240 288 
rect 237 288 240 291 
rect 237 291 240 294 
rect 237 294 240 297 
rect 237 297 240 300 
rect 237 300 240 303 
rect 237 303 240 306 
rect 237 306 240 309 
rect 237 309 240 312 
rect 237 312 240 315 
rect 237 315 240 318 
rect 237 318 240 321 
rect 237 321 240 324 
rect 237 324 240 327 
rect 237 327 240 330 
rect 237 330 240 333 
rect 237 333 240 336 
rect 237 336 240 339 
rect 237 339 240 342 
rect 237 342 240 345 
rect 237 345 240 348 
rect 237 348 240 351 
rect 237 351 240 354 
rect 237 354 240 357 
rect 237 357 240 360 
rect 237 360 240 363 
rect 237 363 240 366 
rect 237 366 240 369 
rect 237 369 240 372 
rect 237 372 240 375 
rect 237 375 240 378 
rect 237 378 240 381 
rect 237 381 240 384 
rect 237 384 240 387 
rect 237 387 240 390 
rect 237 390 240 393 
rect 237 393 240 396 
rect 237 396 240 399 
rect 237 399 240 402 
rect 237 402 240 405 
rect 237 405 240 408 
rect 237 408 240 411 
rect 237 411 240 414 
rect 237 414 240 417 
rect 237 417 240 420 
rect 237 420 240 423 
rect 237 423 240 426 
rect 237 426 240 429 
rect 237 429 240 432 
rect 237 432 240 435 
rect 237 435 240 438 
rect 237 438 240 441 
rect 237 441 240 444 
rect 237 444 240 447 
rect 237 447 240 450 
rect 237 450 240 453 
rect 237 453 240 456 
rect 237 456 240 459 
rect 237 459 240 462 
rect 237 462 240 465 
rect 237 465 240 468 
rect 237 468 240 471 
rect 237 471 240 474 
rect 237 474 240 477 
rect 237 477 240 480 
rect 237 480 240 483 
rect 237 483 240 486 
rect 237 486 240 489 
rect 237 489 240 492 
rect 237 492 240 495 
rect 237 495 240 498 
rect 237 498 240 501 
rect 237 501 240 504 
rect 237 504 240 507 
rect 237 507 240 510 
rect 240 0 243 3 
rect 240 3 243 6 
rect 240 6 243 9 
rect 240 9 243 12 
rect 240 12 243 15 
rect 240 15 243 18 
rect 240 18 243 21 
rect 240 21 243 24 
rect 240 24 243 27 
rect 240 27 243 30 
rect 240 30 243 33 
rect 240 33 243 36 
rect 240 36 243 39 
rect 240 39 243 42 
rect 240 42 243 45 
rect 240 45 243 48 
rect 240 48 243 51 
rect 240 51 243 54 
rect 240 54 243 57 
rect 240 57 243 60 
rect 240 60 243 63 
rect 240 63 243 66 
rect 240 66 243 69 
rect 240 69 243 72 
rect 240 72 243 75 
rect 240 75 243 78 
rect 240 78 243 81 
rect 240 81 243 84 
rect 240 84 243 87 
rect 240 87 243 90 
rect 240 90 243 93 
rect 240 93 243 96 
rect 240 96 243 99 
rect 240 99 243 102 
rect 240 102 243 105 
rect 240 105 243 108 
rect 240 108 243 111 
rect 240 111 243 114 
rect 240 114 243 117 
rect 240 117 243 120 
rect 240 120 243 123 
rect 240 123 243 126 
rect 240 126 243 129 
rect 240 129 243 132 
rect 240 132 243 135 
rect 240 135 243 138 
rect 240 138 243 141 
rect 240 141 243 144 
rect 240 144 243 147 
rect 240 147 243 150 
rect 240 150 243 153 
rect 240 153 243 156 
rect 240 156 243 159 
rect 240 159 243 162 
rect 240 162 243 165 
rect 240 165 243 168 
rect 240 168 243 171 
rect 240 171 243 174 
rect 240 174 243 177 
rect 240 177 243 180 
rect 240 180 243 183 
rect 240 183 243 186 
rect 240 186 243 189 
rect 240 189 243 192 
rect 240 192 243 195 
rect 240 195 243 198 
rect 240 198 243 201 
rect 240 201 243 204 
rect 240 204 243 207 
rect 240 207 243 210 
rect 240 210 243 213 
rect 240 213 243 216 
rect 240 216 243 219 
rect 240 219 243 222 
rect 240 222 243 225 
rect 240 225 243 228 
rect 240 228 243 231 
rect 240 231 243 234 
rect 240 234 243 237 
rect 240 237 243 240 
rect 240 240 243 243 
rect 240 243 243 246 
rect 240 246 243 249 
rect 240 249 243 252 
rect 240 252 243 255 
rect 240 255 243 258 
rect 240 258 243 261 
rect 240 261 243 264 
rect 240 264 243 267 
rect 240 267 243 270 
rect 240 270 243 273 
rect 240 273 243 276 
rect 240 276 243 279 
rect 240 279 243 282 
rect 240 282 243 285 
rect 240 285 243 288 
rect 240 288 243 291 
rect 240 291 243 294 
rect 240 294 243 297 
rect 240 297 243 300 
rect 240 300 243 303 
rect 240 303 243 306 
rect 240 306 243 309 
rect 240 309 243 312 
rect 240 312 243 315 
rect 240 315 243 318 
rect 240 318 243 321 
rect 240 321 243 324 
rect 240 324 243 327 
rect 240 327 243 330 
rect 240 330 243 333 
rect 240 333 243 336 
rect 240 336 243 339 
rect 240 339 243 342 
rect 240 342 243 345 
rect 240 345 243 348 
rect 240 348 243 351 
rect 240 351 243 354 
rect 240 354 243 357 
rect 240 357 243 360 
rect 240 360 243 363 
rect 240 363 243 366 
rect 240 366 243 369 
rect 240 369 243 372 
rect 240 372 243 375 
rect 240 375 243 378 
rect 240 378 243 381 
rect 240 381 243 384 
rect 240 384 243 387 
rect 240 387 243 390 
rect 240 390 243 393 
rect 240 393 243 396 
rect 240 396 243 399 
rect 240 399 243 402 
rect 240 402 243 405 
rect 240 405 243 408 
rect 240 408 243 411 
rect 240 411 243 414 
rect 240 414 243 417 
rect 240 417 243 420 
rect 240 420 243 423 
rect 240 423 243 426 
rect 240 426 243 429 
rect 240 429 243 432 
rect 240 432 243 435 
rect 240 435 243 438 
rect 240 438 243 441 
rect 240 441 243 444 
rect 240 444 243 447 
rect 240 447 243 450 
rect 240 450 243 453 
rect 240 453 243 456 
rect 240 456 243 459 
rect 240 459 243 462 
rect 240 462 243 465 
rect 240 465 243 468 
rect 240 468 243 471 
rect 240 471 243 474 
rect 240 474 243 477 
rect 240 477 243 480 
rect 240 480 243 483 
rect 240 483 243 486 
rect 240 486 243 489 
rect 240 489 243 492 
rect 240 492 243 495 
rect 240 495 243 498 
rect 240 498 243 501 
rect 240 501 243 504 
rect 240 504 243 507 
rect 240 507 243 510 
rect 243 0 246 3 
rect 243 3 246 6 
rect 243 6 246 9 
rect 243 9 246 12 
rect 243 12 246 15 
rect 243 15 246 18 
rect 243 18 246 21 
rect 243 21 246 24 
rect 243 24 246 27 
rect 243 27 246 30 
rect 243 30 246 33 
rect 243 33 246 36 
rect 243 36 246 39 
rect 243 39 246 42 
rect 243 42 246 45 
rect 243 45 246 48 
rect 243 48 246 51 
rect 243 51 246 54 
rect 243 54 246 57 
rect 243 57 246 60 
rect 243 60 246 63 
rect 243 63 246 66 
rect 243 66 246 69 
rect 243 69 246 72 
rect 243 72 246 75 
rect 243 75 246 78 
rect 243 78 246 81 
rect 243 81 246 84 
rect 243 84 246 87 
rect 243 87 246 90 
rect 243 90 246 93 
rect 243 93 246 96 
rect 243 96 246 99 
rect 243 99 246 102 
rect 243 102 246 105 
rect 243 105 246 108 
rect 243 108 246 111 
rect 243 111 246 114 
rect 243 114 246 117 
rect 243 117 246 120 
rect 243 120 246 123 
rect 243 123 246 126 
rect 243 126 246 129 
rect 243 129 246 132 
rect 243 132 246 135 
rect 243 135 246 138 
rect 243 138 246 141 
rect 243 141 246 144 
rect 243 144 246 147 
rect 243 147 246 150 
rect 243 150 246 153 
rect 243 153 246 156 
rect 243 156 246 159 
rect 243 159 246 162 
rect 243 162 246 165 
rect 243 165 246 168 
rect 243 168 246 171 
rect 243 171 246 174 
rect 243 174 246 177 
rect 243 177 246 180 
rect 243 180 246 183 
rect 243 183 246 186 
rect 243 186 246 189 
rect 243 189 246 192 
rect 243 192 246 195 
rect 243 195 246 198 
rect 243 198 246 201 
rect 243 201 246 204 
rect 243 204 246 207 
rect 243 207 246 210 
rect 243 210 246 213 
rect 243 213 246 216 
rect 243 216 246 219 
rect 243 219 246 222 
rect 243 222 246 225 
rect 243 225 246 228 
rect 243 228 246 231 
rect 243 231 246 234 
rect 243 234 246 237 
rect 243 237 246 240 
rect 243 240 246 243 
rect 243 243 246 246 
rect 243 246 246 249 
rect 243 249 246 252 
rect 243 252 246 255 
rect 243 255 246 258 
rect 243 258 246 261 
rect 243 261 246 264 
rect 243 264 246 267 
rect 243 267 246 270 
rect 243 270 246 273 
rect 243 273 246 276 
rect 243 276 246 279 
rect 243 279 246 282 
rect 243 282 246 285 
rect 243 285 246 288 
rect 243 288 246 291 
rect 243 291 246 294 
rect 243 294 246 297 
rect 243 297 246 300 
rect 243 300 246 303 
rect 243 303 246 306 
rect 243 306 246 309 
rect 243 309 246 312 
rect 243 312 246 315 
rect 243 315 246 318 
rect 243 318 246 321 
rect 243 321 246 324 
rect 243 324 246 327 
rect 243 327 246 330 
rect 243 330 246 333 
rect 243 333 246 336 
rect 243 336 246 339 
rect 243 339 246 342 
rect 243 342 246 345 
rect 243 345 246 348 
rect 243 348 246 351 
rect 243 351 246 354 
rect 243 354 246 357 
rect 243 357 246 360 
rect 243 360 246 363 
rect 243 363 246 366 
rect 243 366 246 369 
rect 243 369 246 372 
rect 243 372 246 375 
rect 243 375 246 378 
rect 243 378 246 381 
rect 243 381 246 384 
rect 243 384 246 387 
rect 243 387 246 390 
rect 243 390 246 393 
rect 243 393 246 396 
rect 243 396 246 399 
rect 243 399 246 402 
rect 243 402 246 405 
rect 243 405 246 408 
rect 243 408 246 411 
rect 243 411 246 414 
rect 243 414 246 417 
rect 243 417 246 420 
rect 243 420 246 423 
rect 243 423 246 426 
rect 243 426 246 429 
rect 243 429 246 432 
rect 243 432 246 435 
rect 243 435 246 438 
rect 243 438 246 441 
rect 243 441 246 444 
rect 243 444 246 447 
rect 243 447 246 450 
rect 243 450 246 453 
rect 243 453 246 456 
rect 243 456 246 459 
rect 243 459 246 462 
rect 243 462 246 465 
rect 243 465 246 468 
rect 243 468 246 471 
rect 243 471 246 474 
rect 243 474 246 477 
rect 243 477 246 480 
rect 243 480 246 483 
rect 243 483 246 486 
rect 243 486 246 489 
rect 243 489 246 492 
rect 243 492 246 495 
rect 243 495 246 498 
rect 243 498 246 501 
rect 243 501 246 504 
rect 243 504 246 507 
rect 243 507 246 510 
rect 246 0 249 3 
rect 246 3 249 6 
rect 246 6 249 9 
rect 246 9 249 12 
rect 246 12 249 15 
rect 246 15 249 18 
rect 246 18 249 21 
rect 246 21 249 24 
rect 246 24 249 27 
rect 246 27 249 30 
rect 246 30 249 33 
rect 246 33 249 36 
rect 246 36 249 39 
rect 246 39 249 42 
rect 246 42 249 45 
rect 246 45 249 48 
rect 246 48 249 51 
rect 246 51 249 54 
rect 246 54 249 57 
rect 246 57 249 60 
rect 246 60 249 63 
rect 246 63 249 66 
rect 246 66 249 69 
rect 246 69 249 72 
rect 246 72 249 75 
rect 246 75 249 78 
rect 246 78 249 81 
rect 246 81 249 84 
rect 246 84 249 87 
rect 246 87 249 90 
rect 246 90 249 93 
rect 246 93 249 96 
rect 246 96 249 99 
rect 246 99 249 102 
rect 246 102 249 105 
rect 246 105 249 108 
rect 246 108 249 111 
rect 246 111 249 114 
rect 246 114 249 117 
rect 246 117 249 120 
rect 246 120 249 123 
rect 246 123 249 126 
rect 246 126 249 129 
rect 246 129 249 132 
rect 246 132 249 135 
rect 246 135 249 138 
rect 246 138 249 141 
rect 246 141 249 144 
rect 246 144 249 147 
rect 246 147 249 150 
rect 246 150 249 153 
rect 246 153 249 156 
rect 246 156 249 159 
rect 246 159 249 162 
rect 246 162 249 165 
rect 246 165 249 168 
rect 246 168 249 171 
rect 246 171 249 174 
rect 246 174 249 177 
rect 246 177 249 180 
rect 246 180 249 183 
rect 246 183 249 186 
rect 246 186 249 189 
rect 246 189 249 192 
rect 246 192 249 195 
rect 246 195 249 198 
rect 246 198 249 201 
rect 246 201 249 204 
rect 246 204 249 207 
rect 246 207 249 210 
rect 246 210 249 213 
rect 246 213 249 216 
rect 246 216 249 219 
rect 246 219 249 222 
rect 246 222 249 225 
rect 246 225 249 228 
rect 246 228 249 231 
rect 246 231 249 234 
rect 246 234 249 237 
rect 246 237 249 240 
rect 246 240 249 243 
rect 246 243 249 246 
rect 246 246 249 249 
rect 246 249 249 252 
rect 246 252 249 255 
rect 246 255 249 258 
rect 246 258 249 261 
rect 246 261 249 264 
rect 246 264 249 267 
rect 246 267 249 270 
rect 246 270 249 273 
rect 246 273 249 276 
rect 246 276 249 279 
rect 246 279 249 282 
rect 246 282 249 285 
rect 246 285 249 288 
rect 246 288 249 291 
rect 246 291 249 294 
rect 246 294 249 297 
rect 246 297 249 300 
rect 246 300 249 303 
rect 246 303 249 306 
rect 246 306 249 309 
rect 246 309 249 312 
rect 246 312 249 315 
rect 246 315 249 318 
rect 246 318 249 321 
rect 246 321 249 324 
rect 246 324 249 327 
rect 246 327 249 330 
rect 246 330 249 333 
rect 246 333 249 336 
rect 246 336 249 339 
rect 246 339 249 342 
rect 246 342 249 345 
rect 246 345 249 348 
rect 246 348 249 351 
rect 246 351 249 354 
rect 246 354 249 357 
rect 246 357 249 360 
rect 246 360 249 363 
rect 246 363 249 366 
rect 246 366 249 369 
rect 246 369 249 372 
rect 246 372 249 375 
rect 246 375 249 378 
rect 246 378 249 381 
rect 246 381 249 384 
rect 246 384 249 387 
rect 246 387 249 390 
rect 246 390 249 393 
rect 246 393 249 396 
rect 246 396 249 399 
rect 246 399 249 402 
rect 246 402 249 405 
rect 246 405 249 408 
rect 246 408 249 411 
rect 246 411 249 414 
rect 246 414 249 417 
rect 246 417 249 420 
rect 246 420 249 423 
rect 246 423 249 426 
rect 246 426 249 429 
rect 246 429 249 432 
rect 246 432 249 435 
rect 246 435 249 438 
rect 246 438 249 441 
rect 246 441 249 444 
rect 246 444 249 447 
rect 246 447 249 450 
rect 246 450 249 453 
rect 246 453 249 456 
rect 246 456 249 459 
rect 246 459 249 462 
rect 246 462 249 465 
rect 246 465 249 468 
rect 246 468 249 471 
rect 246 471 249 474 
rect 246 474 249 477 
rect 246 477 249 480 
rect 246 480 249 483 
rect 246 483 249 486 
rect 246 486 249 489 
rect 246 489 249 492 
rect 246 492 249 495 
rect 246 495 249 498 
rect 246 498 249 501 
rect 246 501 249 504 
rect 246 504 249 507 
rect 246 507 249 510 
rect 249 0 252 3 
rect 249 3 252 6 
rect 249 6 252 9 
rect 249 9 252 12 
rect 249 12 252 15 
rect 249 15 252 18 
rect 249 18 252 21 
rect 249 21 252 24 
rect 249 24 252 27 
rect 249 27 252 30 
rect 249 30 252 33 
rect 249 33 252 36 
rect 249 36 252 39 
rect 249 39 252 42 
rect 249 42 252 45 
rect 249 45 252 48 
rect 249 48 252 51 
rect 249 51 252 54 
rect 249 54 252 57 
rect 249 57 252 60 
rect 249 60 252 63 
rect 249 63 252 66 
rect 249 66 252 69 
rect 249 69 252 72 
rect 249 72 252 75 
rect 249 75 252 78 
rect 249 78 252 81 
rect 249 81 252 84 
rect 249 84 252 87 
rect 249 87 252 90 
rect 249 90 252 93 
rect 249 93 252 96 
rect 249 96 252 99 
rect 249 99 252 102 
rect 249 102 252 105 
rect 249 105 252 108 
rect 249 108 252 111 
rect 249 111 252 114 
rect 249 114 252 117 
rect 249 117 252 120 
rect 249 120 252 123 
rect 249 123 252 126 
rect 249 126 252 129 
rect 249 129 252 132 
rect 249 132 252 135 
rect 249 135 252 138 
rect 249 138 252 141 
rect 249 141 252 144 
rect 249 144 252 147 
rect 249 147 252 150 
rect 249 150 252 153 
rect 249 153 252 156 
rect 249 156 252 159 
rect 249 159 252 162 
rect 249 162 252 165 
rect 249 165 252 168 
rect 249 168 252 171 
rect 249 171 252 174 
rect 249 174 252 177 
rect 249 177 252 180 
rect 249 180 252 183 
rect 249 183 252 186 
rect 249 186 252 189 
rect 249 189 252 192 
rect 249 192 252 195 
rect 249 195 252 198 
rect 249 198 252 201 
rect 249 201 252 204 
rect 249 204 252 207 
rect 249 207 252 210 
rect 249 210 252 213 
rect 249 213 252 216 
rect 249 216 252 219 
rect 249 219 252 222 
rect 249 222 252 225 
rect 249 225 252 228 
rect 249 228 252 231 
rect 249 231 252 234 
rect 249 234 252 237 
rect 249 237 252 240 
rect 249 240 252 243 
rect 249 243 252 246 
rect 249 246 252 249 
rect 249 249 252 252 
rect 249 252 252 255 
rect 249 255 252 258 
rect 249 258 252 261 
rect 249 261 252 264 
rect 249 264 252 267 
rect 249 267 252 270 
rect 249 270 252 273 
rect 249 273 252 276 
rect 249 276 252 279 
rect 249 279 252 282 
rect 249 282 252 285 
rect 249 285 252 288 
rect 249 288 252 291 
rect 249 291 252 294 
rect 249 294 252 297 
rect 249 297 252 300 
rect 249 300 252 303 
rect 249 303 252 306 
rect 249 306 252 309 
rect 249 309 252 312 
rect 249 312 252 315 
rect 249 315 252 318 
rect 249 318 252 321 
rect 249 321 252 324 
rect 249 324 252 327 
rect 249 327 252 330 
rect 249 330 252 333 
rect 249 333 252 336 
rect 249 336 252 339 
rect 249 339 252 342 
rect 249 342 252 345 
rect 249 345 252 348 
rect 249 348 252 351 
rect 249 351 252 354 
rect 249 354 252 357 
rect 249 357 252 360 
rect 249 360 252 363 
rect 249 363 252 366 
rect 249 366 252 369 
rect 249 369 252 372 
rect 249 372 252 375 
rect 249 375 252 378 
rect 249 378 252 381 
rect 249 381 252 384 
rect 249 384 252 387 
rect 249 387 252 390 
rect 249 390 252 393 
rect 249 393 252 396 
rect 249 396 252 399 
rect 249 399 252 402 
rect 249 402 252 405 
rect 249 405 252 408 
rect 249 408 252 411 
rect 249 411 252 414 
rect 249 414 252 417 
rect 249 417 252 420 
rect 249 420 252 423 
rect 249 423 252 426 
rect 249 426 252 429 
rect 249 429 252 432 
rect 249 432 252 435 
rect 249 435 252 438 
rect 249 438 252 441 
rect 249 441 252 444 
rect 249 444 252 447 
rect 249 447 252 450 
rect 249 450 252 453 
rect 249 453 252 456 
rect 249 456 252 459 
rect 249 459 252 462 
rect 249 462 252 465 
rect 249 465 252 468 
rect 249 468 252 471 
rect 249 471 252 474 
rect 249 474 252 477 
rect 249 477 252 480 
rect 249 480 252 483 
rect 249 483 252 486 
rect 249 486 252 489 
rect 249 489 252 492 
rect 249 492 252 495 
rect 249 495 252 498 
rect 249 498 252 501 
rect 249 501 252 504 
rect 249 504 252 507 
rect 249 507 252 510 
rect 252 0 255 3 
rect 252 3 255 6 
rect 252 6 255 9 
rect 252 9 255 12 
rect 252 12 255 15 
rect 252 15 255 18 
rect 252 18 255 21 
rect 252 21 255 24 
rect 252 24 255 27 
rect 252 27 255 30 
rect 252 30 255 33 
rect 252 33 255 36 
rect 252 36 255 39 
rect 252 39 255 42 
rect 252 42 255 45 
rect 252 45 255 48 
rect 252 48 255 51 
rect 252 51 255 54 
rect 252 54 255 57 
rect 252 57 255 60 
rect 252 60 255 63 
rect 252 63 255 66 
rect 252 66 255 69 
rect 252 69 255 72 
rect 252 72 255 75 
rect 252 75 255 78 
rect 252 78 255 81 
rect 252 81 255 84 
rect 252 84 255 87 
rect 252 87 255 90 
rect 252 90 255 93 
rect 252 93 255 96 
rect 252 96 255 99 
rect 252 99 255 102 
rect 252 102 255 105 
rect 252 105 255 108 
rect 252 108 255 111 
rect 252 111 255 114 
rect 252 114 255 117 
rect 252 117 255 120 
rect 252 120 255 123 
rect 252 123 255 126 
rect 252 126 255 129 
rect 252 129 255 132 
rect 252 132 255 135 
rect 252 135 255 138 
rect 252 138 255 141 
rect 252 141 255 144 
rect 252 144 255 147 
rect 252 147 255 150 
rect 252 150 255 153 
rect 252 153 255 156 
rect 252 156 255 159 
rect 252 159 255 162 
rect 252 162 255 165 
rect 252 165 255 168 
rect 252 168 255 171 
rect 252 171 255 174 
rect 252 174 255 177 
rect 252 177 255 180 
rect 252 180 255 183 
rect 252 183 255 186 
rect 252 186 255 189 
rect 252 189 255 192 
rect 252 192 255 195 
rect 252 195 255 198 
rect 252 198 255 201 
rect 252 201 255 204 
rect 252 204 255 207 
rect 252 207 255 210 
rect 252 210 255 213 
rect 252 213 255 216 
rect 252 216 255 219 
rect 252 219 255 222 
rect 252 222 255 225 
rect 252 225 255 228 
rect 252 228 255 231 
rect 252 231 255 234 
rect 252 234 255 237 
rect 252 237 255 240 
rect 252 240 255 243 
rect 252 243 255 246 
rect 252 246 255 249 
rect 252 249 255 252 
rect 252 252 255 255 
rect 252 255 255 258 
rect 252 258 255 261 
rect 252 261 255 264 
rect 252 264 255 267 
rect 252 267 255 270 
rect 252 270 255 273 
rect 252 273 255 276 
rect 252 276 255 279 
rect 252 279 255 282 
rect 252 282 255 285 
rect 252 285 255 288 
rect 252 288 255 291 
rect 252 291 255 294 
rect 252 294 255 297 
rect 252 297 255 300 
rect 252 300 255 303 
rect 252 303 255 306 
rect 252 306 255 309 
rect 252 309 255 312 
rect 252 312 255 315 
rect 252 315 255 318 
rect 252 318 255 321 
rect 252 321 255 324 
rect 252 324 255 327 
rect 252 327 255 330 
rect 252 330 255 333 
rect 252 333 255 336 
rect 252 336 255 339 
rect 252 339 255 342 
rect 252 342 255 345 
rect 252 345 255 348 
rect 252 348 255 351 
rect 252 351 255 354 
rect 252 354 255 357 
rect 252 357 255 360 
rect 252 360 255 363 
rect 252 363 255 366 
rect 252 366 255 369 
rect 252 369 255 372 
rect 252 372 255 375 
rect 252 375 255 378 
rect 252 378 255 381 
rect 252 381 255 384 
rect 252 384 255 387 
rect 252 387 255 390 
rect 252 390 255 393 
rect 252 393 255 396 
rect 252 396 255 399 
rect 252 399 255 402 
rect 252 402 255 405 
rect 252 405 255 408 
rect 252 408 255 411 
rect 252 411 255 414 
rect 252 414 255 417 
rect 252 417 255 420 
rect 252 420 255 423 
rect 252 423 255 426 
rect 252 426 255 429 
rect 252 429 255 432 
rect 252 432 255 435 
rect 252 435 255 438 
rect 252 438 255 441 
rect 252 441 255 444 
rect 252 444 255 447 
rect 252 447 255 450 
rect 252 450 255 453 
rect 252 453 255 456 
rect 252 456 255 459 
rect 252 459 255 462 
rect 252 462 255 465 
rect 252 465 255 468 
rect 252 468 255 471 
rect 252 471 255 474 
rect 252 474 255 477 
rect 252 477 255 480 
rect 252 480 255 483 
rect 252 483 255 486 
rect 252 486 255 489 
rect 252 489 255 492 
rect 252 492 255 495 
rect 252 495 255 498 
rect 252 498 255 501 
rect 252 501 255 504 
rect 252 504 255 507 
rect 252 507 255 510 
rect 255 0 258 3 
rect 255 3 258 6 
rect 255 6 258 9 
rect 255 9 258 12 
rect 255 12 258 15 
rect 255 15 258 18 
rect 255 18 258 21 
rect 255 21 258 24 
rect 255 24 258 27 
rect 255 27 258 30 
rect 255 30 258 33 
rect 255 33 258 36 
rect 255 36 258 39 
rect 255 39 258 42 
rect 255 42 258 45 
rect 255 45 258 48 
rect 255 48 258 51 
rect 255 51 258 54 
rect 255 54 258 57 
rect 255 57 258 60 
rect 255 60 258 63 
rect 255 63 258 66 
rect 255 66 258 69 
rect 255 69 258 72 
rect 255 72 258 75 
rect 255 75 258 78 
rect 255 78 258 81 
rect 255 81 258 84 
rect 255 84 258 87 
rect 255 87 258 90 
rect 255 90 258 93 
rect 255 93 258 96 
rect 255 96 258 99 
rect 255 99 258 102 
rect 255 102 258 105 
rect 255 105 258 108 
rect 255 108 258 111 
rect 255 111 258 114 
rect 255 114 258 117 
rect 255 117 258 120 
rect 255 120 258 123 
rect 255 123 258 126 
rect 255 126 258 129 
rect 255 129 258 132 
rect 255 132 258 135 
rect 255 135 258 138 
rect 255 138 258 141 
rect 255 141 258 144 
rect 255 144 258 147 
rect 255 147 258 150 
rect 255 150 258 153 
rect 255 153 258 156 
rect 255 156 258 159 
rect 255 159 258 162 
rect 255 162 258 165 
rect 255 165 258 168 
rect 255 168 258 171 
rect 255 171 258 174 
rect 255 174 258 177 
rect 255 177 258 180 
rect 255 180 258 183 
rect 255 183 258 186 
rect 255 186 258 189 
rect 255 189 258 192 
rect 255 192 258 195 
rect 255 195 258 198 
rect 255 198 258 201 
rect 255 201 258 204 
rect 255 204 258 207 
rect 255 207 258 210 
rect 255 210 258 213 
rect 255 213 258 216 
rect 255 216 258 219 
rect 255 219 258 222 
rect 255 222 258 225 
rect 255 225 258 228 
rect 255 228 258 231 
rect 255 231 258 234 
rect 255 234 258 237 
rect 255 237 258 240 
rect 255 240 258 243 
rect 255 243 258 246 
rect 255 246 258 249 
rect 255 249 258 252 
rect 255 252 258 255 
rect 255 255 258 258 
rect 255 258 258 261 
rect 255 261 258 264 
rect 255 264 258 267 
rect 255 267 258 270 
rect 255 270 258 273 
rect 255 273 258 276 
rect 255 276 258 279 
rect 255 279 258 282 
rect 255 282 258 285 
rect 255 285 258 288 
rect 255 288 258 291 
rect 255 291 258 294 
rect 255 294 258 297 
rect 255 297 258 300 
rect 255 300 258 303 
rect 255 303 258 306 
rect 255 306 258 309 
rect 255 309 258 312 
rect 255 312 258 315 
rect 255 315 258 318 
rect 255 318 258 321 
rect 255 321 258 324 
rect 255 324 258 327 
rect 255 327 258 330 
rect 255 330 258 333 
rect 255 333 258 336 
rect 255 336 258 339 
rect 255 339 258 342 
rect 255 342 258 345 
rect 255 345 258 348 
rect 255 348 258 351 
rect 255 351 258 354 
rect 255 354 258 357 
rect 255 357 258 360 
rect 255 360 258 363 
rect 255 363 258 366 
rect 255 366 258 369 
rect 255 369 258 372 
rect 255 372 258 375 
rect 255 375 258 378 
rect 255 378 258 381 
rect 255 381 258 384 
rect 255 384 258 387 
rect 255 387 258 390 
rect 255 390 258 393 
rect 255 393 258 396 
rect 255 396 258 399 
rect 255 399 258 402 
rect 255 402 258 405 
rect 255 405 258 408 
rect 255 408 258 411 
rect 255 411 258 414 
rect 255 414 258 417 
rect 255 417 258 420 
rect 255 420 258 423 
rect 255 423 258 426 
rect 255 426 258 429 
rect 255 429 258 432 
rect 255 432 258 435 
rect 255 435 258 438 
rect 255 438 258 441 
rect 255 441 258 444 
rect 255 444 258 447 
rect 255 447 258 450 
rect 255 450 258 453 
rect 255 453 258 456 
rect 255 456 258 459 
rect 255 459 258 462 
rect 255 462 258 465 
rect 255 465 258 468 
rect 255 468 258 471 
rect 255 471 258 474 
rect 255 474 258 477 
rect 255 477 258 480 
rect 255 480 258 483 
rect 255 483 258 486 
rect 255 486 258 489 
rect 255 489 258 492 
rect 255 492 258 495 
rect 255 495 258 498 
rect 255 498 258 501 
rect 255 501 258 504 
rect 255 504 258 507 
rect 255 507 258 510 
rect 258 0 261 3 
rect 258 3 261 6 
rect 258 6 261 9 
rect 258 9 261 12 
rect 258 12 261 15 
rect 258 15 261 18 
rect 258 18 261 21 
rect 258 21 261 24 
rect 258 24 261 27 
rect 258 27 261 30 
rect 258 30 261 33 
rect 258 33 261 36 
rect 258 36 261 39 
rect 258 39 261 42 
rect 258 42 261 45 
rect 258 45 261 48 
rect 258 48 261 51 
rect 258 51 261 54 
rect 258 54 261 57 
rect 258 57 261 60 
rect 258 60 261 63 
rect 258 63 261 66 
rect 258 66 261 69 
rect 258 69 261 72 
rect 258 72 261 75 
rect 258 75 261 78 
rect 258 78 261 81 
rect 258 81 261 84 
rect 258 84 261 87 
rect 258 87 261 90 
rect 258 90 261 93 
rect 258 93 261 96 
rect 258 96 261 99 
rect 258 99 261 102 
rect 258 102 261 105 
rect 258 105 261 108 
rect 258 108 261 111 
rect 258 111 261 114 
rect 258 114 261 117 
rect 258 117 261 120 
rect 258 120 261 123 
rect 258 123 261 126 
rect 258 126 261 129 
rect 258 129 261 132 
rect 258 132 261 135 
rect 258 135 261 138 
rect 258 138 261 141 
rect 258 141 261 144 
rect 258 144 261 147 
rect 258 147 261 150 
rect 258 150 261 153 
rect 258 153 261 156 
rect 258 156 261 159 
rect 258 159 261 162 
rect 258 162 261 165 
rect 258 165 261 168 
rect 258 168 261 171 
rect 258 171 261 174 
rect 258 174 261 177 
rect 258 177 261 180 
rect 258 180 261 183 
rect 258 183 261 186 
rect 258 186 261 189 
rect 258 189 261 192 
rect 258 192 261 195 
rect 258 195 261 198 
rect 258 198 261 201 
rect 258 201 261 204 
rect 258 204 261 207 
rect 258 207 261 210 
rect 258 210 261 213 
rect 258 213 261 216 
rect 258 216 261 219 
rect 258 219 261 222 
rect 258 222 261 225 
rect 258 225 261 228 
rect 258 228 261 231 
rect 258 231 261 234 
rect 258 234 261 237 
rect 258 237 261 240 
rect 258 240 261 243 
rect 258 243 261 246 
rect 258 246 261 249 
rect 258 249 261 252 
rect 258 252 261 255 
rect 258 255 261 258 
rect 258 258 261 261 
rect 258 261 261 264 
rect 258 264 261 267 
rect 258 267 261 270 
rect 258 270 261 273 
rect 258 273 261 276 
rect 258 276 261 279 
rect 258 279 261 282 
rect 258 282 261 285 
rect 258 285 261 288 
rect 258 288 261 291 
rect 258 291 261 294 
rect 258 294 261 297 
rect 258 297 261 300 
rect 258 300 261 303 
rect 258 303 261 306 
rect 258 306 261 309 
rect 258 309 261 312 
rect 258 312 261 315 
rect 258 315 261 318 
rect 258 318 261 321 
rect 258 321 261 324 
rect 258 324 261 327 
rect 258 327 261 330 
rect 258 330 261 333 
rect 258 333 261 336 
rect 258 336 261 339 
rect 258 339 261 342 
rect 258 342 261 345 
rect 258 345 261 348 
rect 258 348 261 351 
rect 258 351 261 354 
rect 258 354 261 357 
rect 258 357 261 360 
rect 258 360 261 363 
rect 258 363 261 366 
rect 258 366 261 369 
rect 258 369 261 372 
rect 258 372 261 375 
rect 258 375 261 378 
rect 258 378 261 381 
rect 258 381 261 384 
rect 258 384 261 387 
rect 258 387 261 390 
rect 258 390 261 393 
rect 258 393 261 396 
rect 258 396 261 399 
rect 258 399 261 402 
rect 258 402 261 405 
rect 258 405 261 408 
rect 258 408 261 411 
rect 258 411 261 414 
rect 258 414 261 417 
rect 258 417 261 420 
rect 258 420 261 423 
rect 258 423 261 426 
rect 258 426 261 429 
rect 258 429 261 432 
rect 258 432 261 435 
rect 258 435 261 438 
rect 258 438 261 441 
rect 258 441 261 444 
rect 258 444 261 447 
rect 258 447 261 450 
rect 258 450 261 453 
rect 258 453 261 456 
rect 258 456 261 459 
rect 258 459 261 462 
rect 258 462 261 465 
rect 258 465 261 468 
rect 258 468 261 471 
rect 258 471 261 474 
rect 258 474 261 477 
rect 258 477 261 480 
rect 258 480 261 483 
rect 258 483 261 486 
rect 258 486 261 489 
rect 258 489 261 492 
rect 258 492 261 495 
rect 258 495 261 498 
rect 258 498 261 501 
rect 258 501 261 504 
rect 258 504 261 507 
rect 258 507 261 510 
rect 261 0 264 3 
rect 261 3 264 6 
rect 261 6 264 9 
rect 261 9 264 12 
rect 261 12 264 15 
rect 261 15 264 18 
rect 261 18 264 21 
rect 261 21 264 24 
rect 261 24 264 27 
rect 261 27 264 30 
rect 261 30 264 33 
rect 261 33 264 36 
rect 261 36 264 39 
rect 261 39 264 42 
rect 261 42 264 45 
rect 261 45 264 48 
rect 261 48 264 51 
rect 261 51 264 54 
rect 261 54 264 57 
rect 261 57 264 60 
rect 261 60 264 63 
rect 261 63 264 66 
rect 261 66 264 69 
rect 261 69 264 72 
rect 261 72 264 75 
rect 261 75 264 78 
rect 261 78 264 81 
rect 261 81 264 84 
rect 261 84 264 87 
rect 261 87 264 90 
rect 261 90 264 93 
rect 261 93 264 96 
rect 261 96 264 99 
rect 261 99 264 102 
rect 261 102 264 105 
rect 261 105 264 108 
rect 261 108 264 111 
rect 261 111 264 114 
rect 261 114 264 117 
rect 261 117 264 120 
rect 261 120 264 123 
rect 261 123 264 126 
rect 261 126 264 129 
rect 261 129 264 132 
rect 261 132 264 135 
rect 261 135 264 138 
rect 261 138 264 141 
rect 261 141 264 144 
rect 261 144 264 147 
rect 261 147 264 150 
rect 261 150 264 153 
rect 261 153 264 156 
rect 261 156 264 159 
rect 261 159 264 162 
rect 261 162 264 165 
rect 261 165 264 168 
rect 261 168 264 171 
rect 261 171 264 174 
rect 261 174 264 177 
rect 261 177 264 180 
rect 261 180 264 183 
rect 261 183 264 186 
rect 261 186 264 189 
rect 261 189 264 192 
rect 261 192 264 195 
rect 261 195 264 198 
rect 261 198 264 201 
rect 261 201 264 204 
rect 261 204 264 207 
rect 261 207 264 210 
rect 261 210 264 213 
rect 261 213 264 216 
rect 261 216 264 219 
rect 261 219 264 222 
rect 261 222 264 225 
rect 261 225 264 228 
rect 261 228 264 231 
rect 261 231 264 234 
rect 261 234 264 237 
rect 261 237 264 240 
rect 261 240 264 243 
rect 261 243 264 246 
rect 261 246 264 249 
rect 261 249 264 252 
rect 261 252 264 255 
rect 261 255 264 258 
rect 261 258 264 261 
rect 261 261 264 264 
rect 261 264 264 267 
rect 261 267 264 270 
rect 261 270 264 273 
rect 261 273 264 276 
rect 261 276 264 279 
rect 261 279 264 282 
rect 261 282 264 285 
rect 261 285 264 288 
rect 261 288 264 291 
rect 261 291 264 294 
rect 261 294 264 297 
rect 261 297 264 300 
rect 261 300 264 303 
rect 261 303 264 306 
rect 261 306 264 309 
rect 261 309 264 312 
rect 261 312 264 315 
rect 261 315 264 318 
rect 261 318 264 321 
rect 261 321 264 324 
rect 261 324 264 327 
rect 261 327 264 330 
rect 261 330 264 333 
rect 261 333 264 336 
rect 261 336 264 339 
rect 261 339 264 342 
rect 261 342 264 345 
rect 261 345 264 348 
rect 261 348 264 351 
rect 261 351 264 354 
rect 261 354 264 357 
rect 261 357 264 360 
rect 261 360 264 363 
rect 261 363 264 366 
rect 261 366 264 369 
rect 261 369 264 372 
rect 261 372 264 375 
rect 261 375 264 378 
rect 261 378 264 381 
rect 261 381 264 384 
rect 261 384 264 387 
rect 261 387 264 390 
rect 261 390 264 393 
rect 261 393 264 396 
rect 261 396 264 399 
rect 261 399 264 402 
rect 261 402 264 405 
rect 261 405 264 408 
rect 261 408 264 411 
rect 261 411 264 414 
rect 261 414 264 417 
rect 261 417 264 420 
rect 261 420 264 423 
rect 261 423 264 426 
rect 261 426 264 429 
rect 261 429 264 432 
rect 261 432 264 435 
rect 261 435 264 438 
rect 261 438 264 441 
rect 261 441 264 444 
rect 261 444 264 447 
rect 261 447 264 450 
rect 261 450 264 453 
rect 261 453 264 456 
rect 261 456 264 459 
rect 261 459 264 462 
rect 261 462 264 465 
rect 261 465 264 468 
rect 261 468 264 471 
rect 261 471 264 474 
rect 261 474 264 477 
rect 261 477 264 480 
rect 261 480 264 483 
rect 261 483 264 486 
rect 261 486 264 489 
rect 261 489 264 492 
rect 261 492 264 495 
rect 261 495 264 498 
rect 261 498 264 501 
rect 261 501 264 504 
rect 261 504 264 507 
rect 261 507 264 510 
rect 264 0 267 3 
rect 264 3 267 6 
rect 264 6 267 9 
rect 264 9 267 12 
rect 264 12 267 15 
rect 264 15 267 18 
rect 264 18 267 21 
rect 264 21 267 24 
rect 264 24 267 27 
rect 264 27 267 30 
rect 264 30 267 33 
rect 264 33 267 36 
rect 264 36 267 39 
rect 264 39 267 42 
rect 264 42 267 45 
rect 264 45 267 48 
rect 264 48 267 51 
rect 264 51 267 54 
rect 264 54 267 57 
rect 264 57 267 60 
rect 264 60 267 63 
rect 264 63 267 66 
rect 264 66 267 69 
rect 264 69 267 72 
rect 264 72 267 75 
rect 264 75 267 78 
rect 264 78 267 81 
rect 264 81 267 84 
rect 264 84 267 87 
rect 264 87 267 90 
rect 264 90 267 93 
rect 264 93 267 96 
rect 264 96 267 99 
rect 264 99 267 102 
rect 264 102 267 105 
rect 264 105 267 108 
rect 264 108 267 111 
rect 264 111 267 114 
rect 264 114 267 117 
rect 264 117 267 120 
rect 264 120 267 123 
rect 264 123 267 126 
rect 264 126 267 129 
rect 264 129 267 132 
rect 264 132 267 135 
rect 264 135 267 138 
rect 264 138 267 141 
rect 264 141 267 144 
rect 264 144 267 147 
rect 264 147 267 150 
rect 264 150 267 153 
rect 264 153 267 156 
rect 264 156 267 159 
rect 264 159 267 162 
rect 264 162 267 165 
rect 264 165 267 168 
rect 264 168 267 171 
rect 264 171 267 174 
rect 264 174 267 177 
rect 264 177 267 180 
rect 264 180 267 183 
rect 264 183 267 186 
rect 264 186 267 189 
rect 264 189 267 192 
rect 264 192 267 195 
rect 264 195 267 198 
rect 264 198 267 201 
rect 264 201 267 204 
rect 264 204 267 207 
rect 264 207 267 210 
rect 264 210 267 213 
rect 264 213 267 216 
rect 264 216 267 219 
rect 264 219 267 222 
rect 264 222 267 225 
rect 264 225 267 228 
rect 264 228 267 231 
rect 264 231 267 234 
rect 264 234 267 237 
rect 264 237 267 240 
rect 264 240 267 243 
rect 264 243 267 246 
rect 264 246 267 249 
rect 264 249 267 252 
rect 264 252 267 255 
rect 264 255 267 258 
rect 264 258 267 261 
rect 264 261 267 264 
rect 264 264 267 267 
rect 264 267 267 270 
rect 264 270 267 273 
rect 264 273 267 276 
rect 264 276 267 279 
rect 264 279 267 282 
rect 264 282 267 285 
rect 264 285 267 288 
rect 264 288 267 291 
rect 264 291 267 294 
rect 264 294 267 297 
rect 264 297 267 300 
rect 264 300 267 303 
rect 264 303 267 306 
rect 264 306 267 309 
rect 264 309 267 312 
rect 264 312 267 315 
rect 264 315 267 318 
rect 264 318 267 321 
rect 264 321 267 324 
rect 264 324 267 327 
rect 264 327 267 330 
rect 264 330 267 333 
rect 264 333 267 336 
rect 264 336 267 339 
rect 264 339 267 342 
rect 264 342 267 345 
rect 264 345 267 348 
rect 264 348 267 351 
rect 264 351 267 354 
rect 264 354 267 357 
rect 264 357 267 360 
rect 264 360 267 363 
rect 264 363 267 366 
rect 264 366 267 369 
rect 264 369 267 372 
rect 264 372 267 375 
rect 264 375 267 378 
rect 264 378 267 381 
rect 264 381 267 384 
rect 264 384 267 387 
rect 264 387 267 390 
rect 264 390 267 393 
rect 264 393 267 396 
rect 264 396 267 399 
rect 264 399 267 402 
rect 264 402 267 405 
rect 264 405 267 408 
rect 264 408 267 411 
rect 264 411 267 414 
rect 264 414 267 417 
rect 264 417 267 420 
rect 264 420 267 423 
rect 264 423 267 426 
rect 264 426 267 429 
rect 264 429 267 432 
rect 264 432 267 435 
rect 264 435 267 438 
rect 264 438 267 441 
rect 264 441 267 444 
rect 264 444 267 447 
rect 264 447 267 450 
rect 264 450 267 453 
rect 264 453 267 456 
rect 264 456 267 459 
rect 264 459 267 462 
rect 264 462 267 465 
rect 264 465 267 468 
rect 264 468 267 471 
rect 264 471 267 474 
rect 264 474 267 477 
rect 264 477 267 480 
rect 264 480 267 483 
rect 264 483 267 486 
rect 264 486 267 489 
rect 264 489 267 492 
rect 264 492 267 495 
rect 264 495 267 498 
rect 264 498 267 501 
rect 264 501 267 504 
rect 264 504 267 507 
rect 264 507 267 510 
rect 267 0 270 3 
rect 267 3 270 6 
rect 267 6 270 9 
rect 267 9 270 12 
rect 267 12 270 15 
rect 267 15 270 18 
rect 267 18 270 21 
rect 267 21 270 24 
rect 267 24 270 27 
rect 267 27 270 30 
rect 267 30 270 33 
rect 267 33 270 36 
rect 267 36 270 39 
rect 267 39 270 42 
rect 267 42 270 45 
rect 267 45 270 48 
rect 267 48 270 51 
rect 267 51 270 54 
rect 267 54 270 57 
rect 267 57 270 60 
rect 267 60 270 63 
rect 267 63 270 66 
rect 267 66 270 69 
rect 267 69 270 72 
rect 267 72 270 75 
rect 267 75 270 78 
rect 267 78 270 81 
rect 267 81 270 84 
rect 267 84 270 87 
rect 267 87 270 90 
rect 267 90 270 93 
rect 267 93 270 96 
rect 267 96 270 99 
rect 267 99 270 102 
rect 267 102 270 105 
rect 267 105 270 108 
rect 267 108 270 111 
rect 267 111 270 114 
rect 267 114 270 117 
rect 267 117 270 120 
rect 267 120 270 123 
rect 267 123 270 126 
rect 267 126 270 129 
rect 267 129 270 132 
rect 267 132 270 135 
rect 267 135 270 138 
rect 267 138 270 141 
rect 267 141 270 144 
rect 267 144 270 147 
rect 267 147 270 150 
rect 267 150 270 153 
rect 267 153 270 156 
rect 267 156 270 159 
rect 267 159 270 162 
rect 267 162 270 165 
rect 267 165 270 168 
rect 267 168 270 171 
rect 267 171 270 174 
rect 267 174 270 177 
rect 267 177 270 180 
rect 267 180 270 183 
rect 267 183 270 186 
rect 267 186 270 189 
rect 267 189 270 192 
rect 267 192 270 195 
rect 267 195 270 198 
rect 267 198 270 201 
rect 267 201 270 204 
rect 267 204 270 207 
rect 267 207 270 210 
rect 267 210 270 213 
rect 267 213 270 216 
rect 267 216 270 219 
rect 267 219 270 222 
rect 267 222 270 225 
rect 267 225 270 228 
rect 267 228 270 231 
rect 267 231 270 234 
rect 267 234 270 237 
rect 267 237 270 240 
rect 267 240 270 243 
rect 267 243 270 246 
rect 267 246 270 249 
rect 267 249 270 252 
rect 267 252 270 255 
rect 267 255 270 258 
rect 267 258 270 261 
rect 267 261 270 264 
rect 267 264 270 267 
rect 267 267 270 270 
rect 267 270 270 273 
rect 267 273 270 276 
rect 267 276 270 279 
rect 267 279 270 282 
rect 267 282 270 285 
rect 267 285 270 288 
rect 267 288 270 291 
rect 267 291 270 294 
rect 267 294 270 297 
rect 267 297 270 300 
rect 267 300 270 303 
rect 267 303 270 306 
rect 267 306 270 309 
rect 267 309 270 312 
rect 267 312 270 315 
rect 267 315 270 318 
rect 267 318 270 321 
rect 267 321 270 324 
rect 267 324 270 327 
rect 267 327 270 330 
rect 267 330 270 333 
rect 267 333 270 336 
rect 267 336 270 339 
rect 267 339 270 342 
rect 267 342 270 345 
rect 267 345 270 348 
rect 267 348 270 351 
rect 267 351 270 354 
rect 267 354 270 357 
rect 267 357 270 360 
rect 267 360 270 363 
rect 267 363 270 366 
rect 267 366 270 369 
rect 267 369 270 372 
rect 267 372 270 375 
rect 267 375 270 378 
rect 267 378 270 381 
rect 267 381 270 384 
rect 267 384 270 387 
rect 267 387 270 390 
rect 267 390 270 393 
rect 267 393 270 396 
rect 267 396 270 399 
rect 267 399 270 402 
rect 267 402 270 405 
rect 267 405 270 408 
rect 267 408 270 411 
rect 267 411 270 414 
rect 267 414 270 417 
rect 267 417 270 420 
rect 267 420 270 423 
rect 267 423 270 426 
rect 267 426 270 429 
rect 267 429 270 432 
rect 267 432 270 435 
rect 267 435 270 438 
rect 267 438 270 441 
rect 267 441 270 444 
rect 267 444 270 447 
rect 267 447 270 450 
rect 267 450 270 453 
rect 267 453 270 456 
rect 267 456 270 459 
rect 267 459 270 462 
rect 267 462 270 465 
rect 267 465 270 468 
rect 267 468 270 471 
rect 267 471 270 474 
rect 267 474 270 477 
rect 267 477 270 480 
rect 267 480 270 483 
rect 267 483 270 486 
rect 267 486 270 489 
rect 267 489 270 492 
rect 267 492 270 495 
rect 267 495 270 498 
rect 267 498 270 501 
rect 267 501 270 504 
rect 267 504 270 507 
rect 267 507 270 510 
rect 270 0 273 3 
rect 270 3 273 6 
rect 270 6 273 9 
rect 270 9 273 12 
rect 270 12 273 15 
rect 270 15 273 18 
rect 270 18 273 21 
rect 270 21 273 24 
rect 270 24 273 27 
rect 270 27 273 30 
rect 270 30 273 33 
rect 270 33 273 36 
rect 270 36 273 39 
rect 270 39 273 42 
rect 270 42 273 45 
rect 270 45 273 48 
rect 270 48 273 51 
rect 270 51 273 54 
rect 270 54 273 57 
rect 270 57 273 60 
rect 270 60 273 63 
rect 270 63 273 66 
rect 270 66 273 69 
rect 270 69 273 72 
rect 270 72 273 75 
rect 270 75 273 78 
rect 270 78 273 81 
rect 270 81 273 84 
rect 270 84 273 87 
rect 270 87 273 90 
rect 270 90 273 93 
rect 270 93 273 96 
rect 270 96 273 99 
rect 270 99 273 102 
rect 270 102 273 105 
rect 270 105 273 108 
rect 270 108 273 111 
rect 270 111 273 114 
rect 270 114 273 117 
rect 270 117 273 120 
rect 270 120 273 123 
rect 270 123 273 126 
rect 270 126 273 129 
rect 270 129 273 132 
rect 270 132 273 135 
rect 270 135 273 138 
rect 270 138 273 141 
rect 270 141 273 144 
rect 270 144 273 147 
rect 270 147 273 150 
rect 270 150 273 153 
rect 270 153 273 156 
rect 270 156 273 159 
rect 270 159 273 162 
rect 270 162 273 165 
rect 270 165 273 168 
rect 270 168 273 171 
rect 270 171 273 174 
rect 270 174 273 177 
rect 270 177 273 180 
rect 270 180 273 183 
rect 270 183 273 186 
rect 270 186 273 189 
rect 270 189 273 192 
rect 270 192 273 195 
rect 270 195 273 198 
rect 270 198 273 201 
rect 270 201 273 204 
rect 270 204 273 207 
rect 270 207 273 210 
rect 270 210 273 213 
rect 270 213 273 216 
rect 270 216 273 219 
rect 270 219 273 222 
rect 270 222 273 225 
rect 270 225 273 228 
rect 270 228 273 231 
rect 270 231 273 234 
rect 270 234 273 237 
rect 270 237 273 240 
rect 270 240 273 243 
rect 270 243 273 246 
rect 270 246 273 249 
rect 270 249 273 252 
rect 270 252 273 255 
rect 270 255 273 258 
rect 270 258 273 261 
rect 270 261 273 264 
rect 270 264 273 267 
rect 270 267 273 270 
rect 270 270 273 273 
rect 270 273 273 276 
rect 270 276 273 279 
rect 270 279 273 282 
rect 270 282 273 285 
rect 270 285 273 288 
rect 270 288 273 291 
rect 270 291 273 294 
rect 270 294 273 297 
rect 270 297 273 300 
rect 270 300 273 303 
rect 270 303 273 306 
rect 270 306 273 309 
rect 270 309 273 312 
rect 270 312 273 315 
rect 270 315 273 318 
rect 270 318 273 321 
rect 270 321 273 324 
rect 270 324 273 327 
rect 270 327 273 330 
rect 270 330 273 333 
rect 270 333 273 336 
rect 270 336 273 339 
rect 270 339 273 342 
rect 270 342 273 345 
rect 270 345 273 348 
rect 270 348 273 351 
rect 270 351 273 354 
rect 270 354 273 357 
rect 270 357 273 360 
rect 270 360 273 363 
rect 270 363 273 366 
rect 270 366 273 369 
rect 270 369 273 372 
rect 270 372 273 375 
rect 270 375 273 378 
rect 270 378 273 381 
rect 270 381 273 384 
rect 270 384 273 387 
rect 270 387 273 390 
rect 270 390 273 393 
rect 270 393 273 396 
rect 270 396 273 399 
rect 270 399 273 402 
rect 270 402 273 405 
rect 270 405 273 408 
rect 270 408 273 411 
rect 270 411 273 414 
rect 270 414 273 417 
rect 270 417 273 420 
rect 270 420 273 423 
rect 270 423 273 426 
rect 270 426 273 429 
rect 270 429 273 432 
rect 270 432 273 435 
rect 270 435 273 438 
rect 270 438 273 441 
rect 270 441 273 444 
rect 270 444 273 447 
rect 270 447 273 450 
rect 270 450 273 453 
rect 270 453 273 456 
rect 270 456 273 459 
rect 270 459 273 462 
rect 270 462 273 465 
rect 270 465 273 468 
rect 270 468 273 471 
rect 270 471 273 474 
rect 270 474 273 477 
rect 270 477 273 480 
rect 270 480 273 483 
rect 270 483 273 486 
rect 270 486 273 489 
rect 270 489 273 492 
rect 270 492 273 495 
rect 270 495 273 498 
rect 270 498 273 501 
rect 270 501 273 504 
rect 270 504 273 507 
rect 270 507 273 510 
rect 273 0 276 3 
rect 273 3 276 6 
rect 273 6 276 9 
rect 273 9 276 12 
rect 273 12 276 15 
rect 273 15 276 18 
rect 273 18 276 21 
rect 273 21 276 24 
rect 273 24 276 27 
rect 273 27 276 30 
rect 273 30 276 33 
rect 273 33 276 36 
rect 273 36 276 39 
rect 273 39 276 42 
rect 273 42 276 45 
rect 273 45 276 48 
rect 273 48 276 51 
rect 273 51 276 54 
rect 273 54 276 57 
rect 273 57 276 60 
rect 273 60 276 63 
rect 273 63 276 66 
rect 273 66 276 69 
rect 273 69 276 72 
rect 273 72 276 75 
rect 273 75 276 78 
rect 273 78 276 81 
rect 273 81 276 84 
rect 273 84 276 87 
rect 273 87 276 90 
rect 273 90 276 93 
rect 273 93 276 96 
rect 273 96 276 99 
rect 273 99 276 102 
rect 273 102 276 105 
rect 273 105 276 108 
rect 273 108 276 111 
rect 273 111 276 114 
rect 273 114 276 117 
rect 273 117 276 120 
rect 273 120 276 123 
rect 273 123 276 126 
rect 273 126 276 129 
rect 273 129 276 132 
rect 273 132 276 135 
rect 273 135 276 138 
rect 273 138 276 141 
rect 273 141 276 144 
rect 273 144 276 147 
rect 273 147 276 150 
rect 273 150 276 153 
rect 273 153 276 156 
rect 273 156 276 159 
rect 273 159 276 162 
rect 273 162 276 165 
rect 273 165 276 168 
rect 273 168 276 171 
rect 273 171 276 174 
rect 273 174 276 177 
rect 273 177 276 180 
rect 273 180 276 183 
rect 273 183 276 186 
rect 273 186 276 189 
rect 273 189 276 192 
rect 273 192 276 195 
rect 273 195 276 198 
rect 273 198 276 201 
rect 273 201 276 204 
rect 273 204 276 207 
rect 273 207 276 210 
rect 273 210 276 213 
rect 273 213 276 216 
rect 273 216 276 219 
rect 273 219 276 222 
rect 273 222 276 225 
rect 273 225 276 228 
rect 273 228 276 231 
rect 273 231 276 234 
rect 273 234 276 237 
rect 273 237 276 240 
rect 273 240 276 243 
rect 273 243 276 246 
rect 273 246 276 249 
rect 273 249 276 252 
rect 273 252 276 255 
rect 273 255 276 258 
rect 273 258 276 261 
rect 273 261 276 264 
rect 273 264 276 267 
rect 273 267 276 270 
rect 273 270 276 273 
rect 273 273 276 276 
rect 273 276 276 279 
rect 273 279 276 282 
rect 273 282 276 285 
rect 273 285 276 288 
rect 273 288 276 291 
rect 273 291 276 294 
rect 273 294 276 297 
rect 273 297 276 300 
rect 273 300 276 303 
rect 273 303 276 306 
rect 273 306 276 309 
rect 273 309 276 312 
rect 273 312 276 315 
rect 273 315 276 318 
rect 273 318 276 321 
rect 273 321 276 324 
rect 273 324 276 327 
rect 273 327 276 330 
rect 273 330 276 333 
rect 273 333 276 336 
rect 273 336 276 339 
rect 273 339 276 342 
rect 273 342 276 345 
rect 273 345 276 348 
rect 273 348 276 351 
rect 273 351 276 354 
rect 273 354 276 357 
rect 273 357 276 360 
rect 273 360 276 363 
rect 273 363 276 366 
rect 273 366 276 369 
rect 273 369 276 372 
rect 273 372 276 375 
rect 273 375 276 378 
rect 273 378 276 381 
rect 273 381 276 384 
rect 273 384 276 387 
rect 273 387 276 390 
rect 273 390 276 393 
rect 273 393 276 396 
rect 273 396 276 399 
rect 273 399 276 402 
rect 273 402 276 405 
rect 273 405 276 408 
rect 273 408 276 411 
rect 273 411 276 414 
rect 273 414 276 417 
rect 273 417 276 420 
rect 273 420 276 423 
rect 273 423 276 426 
rect 273 426 276 429 
rect 273 429 276 432 
rect 273 432 276 435 
rect 273 435 276 438 
rect 273 438 276 441 
rect 273 441 276 444 
rect 273 444 276 447 
rect 273 447 276 450 
rect 273 450 276 453 
rect 273 453 276 456 
rect 273 456 276 459 
rect 273 459 276 462 
rect 273 462 276 465 
rect 273 465 276 468 
rect 273 468 276 471 
rect 273 471 276 474 
rect 273 474 276 477 
rect 273 477 276 480 
rect 273 480 276 483 
rect 273 483 276 486 
rect 273 486 276 489 
rect 273 489 276 492 
rect 273 492 276 495 
rect 273 495 276 498 
rect 273 498 276 501 
rect 273 501 276 504 
rect 273 504 276 507 
rect 273 507 276 510 
rect 276 0 279 3 
rect 276 3 279 6 
rect 276 6 279 9 
rect 276 9 279 12 
rect 276 12 279 15 
rect 276 15 279 18 
rect 276 18 279 21 
rect 276 21 279 24 
rect 276 24 279 27 
rect 276 27 279 30 
rect 276 30 279 33 
rect 276 33 279 36 
rect 276 36 279 39 
rect 276 39 279 42 
rect 276 42 279 45 
rect 276 45 279 48 
rect 276 48 279 51 
rect 276 51 279 54 
rect 276 54 279 57 
rect 276 57 279 60 
rect 276 60 279 63 
rect 276 63 279 66 
rect 276 66 279 69 
rect 276 69 279 72 
rect 276 72 279 75 
rect 276 75 279 78 
rect 276 78 279 81 
rect 276 81 279 84 
rect 276 84 279 87 
rect 276 87 279 90 
rect 276 90 279 93 
rect 276 93 279 96 
rect 276 96 279 99 
rect 276 99 279 102 
rect 276 102 279 105 
rect 276 105 279 108 
rect 276 108 279 111 
rect 276 111 279 114 
rect 276 114 279 117 
rect 276 117 279 120 
rect 276 120 279 123 
rect 276 123 279 126 
rect 276 126 279 129 
rect 276 129 279 132 
rect 276 132 279 135 
rect 276 135 279 138 
rect 276 138 279 141 
rect 276 141 279 144 
rect 276 144 279 147 
rect 276 147 279 150 
rect 276 150 279 153 
rect 276 153 279 156 
rect 276 156 279 159 
rect 276 159 279 162 
rect 276 162 279 165 
rect 276 165 279 168 
rect 276 168 279 171 
rect 276 171 279 174 
rect 276 174 279 177 
rect 276 177 279 180 
rect 276 180 279 183 
rect 276 183 279 186 
rect 276 186 279 189 
rect 276 189 279 192 
rect 276 192 279 195 
rect 276 195 279 198 
rect 276 198 279 201 
rect 276 201 279 204 
rect 276 204 279 207 
rect 276 207 279 210 
rect 276 210 279 213 
rect 276 213 279 216 
rect 276 216 279 219 
rect 276 219 279 222 
rect 276 222 279 225 
rect 276 225 279 228 
rect 276 228 279 231 
rect 276 231 279 234 
rect 276 234 279 237 
rect 276 237 279 240 
rect 276 240 279 243 
rect 276 243 279 246 
rect 276 246 279 249 
rect 276 249 279 252 
rect 276 252 279 255 
rect 276 255 279 258 
rect 276 258 279 261 
rect 276 261 279 264 
rect 276 264 279 267 
rect 276 267 279 270 
rect 276 270 279 273 
rect 276 273 279 276 
rect 276 276 279 279 
rect 276 279 279 282 
rect 276 282 279 285 
rect 276 285 279 288 
rect 276 288 279 291 
rect 276 291 279 294 
rect 276 294 279 297 
rect 276 297 279 300 
rect 276 300 279 303 
rect 276 303 279 306 
rect 276 306 279 309 
rect 276 309 279 312 
rect 276 312 279 315 
rect 276 315 279 318 
rect 276 318 279 321 
rect 276 321 279 324 
rect 276 324 279 327 
rect 276 327 279 330 
rect 276 330 279 333 
rect 276 333 279 336 
rect 276 336 279 339 
rect 276 339 279 342 
rect 276 342 279 345 
rect 276 345 279 348 
rect 276 348 279 351 
rect 276 351 279 354 
rect 276 354 279 357 
rect 276 357 279 360 
rect 276 360 279 363 
rect 276 363 279 366 
rect 276 366 279 369 
rect 276 369 279 372 
rect 276 372 279 375 
rect 276 375 279 378 
rect 276 378 279 381 
rect 276 381 279 384 
rect 276 384 279 387 
rect 276 387 279 390 
rect 276 390 279 393 
rect 276 393 279 396 
rect 276 396 279 399 
rect 276 399 279 402 
rect 276 402 279 405 
rect 276 405 279 408 
rect 276 408 279 411 
rect 276 411 279 414 
rect 276 414 279 417 
rect 276 417 279 420 
rect 276 420 279 423 
rect 276 423 279 426 
rect 276 426 279 429 
rect 276 429 279 432 
rect 276 432 279 435 
rect 276 435 279 438 
rect 276 438 279 441 
rect 276 441 279 444 
rect 276 444 279 447 
rect 276 447 279 450 
rect 276 450 279 453 
rect 276 453 279 456 
rect 276 456 279 459 
rect 276 459 279 462 
rect 276 462 279 465 
rect 276 465 279 468 
rect 276 468 279 471 
rect 276 471 279 474 
rect 276 474 279 477 
rect 276 477 279 480 
rect 276 480 279 483 
rect 276 483 279 486 
rect 276 486 279 489 
rect 276 489 279 492 
rect 276 492 279 495 
rect 276 495 279 498 
rect 276 498 279 501 
rect 276 501 279 504 
rect 276 504 279 507 
rect 276 507 279 510 
rect 279 0 282 3 
rect 279 3 282 6 
rect 279 6 282 9 
rect 279 9 282 12 
rect 279 12 282 15 
rect 279 15 282 18 
rect 279 18 282 21 
rect 279 21 282 24 
rect 279 24 282 27 
rect 279 27 282 30 
rect 279 30 282 33 
rect 279 33 282 36 
rect 279 36 282 39 
rect 279 39 282 42 
rect 279 42 282 45 
rect 279 45 282 48 
rect 279 48 282 51 
rect 279 51 282 54 
rect 279 54 282 57 
rect 279 57 282 60 
rect 279 60 282 63 
rect 279 63 282 66 
rect 279 66 282 69 
rect 279 69 282 72 
rect 279 72 282 75 
rect 279 75 282 78 
rect 279 78 282 81 
rect 279 81 282 84 
rect 279 84 282 87 
rect 279 87 282 90 
rect 279 90 282 93 
rect 279 93 282 96 
rect 279 96 282 99 
rect 279 99 282 102 
rect 279 102 282 105 
rect 279 105 282 108 
rect 279 108 282 111 
rect 279 111 282 114 
rect 279 114 282 117 
rect 279 117 282 120 
rect 279 120 282 123 
rect 279 123 282 126 
rect 279 126 282 129 
rect 279 129 282 132 
rect 279 132 282 135 
rect 279 135 282 138 
rect 279 138 282 141 
rect 279 141 282 144 
rect 279 144 282 147 
rect 279 147 282 150 
rect 279 150 282 153 
rect 279 153 282 156 
rect 279 156 282 159 
rect 279 159 282 162 
rect 279 162 282 165 
rect 279 165 282 168 
rect 279 168 282 171 
rect 279 171 282 174 
rect 279 174 282 177 
rect 279 177 282 180 
rect 279 180 282 183 
rect 279 183 282 186 
rect 279 186 282 189 
rect 279 189 282 192 
rect 279 192 282 195 
rect 279 195 282 198 
rect 279 198 282 201 
rect 279 201 282 204 
rect 279 204 282 207 
rect 279 207 282 210 
rect 279 210 282 213 
rect 279 213 282 216 
rect 279 216 282 219 
rect 279 219 282 222 
rect 279 222 282 225 
rect 279 225 282 228 
rect 279 228 282 231 
rect 279 231 282 234 
rect 279 234 282 237 
rect 279 237 282 240 
rect 279 240 282 243 
rect 279 243 282 246 
rect 279 246 282 249 
rect 279 249 282 252 
rect 279 252 282 255 
rect 279 255 282 258 
rect 279 258 282 261 
rect 279 261 282 264 
rect 279 264 282 267 
rect 279 267 282 270 
rect 279 270 282 273 
rect 279 273 282 276 
rect 279 276 282 279 
rect 279 279 282 282 
rect 279 282 282 285 
rect 279 285 282 288 
rect 279 288 282 291 
rect 279 291 282 294 
rect 279 294 282 297 
rect 279 297 282 300 
rect 279 300 282 303 
rect 279 303 282 306 
rect 279 306 282 309 
rect 279 309 282 312 
rect 279 312 282 315 
rect 279 315 282 318 
rect 279 318 282 321 
rect 279 321 282 324 
rect 279 324 282 327 
rect 279 327 282 330 
rect 279 330 282 333 
rect 279 333 282 336 
rect 279 336 282 339 
rect 279 339 282 342 
rect 279 342 282 345 
rect 279 345 282 348 
rect 279 348 282 351 
rect 279 351 282 354 
rect 279 354 282 357 
rect 279 357 282 360 
rect 279 360 282 363 
rect 279 363 282 366 
rect 279 366 282 369 
rect 279 369 282 372 
rect 279 372 282 375 
rect 279 375 282 378 
rect 279 378 282 381 
rect 279 381 282 384 
rect 279 384 282 387 
rect 279 387 282 390 
rect 279 390 282 393 
rect 279 393 282 396 
rect 279 396 282 399 
rect 279 399 282 402 
rect 279 402 282 405 
rect 279 405 282 408 
rect 279 408 282 411 
rect 279 411 282 414 
rect 279 414 282 417 
rect 279 417 282 420 
rect 279 420 282 423 
rect 279 423 282 426 
rect 279 426 282 429 
rect 279 429 282 432 
rect 279 432 282 435 
rect 279 435 282 438 
rect 279 438 282 441 
rect 279 441 282 444 
rect 279 444 282 447 
rect 279 447 282 450 
rect 279 450 282 453 
rect 279 453 282 456 
rect 279 456 282 459 
rect 279 459 282 462 
rect 279 462 282 465 
rect 279 465 282 468 
rect 279 468 282 471 
rect 279 471 282 474 
rect 279 474 282 477 
rect 279 477 282 480 
rect 279 480 282 483 
rect 279 483 282 486 
rect 279 486 282 489 
rect 279 489 282 492 
rect 279 492 282 495 
rect 279 495 282 498 
rect 279 498 282 501 
rect 279 501 282 504 
rect 279 504 282 507 
rect 279 507 282 510 
rect 282 0 285 3 
rect 282 3 285 6 
rect 282 6 285 9 
rect 282 9 285 12 
rect 282 12 285 15 
rect 282 15 285 18 
rect 282 18 285 21 
rect 282 21 285 24 
rect 282 24 285 27 
rect 282 27 285 30 
rect 282 30 285 33 
rect 282 33 285 36 
rect 282 36 285 39 
rect 282 39 285 42 
rect 282 42 285 45 
rect 282 45 285 48 
rect 282 48 285 51 
rect 282 51 285 54 
rect 282 54 285 57 
rect 282 57 285 60 
rect 282 60 285 63 
rect 282 63 285 66 
rect 282 66 285 69 
rect 282 69 285 72 
rect 282 72 285 75 
rect 282 75 285 78 
rect 282 78 285 81 
rect 282 81 285 84 
rect 282 84 285 87 
rect 282 87 285 90 
rect 282 90 285 93 
rect 282 93 285 96 
rect 282 96 285 99 
rect 282 99 285 102 
rect 282 102 285 105 
rect 282 105 285 108 
rect 282 108 285 111 
rect 282 111 285 114 
rect 282 114 285 117 
rect 282 117 285 120 
rect 282 120 285 123 
rect 282 123 285 126 
rect 282 126 285 129 
rect 282 129 285 132 
rect 282 132 285 135 
rect 282 135 285 138 
rect 282 138 285 141 
rect 282 141 285 144 
rect 282 144 285 147 
rect 282 147 285 150 
rect 282 150 285 153 
rect 282 153 285 156 
rect 282 156 285 159 
rect 282 159 285 162 
rect 282 162 285 165 
rect 282 165 285 168 
rect 282 168 285 171 
rect 282 171 285 174 
rect 282 174 285 177 
rect 282 177 285 180 
rect 282 180 285 183 
rect 282 183 285 186 
rect 282 186 285 189 
rect 282 189 285 192 
rect 282 192 285 195 
rect 282 195 285 198 
rect 282 198 285 201 
rect 282 201 285 204 
rect 282 204 285 207 
rect 282 207 285 210 
rect 282 210 285 213 
rect 282 213 285 216 
rect 282 216 285 219 
rect 282 219 285 222 
rect 282 222 285 225 
rect 282 225 285 228 
rect 282 228 285 231 
rect 282 231 285 234 
rect 282 234 285 237 
rect 282 237 285 240 
rect 282 240 285 243 
rect 282 243 285 246 
rect 282 246 285 249 
rect 282 249 285 252 
rect 282 252 285 255 
rect 282 255 285 258 
rect 282 258 285 261 
rect 282 261 285 264 
rect 282 264 285 267 
rect 282 267 285 270 
rect 282 270 285 273 
rect 282 273 285 276 
rect 282 276 285 279 
rect 282 279 285 282 
rect 282 282 285 285 
rect 282 285 285 288 
rect 282 288 285 291 
rect 282 291 285 294 
rect 282 294 285 297 
rect 282 297 285 300 
rect 282 300 285 303 
rect 282 303 285 306 
rect 282 306 285 309 
rect 282 309 285 312 
rect 282 312 285 315 
rect 282 315 285 318 
rect 282 318 285 321 
rect 282 321 285 324 
rect 282 324 285 327 
rect 282 327 285 330 
rect 282 330 285 333 
rect 282 333 285 336 
rect 282 336 285 339 
rect 282 339 285 342 
rect 282 342 285 345 
rect 282 345 285 348 
rect 282 348 285 351 
rect 282 351 285 354 
rect 282 354 285 357 
rect 282 357 285 360 
rect 282 360 285 363 
rect 282 363 285 366 
rect 282 366 285 369 
rect 282 369 285 372 
rect 282 372 285 375 
rect 282 375 285 378 
rect 282 378 285 381 
rect 282 381 285 384 
rect 282 384 285 387 
rect 282 387 285 390 
rect 282 390 285 393 
rect 282 393 285 396 
rect 282 396 285 399 
rect 282 399 285 402 
rect 282 402 285 405 
rect 282 405 285 408 
rect 282 408 285 411 
rect 282 411 285 414 
rect 282 414 285 417 
rect 282 417 285 420 
rect 282 420 285 423 
rect 282 423 285 426 
rect 282 426 285 429 
rect 282 429 285 432 
rect 282 432 285 435 
rect 282 435 285 438 
rect 282 438 285 441 
rect 282 441 285 444 
rect 282 444 285 447 
rect 282 447 285 450 
rect 282 450 285 453 
rect 282 453 285 456 
rect 282 456 285 459 
rect 282 459 285 462 
rect 282 462 285 465 
rect 282 465 285 468 
rect 282 468 285 471 
rect 282 471 285 474 
rect 282 474 285 477 
rect 282 477 285 480 
rect 282 480 285 483 
rect 282 483 285 486 
rect 282 486 285 489 
rect 282 489 285 492 
rect 282 492 285 495 
rect 282 495 285 498 
rect 282 498 285 501 
rect 282 501 285 504 
rect 282 504 285 507 
rect 282 507 285 510 
rect 285 0 288 3 
rect 285 3 288 6 
rect 285 6 288 9 
rect 285 9 288 12 
rect 285 12 288 15 
rect 285 15 288 18 
rect 285 18 288 21 
rect 285 21 288 24 
rect 285 24 288 27 
rect 285 27 288 30 
rect 285 30 288 33 
rect 285 33 288 36 
rect 285 36 288 39 
rect 285 39 288 42 
rect 285 42 288 45 
rect 285 45 288 48 
rect 285 48 288 51 
rect 285 51 288 54 
rect 285 54 288 57 
rect 285 57 288 60 
rect 285 60 288 63 
rect 285 63 288 66 
rect 285 66 288 69 
rect 285 69 288 72 
rect 285 72 288 75 
rect 285 75 288 78 
rect 285 78 288 81 
rect 285 81 288 84 
rect 285 84 288 87 
rect 285 87 288 90 
rect 285 90 288 93 
rect 285 93 288 96 
rect 285 96 288 99 
rect 285 99 288 102 
rect 285 102 288 105 
rect 285 105 288 108 
rect 285 108 288 111 
rect 285 111 288 114 
rect 285 114 288 117 
rect 285 117 288 120 
rect 285 120 288 123 
rect 285 123 288 126 
rect 285 126 288 129 
rect 285 129 288 132 
rect 285 132 288 135 
rect 285 135 288 138 
rect 285 138 288 141 
rect 285 141 288 144 
rect 285 144 288 147 
rect 285 147 288 150 
rect 285 150 288 153 
rect 285 153 288 156 
rect 285 156 288 159 
rect 285 159 288 162 
rect 285 162 288 165 
rect 285 165 288 168 
rect 285 168 288 171 
rect 285 171 288 174 
rect 285 174 288 177 
rect 285 177 288 180 
rect 285 180 288 183 
rect 285 183 288 186 
rect 285 186 288 189 
rect 285 189 288 192 
rect 285 192 288 195 
rect 285 195 288 198 
rect 285 198 288 201 
rect 285 201 288 204 
rect 285 204 288 207 
rect 285 207 288 210 
rect 285 210 288 213 
rect 285 213 288 216 
rect 285 216 288 219 
rect 285 219 288 222 
rect 285 222 288 225 
rect 285 225 288 228 
rect 285 228 288 231 
rect 285 231 288 234 
rect 285 234 288 237 
rect 285 237 288 240 
rect 285 240 288 243 
rect 285 243 288 246 
rect 285 246 288 249 
rect 285 249 288 252 
rect 285 252 288 255 
rect 285 255 288 258 
rect 285 258 288 261 
rect 285 261 288 264 
rect 285 264 288 267 
rect 285 267 288 270 
rect 285 270 288 273 
rect 285 273 288 276 
rect 285 276 288 279 
rect 285 279 288 282 
rect 285 282 288 285 
rect 285 285 288 288 
rect 285 288 288 291 
rect 285 291 288 294 
rect 285 294 288 297 
rect 285 297 288 300 
rect 285 300 288 303 
rect 285 303 288 306 
rect 285 306 288 309 
rect 285 309 288 312 
rect 285 312 288 315 
rect 285 315 288 318 
rect 285 318 288 321 
rect 285 321 288 324 
rect 285 324 288 327 
rect 285 327 288 330 
rect 285 330 288 333 
rect 285 333 288 336 
rect 285 336 288 339 
rect 285 339 288 342 
rect 285 342 288 345 
rect 285 345 288 348 
rect 285 348 288 351 
rect 285 351 288 354 
rect 285 354 288 357 
rect 285 357 288 360 
rect 285 360 288 363 
rect 285 363 288 366 
rect 285 366 288 369 
rect 285 369 288 372 
rect 285 372 288 375 
rect 285 375 288 378 
rect 285 378 288 381 
rect 285 381 288 384 
rect 285 384 288 387 
rect 285 387 288 390 
rect 285 390 288 393 
rect 285 393 288 396 
rect 285 396 288 399 
rect 285 399 288 402 
rect 285 402 288 405 
rect 285 405 288 408 
rect 285 408 288 411 
rect 285 411 288 414 
rect 285 414 288 417 
rect 285 417 288 420 
rect 285 420 288 423 
rect 285 423 288 426 
rect 285 426 288 429 
rect 285 429 288 432 
rect 285 432 288 435 
rect 285 435 288 438 
rect 285 438 288 441 
rect 285 441 288 444 
rect 285 444 288 447 
rect 285 447 288 450 
rect 285 450 288 453 
rect 285 453 288 456 
rect 285 456 288 459 
rect 285 459 288 462 
rect 285 462 288 465 
rect 285 465 288 468 
rect 285 468 288 471 
rect 285 471 288 474 
rect 285 474 288 477 
rect 285 477 288 480 
rect 285 480 288 483 
rect 285 483 288 486 
rect 285 486 288 489 
rect 285 489 288 492 
rect 285 492 288 495 
rect 285 495 288 498 
rect 285 498 288 501 
rect 285 501 288 504 
rect 285 504 288 507 
rect 285 507 288 510 
rect 288 0 291 3 
rect 288 3 291 6 
rect 288 6 291 9 
rect 288 9 291 12 
rect 288 12 291 15 
rect 288 15 291 18 
rect 288 18 291 21 
rect 288 21 291 24 
rect 288 24 291 27 
rect 288 27 291 30 
rect 288 30 291 33 
rect 288 33 291 36 
rect 288 36 291 39 
rect 288 39 291 42 
rect 288 42 291 45 
rect 288 45 291 48 
rect 288 48 291 51 
rect 288 51 291 54 
rect 288 54 291 57 
rect 288 57 291 60 
rect 288 60 291 63 
rect 288 63 291 66 
rect 288 66 291 69 
rect 288 69 291 72 
rect 288 72 291 75 
rect 288 75 291 78 
rect 288 78 291 81 
rect 288 81 291 84 
rect 288 84 291 87 
rect 288 87 291 90 
rect 288 90 291 93 
rect 288 93 291 96 
rect 288 96 291 99 
rect 288 99 291 102 
rect 288 102 291 105 
rect 288 105 291 108 
rect 288 108 291 111 
rect 288 111 291 114 
rect 288 114 291 117 
rect 288 117 291 120 
rect 288 120 291 123 
rect 288 123 291 126 
rect 288 126 291 129 
rect 288 129 291 132 
rect 288 132 291 135 
rect 288 135 291 138 
rect 288 138 291 141 
rect 288 141 291 144 
rect 288 144 291 147 
rect 288 147 291 150 
rect 288 150 291 153 
rect 288 153 291 156 
rect 288 156 291 159 
rect 288 159 291 162 
rect 288 162 291 165 
rect 288 165 291 168 
rect 288 168 291 171 
rect 288 171 291 174 
rect 288 174 291 177 
rect 288 177 291 180 
rect 288 180 291 183 
rect 288 183 291 186 
rect 288 186 291 189 
rect 288 189 291 192 
rect 288 192 291 195 
rect 288 195 291 198 
rect 288 198 291 201 
rect 288 201 291 204 
rect 288 204 291 207 
rect 288 207 291 210 
rect 288 210 291 213 
rect 288 213 291 216 
rect 288 216 291 219 
rect 288 219 291 222 
rect 288 222 291 225 
rect 288 225 291 228 
rect 288 228 291 231 
rect 288 231 291 234 
rect 288 234 291 237 
rect 288 237 291 240 
rect 288 240 291 243 
rect 288 243 291 246 
rect 288 246 291 249 
rect 288 249 291 252 
rect 288 252 291 255 
rect 288 255 291 258 
rect 288 258 291 261 
rect 288 261 291 264 
rect 288 264 291 267 
rect 288 267 291 270 
rect 288 270 291 273 
rect 288 273 291 276 
rect 288 276 291 279 
rect 288 279 291 282 
rect 288 282 291 285 
rect 288 285 291 288 
rect 288 288 291 291 
rect 288 291 291 294 
rect 288 294 291 297 
rect 288 297 291 300 
rect 288 300 291 303 
rect 288 303 291 306 
rect 288 306 291 309 
rect 288 309 291 312 
rect 288 312 291 315 
rect 288 315 291 318 
rect 288 318 291 321 
rect 288 321 291 324 
rect 288 324 291 327 
rect 288 327 291 330 
rect 288 330 291 333 
rect 288 333 291 336 
rect 288 336 291 339 
rect 288 339 291 342 
rect 288 342 291 345 
rect 288 345 291 348 
rect 288 348 291 351 
rect 288 351 291 354 
rect 288 354 291 357 
rect 288 357 291 360 
rect 288 360 291 363 
rect 288 363 291 366 
rect 288 366 291 369 
rect 288 369 291 372 
rect 288 372 291 375 
rect 288 375 291 378 
rect 288 378 291 381 
rect 288 381 291 384 
rect 288 384 291 387 
rect 288 387 291 390 
rect 288 390 291 393 
rect 288 393 291 396 
rect 288 396 291 399 
rect 288 399 291 402 
rect 288 402 291 405 
rect 288 405 291 408 
rect 288 408 291 411 
rect 288 411 291 414 
rect 288 414 291 417 
rect 288 417 291 420 
rect 288 420 291 423 
rect 288 423 291 426 
rect 288 426 291 429 
rect 288 429 291 432 
rect 288 432 291 435 
rect 288 435 291 438 
rect 288 438 291 441 
rect 288 441 291 444 
rect 288 444 291 447 
rect 288 447 291 450 
rect 288 450 291 453 
rect 288 453 291 456 
rect 288 456 291 459 
rect 288 459 291 462 
rect 288 462 291 465 
rect 288 465 291 468 
rect 288 468 291 471 
rect 288 471 291 474 
rect 288 474 291 477 
rect 288 477 291 480 
rect 288 480 291 483 
rect 288 483 291 486 
rect 288 486 291 489 
rect 288 489 291 492 
rect 288 492 291 495 
rect 288 495 291 498 
rect 288 498 291 501 
rect 288 501 291 504 
rect 288 504 291 507 
rect 288 507 291 510 
rect 291 0 294 3 
rect 291 3 294 6 
rect 291 6 294 9 
rect 291 9 294 12 
rect 291 12 294 15 
rect 291 15 294 18 
rect 291 18 294 21 
rect 291 21 294 24 
rect 291 24 294 27 
rect 291 27 294 30 
rect 291 30 294 33 
rect 291 33 294 36 
rect 291 36 294 39 
rect 291 39 294 42 
rect 291 42 294 45 
rect 291 45 294 48 
rect 291 48 294 51 
rect 291 51 294 54 
rect 291 54 294 57 
rect 291 57 294 60 
rect 291 60 294 63 
rect 291 63 294 66 
rect 291 66 294 69 
rect 291 69 294 72 
rect 291 72 294 75 
rect 291 75 294 78 
rect 291 78 294 81 
rect 291 81 294 84 
rect 291 84 294 87 
rect 291 87 294 90 
rect 291 90 294 93 
rect 291 93 294 96 
rect 291 96 294 99 
rect 291 99 294 102 
rect 291 102 294 105 
rect 291 105 294 108 
rect 291 108 294 111 
rect 291 111 294 114 
rect 291 114 294 117 
rect 291 117 294 120 
rect 291 120 294 123 
rect 291 123 294 126 
rect 291 126 294 129 
rect 291 129 294 132 
rect 291 132 294 135 
rect 291 135 294 138 
rect 291 138 294 141 
rect 291 141 294 144 
rect 291 144 294 147 
rect 291 147 294 150 
rect 291 150 294 153 
rect 291 153 294 156 
rect 291 156 294 159 
rect 291 159 294 162 
rect 291 162 294 165 
rect 291 165 294 168 
rect 291 168 294 171 
rect 291 171 294 174 
rect 291 174 294 177 
rect 291 177 294 180 
rect 291 180 294 183 
rect 291 183 294 186 
rect 291 186 294 189 
rect 291 189 294 192 
rect 291 192 294 195 
rect 291 195 294 198 
rect 291 198 294 201 
rect 291 201 294 204 
rect 291 204 294 207 
rect 291 207 294 210 
rect 291 210 294 213 
rect 291 213 294 216 
rect 291 216 294 219 
rect 291 219 294 222 
rect 291 222 294 225 
rect 291 225 294 228 
rect 291 228 294 231 
rect 291 231 294 234 
rect 291 234 294 237 
rect 291 237 294 240 
rect 291 240 294 243 
rect 291 243 294 246 
rect 291 246 294 249 
rect 291 249 294 252 
rect 291 252 294 255 
rect 291 255 294 258 
rect 291 258 294 261 
rect 291 261 294 264 
rect 291 264 294 267 
rect 291 267 294 270 
rect 291 270 294 273 
rect 291 273 294 276 
rect 291 276 294 279 
rect 291 279 294 282 
rect 291 282 294 285 
rect 291 285 294 288 
rect 291 288 294 291 
rect 291 291 294 294 
rect 291 294 294 297 
rect 291 297 294 300 
rect 291 300 294 303 
rect 291 303 294 306 
rect 291 306 294 309 
rect 291 309 294 312 
rect 291 312 294 315 
rect 291 315 294 318 
rect 291 318 294 321 
rect 291 321 294 324 
rect 291 324 294 327 
rect 291 327 294 330 
rect 291 330 294 333 
rect 291 333 294 336 
rect 291 336 294 339 
rect 291 339 294 342 
rect 291 342 294 345 
rect 291 345 294 348 
rect 291 348 294 351 
rect 291 351 294 354 
rect 291 354 294 357 
rect 291 357 294 360 
rect 291 360 294 363 
rect 291 363 294 366 
rect 291 366 294 369 
rect 291 369 294 372 
rect 291 372 294 375 
rect 291 375 294 378 
rect 291 378 294 381 
rect 291 381 294 384 
rect 291 384 294 387 
rect 291 387 294 390 
rect 291 390 294 393 
rect 291 393 294 396 
rect 291 396 294 399 
rect 291 399 294 402 
rect 291 402 294 405 
rect 291 405 294 408 
rect 291 408 294 411 
rect 291 411 294 414 
rect 291 414 294 417 
rect 291 417 294 420 
rect 291 420 294 423 
rect 291 423 294 426 
rect 291 426 294 429 
rect 291 429 294 432 
rect 291 432 294 435 
rect 291 435 294 438 
rect 291 438 294 441 
rect 291 441 294 444 
rect 291 444 294 447 
rect 291 447 294 450 
rect 291 450 294 453 
rect 291 453 294 456 
rect 291 456 294 459 
rect 291 459 294 462 
rect 291 462 294 465 
rect 291 465 294 468 
rect 291 468 294 471 
rect 291 471 294 474 
rect 291 474 294 477 
rect 291 477 294 480 
rect 291 480 294 483 
rect 291 483 294 486 
rect 291 486 294 489 
rect 291 489 294 492 
rect 291 492 294 495 
rect 291 495 294 498 
rect 291 498 294 501 
rect 291 501 294 504 
rect 291 504 294 507 
rect 291 507 294 510 
rect 294 0 297 3 
rect 294 3 297 6 
rect 294 6 297 9 
rect 294 9 297 12 
rect 294 12 297 15 
rect 294 15 297 18 
rect 294 18 297 21 
rect 294 21 297 24 
rect 294 24 297 27 
rect 294 27 297 30 
rect 294 30 297 33 
rect 294 33 297 36 
rect 294 36 297 39 
rect 294 39 297 42 
rect 294 42 297 45 
rect 294 45 297 48 
rect 294 48 297 51 
rect 294 51 297 54 
rect 294 54 297 57 
rect 294 57 297 60 
rect 294 60 297 63 
rect 294 63 297 66 
rect 294 66 297 69 
rect 294 69 297 72 
rect 294 72 297 75 
rect 294 75 297 78 
rect 294 78 297 81 
rect 294 81 297 84 
rect 294 84 297 87 
rect 294 87 297 90 
rect 294 90 297 93 
rect 294 93 297 96 
rect 294 96 297 99 
rect 294 99 297 102 
rect 294 102 297 105 
rect 294 105 297 108 
rect 294 108 297 111 
rect 294 111 297 114 
rect 294 114 297 117 
rect 294 117 297 120 
rect 294 120 297 123 
rect 294 123 297 126 
rect 294 126 297 129 
rect 294 129 297 132 
rect 294 132 297 135 
rect 294 135 297 138 
rect 294 138 297 141 
rect 294 141 297 144 
rect 294 144 297 147 
rect 294 147 297 150 
rect 294 150 297 153 
rect 294 153 297 156 
rect 294 156 297 159 
rect 294 159 297 162 
rect 294 162 297 165 
rect 294 165 297 168 
rect 294 168 297 171 
rect 294 171 297 174 
rect 294 174 297 177 
rect 294 177 297 180 
rect 294 180 297 183 
rect 294 183 297 186 
rect 294 186 297 189 
rect 294 189 297 192 
rect 294 192 297 195 
rect 294 195 297 198 
rect 294 198 297 201 
rect 294 201 297 204 
rect 294 204 297 207 
rect 294 207 297 210 
rect 294 210 297 213 
rect 294 213 297 216 
rect 294 216 297 219 
rect 294 219 297 222 
rect 294 222 297 225 
rect 294 225 297 228 
rect 294 228 297 231 
rect 294 231 297 234 
rect 294 234 297 237 
rect 294 237 297 240 
rect 294 240 297 243 
rect 294 243 297 246 
rect 294 246 297 249 
rect 294 249 297 252 
rect 294 252 297 255 
rect 294 255 297 258 
rect 294 258 297 261 
rect 294 261 297 264 
rect 294 264 297 267 
rect 294 267 297 270 
rect 294 270 297 273 
rect 294 273 297 276 
rect 294 276 297 279 
rect 294 279 297 282 
rect 294 282 297 285 
rect 294 285 297 288 
rect 294 288 297 291 
rect 294 291 297 294 
rect 294 294 297 297 
rect 294 297 297 300 
rect 294 300 297 303 
rect 294 303 297 306 
rect 294 306 297 309 
rect 294 309 297 312 
rect 294 312 297 315 
rect 294 315 297 318 
rect 294 318 297 321 
rect 294 321 297 324 
rect 294 324 297 327 
rect 294 327 297 330 
rect 294 330 297 333 
rect 294 333 297 336 
rect 294 336 297 339 
rect 294 339 297 342 
rect 294 342 297 345 
rect 294 345 297 348 
rect 294 348 297 351 
rect 294 351 297 354 
rect 294 354 297 357 
rect 294 357 297 360 
rect 294 360 297 363 
rect 294 363 297 366 
rect 294 366 297 369 
rect 294 369 297 372 
rect 294 372 297 375 
rect 294 375 297 378 
rect 294 378 297 381 
rect 294 381 297 384 
rect 294 384 297 387 
rect 294 387 297 390 
rect 294 390 297 393 
rect 294 393 297 396 
rect 294 396 297 399 
rect 294 399 297 402 
rect 294 402 297 405 
rect 294 405 297 408 
rect 294 408 297 411 
rect 294 411 297 414 
rect 294 414 297 417 
rect 294 417 297 420 
rect 294 420 297 423 
rect 294 423 297 426 
rect 294 426 297 429 
rect 294 429 297 432 
rect 294 432 297 435 
rect 294 435 297 438 
rect 294 438 297 441 
rect 294 441 297 444 
rect 294 444 297 447 
rect 294 447 297 450 
rect 294 450 297 453 
rect 294 453 297 456 
rect 294 456 297 459 
rect 294 459 297 462 
rect 294 462 297 465 
rect 294 465 297 468 
rect 294 468 297 471 
rect 294 471 297 474 
rect 294 474 297 477 
rect 294 477 297 480 
rect 294 480 297 483 
rect 294 483 297 486 
rect 294 486 297 489 
rect 294 489 297 492 
rect 294 492 297 495 
rect 294 495 297 498 
rect 294 498 297 501 
rect 294 501 297 504 
rect 294 504 297 507 
rect 294 507 297 510 
rect 297 0 300 3 
rect 297 3 300 6 
rect 297 6 300 9 
rect 297 9 300 12 
rect 297 12 300 15 
rect 297 15 300 18 
rect 297 18 300 21 
rect 297 21 300 24 
rect 297 24 300 27 
rect 297 27 300 30 
rect 297 30 300 33 
rect 297 33 300 36 
rect 297 36 300 39 
rect 297 39 300 42 
rect 297 42 300 45 
rect 297 45 300 48 
rect 297 48 300 51 
rect 297 51 300 54 
rect 297 54 300 57 
rect 297 57 300 60 
rect 297 60 300 63 
rect 297 63 300 66 
rect 297 66 300 69 
rect 297 69 300 72 
rect 297 72 300 75 
rect 297 75 300 78 
rect 297 78 300 81 
rect 297 81 300 84 
rect 297 84 300 87 
rect 297 87 300 90 
rect 297 90 300 93 
rect 297 93 300 96 
rect 297 96 300 99 
rect 297 99 300 102 
rect 297 102 300 105 
rect 297 105 300 108 
rect 297 108 300 111 
rect 297 111 300 114 
rect 297 114 300 117 
rect 297 117 300 120 
rect 297 120 300 123 
rect 297 123 300 126 
rect 297 126 300 129 
rect 297 129 300 132 
rect 297 132 300 135 
rect 297 135 300 138 
rect 297 138 300 141 
rect 297 141 300 144 
rect 297 144 300 147 
rect 297 147 300 150 
rect 297 150 300 153 
rect 297 153 300 156 
rect 297 156 300 159 
rect 297 159 300 162 
rect 297 162 300 165 
rect 297 165 300 168 
rect 297 168 300 171 
rect 297 171 300 174 
rect 297 174 300 177 
rect 297 177 300 180 
rect 297 180 300 183 
rect 297 183 300 186 
rect 297 186 300 189 
rect 297 189 300 192 
rect 297 192 300 195 
rect 297 195 300 198 
rect 297 198 300 201 
rect 297 201 300 204 
rect 297 204 300 207 
rect 297 207 300 210 
rect 297 210 300 213 
rect 297 213 300 216 
rect 297 216 300 219 
rect 297 219 300 222 
rect 297 222 300 225 
rect 297 225 300 228 
rect 297 228 300 231 
rect 297 231 300 234 
rect 297 234 300 237 
rect 297 237 300 240 
rect 297 240 300 243 
rect 297 243 300 246 
rect 297 246 300 249 
rect 297 249 300 252 
rect 297 252 300 255 
rect 297 255 300 258 
rect 297 258 300 261 
rect 297 261 300 264 
rect 297 264 300 267 
rect 297 267 300 270 
rect 297 270 300 273 
rect 297 273 300 276 
rect 297 276 300 279 
rect 297 279 300 282 
rect 297 282 300 285 
rect 297 285 300 288 
rect 297 288 300 291 
rect 297 291 300 294 
rect 297 294 300 297 
rect 297 297 300 300 
rect 297 300 300 303 
rect 297 303 300 306 
rect 297 306 300 309 
rect 297 309 300 312 
rect 297 312 300 315 
rect 297 315 300 318 
rect 297 318 300 321 
rect 297 321 300 324 
rect 297 324 300 327 
rect 297 327 300 330 
rect 297 330 300 333 
rect 297 333 300 336 
rect 297 336 300 339 
rect 297 339 300 342 
rect 297 342 300 345 
rect 297 345 300 348 
rect 297 348 300 351 
rect 297 351 300 354 
rect 297 354 300 357 
rect 297 357 300 360 
rect 297 360 300 363 
rect 297 363 300 366 
rect 297 366 300 369 
rect 297 369 300 372 
rect 297 372 300 375 
rect 297 375 300 378 
rect 297 378 300 381 
rect 297 381 300 384 
rect 297 384 300 387 
rect 297 387 300 390 
rect 297 390 300 393 
rect 297 393 300 396 
rect 297 396 300 399 
rect 297 399 300 402 
rect 297 402 300 405 
rect 297 405 300 408 
rect 297 408 300 411 
rect 297 411 300 414 
rect 297 414 300 417 
rect 297 417 300 420 
rect 297 420 300 423 
rect 297 423 300 426 
rect 297 426 300 429 
rect 297 429 300 432 
rect 297 432 300 435 
rect 297 435 300 438 
rect 297 438 300 441 
rect 297 441 300 444 
rect 297 444 300 447 
rect 297 447 300 450 
rect 297 450 300 453 
rect 297 453 300 456 
rect 297 456 300 459 
rect 297 459 300 462 
rect 297 462 300 465 
rect 297 465 300 468 
rect 297 468 300 471 
rect 297 471 300 474 
rect 297 474 300 477 
rect 297 477 300 480 
rect 297 480 300 483 
rect 297 483 300 486 
rect 297 486 300 489 
rect 297 489 300 492 
rect 297 492 300 495 
rect 297 495 300 498 
rect 297 498 300 501 
rect 297 501 300 504 
rect 297 504 300 507 
rect 297 507 300 510 
rect 300 0 303 3 
rect 300 3 303 6 
rect 300 6 303 9 
rect 300 9 303 12 
rect 300 12 303 15 
rect 300 15 303 18 
rect 300 18 303 21 
rect 300 21 303 24 
rect 300 24 303 27 
rect 300 27 303 30 
rect 300 30 303 33 
rect 300 33 303 36 
rect 300 36 303 39 
rect 300 39 303 42 
rect 300 42 303 45 
rect 300 45 303 48 
rect 300 48 303 51 
rect 300 51 303 54 
rect 300 54 303 57 
rect 300 57 303 60 
rect 300 60 303 63 
rect 300 63 303 66 
rect 300 66 303 69 
rect 300 69 303 72 
rect 300 72 303 75 
rect 300 75 303 78 
rect 300 78 303 81 
rect 300 81 303 84 
rect 300 84 303 87 
rect 300 87 303 90 
rect 300 90 303 93 
rect 300 93 303 96 
rect 300 96 303 99 
rect 300 99 303 102 
rect 300 102 303 105 
rect 300 105 303 108 
rect 300 108 303 111 
rect 300 111 303 114 
rect 300 114 303 117 
rect 300 117 303 120 
rect 300 120 303 123 
rect 300 123 303 126 
rect 300 126 303 129 
rect 300 129 303 132 
rect 300 132 303 135 
rect 300 135 303 138 
rect 300 138 303 141 
rect 300 141 303 144 
rect 300 144 303 147 
rect 300 147 303 150 
rect 300 150 303 153 
rect 300 153 303 156 
rect 300 156 303 159 
rect 300 159 303 162 
rect 300 162 303 165 
rect 300 165 303 168 
rect 300 168 303 171 
rect 300 171 303 174 
rect 300 174 303 177 
rect 300 177 303 180 
rect 300 180 303 183 
rect 300 183 303 186 
rect 300 186 303 189 
rect 300 189 303 192 
rect 300 192 303 195 
rect 300 195 303 198 
rect 300 198 303 201 
rect 300 201 303 204 
rect 300 204 303 207 
rect 300 207 303 210 
rect 300 210 303 213 
rect 300 213 303 216 
rect 300 216 303 219 
rect 300 219 303 222 
rect 300 222 303 225 
rect 300 225 303 228 
rect 300 228 303 231 
rect 300 231 303 234 
rect 300 234 303 237 
rect 300 237 303 240 
rect 300 240 303 243 
rect 300 243 303 246 
rect 300 246 303 249 
rect 300 249 303 252 
rect 300 252 303 255 
rect 300 255 303 258 
rect 300 258 303 261 
rect 300 261 303 264 
rect 300 264 303 267 
rect 300 267 303 270 
rect 300 270 303 273 
rect 300 273 303 276 
rect 300 276 303 279 
rect 300 279 303 282 
rect 300 282 303 285 
rect 300 285 303 288 
rect 300 288 303 291 
rect 300 291 303 294 
rect 300 294 303 297 
rect 300 297 303 300 
rect 300 300 303 303 
rect 300 303 303 306 
rect 300 306 303 309 
rect 300 309 303 312 
rect 300 312 303 315 
rect 300 315 303 318 
rect 300 318 303 321 
rect 300 321 303 324 
rect 300 324 303 327 
rect 300 327 303 330 
rect 300 330 303 333 
rect 300 333 303 336 
rect 300 336 303 339 
rect 300 339 303 342 
rect 300 342 303 345 
rect 300 345 303 348 
rect 300 348 303 351 
rect 300 351 303 354 
rect 300 354 303 357 
rect 300 357 303 360 
rect 300 360 303 363 
rect 300 363 303 366 
rect 300 366 303 369 
rect 300 369 303 372 
rect 300 372 303 375 
rect 300 375 303 378 
rect 300 378 303 381 
rect 300 381 303 384 
rect 300 384 303 387 
rect 300 387 303 390 
rect 300 390 303 393 
rect 300 393 303 396 
rect 300 396 303 399 
rect 300 399 303 402 
rect 300 402 303 405 
rect 300 405 303 408 
rect 300 408 303 411 
rect 300 411 303 414 
rect 300 414 303 417 
rect 300 417 303 420 
rect 300 420 303 423 
rect 300 423 303 426 
rect 300 426 303 429 
rect 300 429 303 432 
rect 300 432 303 435 
rect 300 435 303 438 
rect 300 438 303 441 
rect 300 441 303 444 
rect 300 444 303 447 
rect 300 447 303 450 
rect 300 450 303 453 
rect 300 453 303 456 
rect 300 456 303 459 
rect 300 459 303 462 
rect 300 462 303 465 
rect 300 465 303 468 
rect 300 468 303 471 
rect 300 471 303 474 
rect 300 474 303 477 
rect 300 477 303 480 
rect 300 480 303 483 
rect 300 483 303 486 
rect 300 486 303 489 
rect 300 489 303 492 
rect 300 492 303 495 
rect 300 495 303 498 
rect 300 498 303 501 
rect 300 501 303 504 
rect 300 504 303 507 
rect 300 507 303 510 
rect 303 0 306 3 
rect 303 3 306 6 
rect 303 6 306 9 
rect 303 9 306 12 
rect 303 12 306 15 
rect 303 15 306 18 
rect 303 18 306 21 
rect 303 21 306 24 
rect 303 24 306 27 
rect 303 27 306 30 
rect 303 30 306 33 
rect 303 33 306 36 
rect 303 36 306 39 
rect 303 39 306 42 
rect 303 42 306 45 
rect 303 45 306 48 
rect 303 48 306 51 
rect 303 51 306 54 
rect 303 54 306 57 
rect 303 57 306 60 
rect 303 60 306 63 
rect 303 63 306 66 
rect 303 66 306 69 
rect 303 69 306 72 
rect 303 72 306 75 
rect 303 75 306 78 
rect 303 78 306 81 
rect 303 81 306 84 
rect 303 84 306 87 
rect 303 87 306 90 
rect 303 90 306 93 
rect 303 93 306 96 
rect 303 96 306 99 
rect 303 99 306 102 
rect 303 102 306 105 
rect 303 105 306 108 
rect 303 108 306 111 
rect 303 111 306 114 
rect 303 114 306 117 
rect 303 117 306 120 
rect 303 120 306 123 
rect 303 123 306 126 
rect 303 126 306 129 
rect 303 129 306 132 
rect 303 132 306 135 
rect 303 135 306 138 
rect 303 138 306 141 
rect 303 141 306 144 
rect 303 144 306 147 
rect 303 147 306 150 
rect 303 150 306 153 
rect 303 153 306 156 
rect 303 156 306 159 
rect 303 159 306 162 
rect 303 162 306 165 
rect 303 165 306 168 
rect 303 168 306 171 
rect 303 171 306 174 
rect 303 174 306 177 
rect 303 177 306 180 
rect 303 180 306 183 
rect 303 183 306 186 
rect 303 186 306 189 
rect 303 189 306 192 
rect 303 192 306 195 
rect 303 195 306 198 
rect 303 198 306 201 
rect 303 201 306 204 
rect 303 204 306 207 
rect 303 207 306 210 
rect 303 210 306 213 
rect 303 213 306 216 
rect 303 216 306 219 
rect 303 219 306 222 
rect 303 222 306 225 
rect 303 225 306 228 
rect 303 228 306 231 
rect 303 231 306 234 
rect 303 234 306 237 
rect 303 237 306 240 
rect 303 240 306 243 
rect 303 243 306 246 
rect 303 246 306 249 
rect 303 249 306 252 
rect 303 252 306 255 
rect 303 255 306 258 
rect 303 258 306 261 
rect 303 261 306 264 
rect 303 264 306 267 
rect 303 267 306 270 
rect 303 270 306 273 
rect 303 273 306 276 
rect 303 276 306 279 
rect 303 279 306 282 
rect 303 282 306 285 
rect 303 285 306 288 
rect 303 288 306 291 
rect 303 291 306 294 
rect 303 294 306 297 
rect 303 297 306 300 
rect 303 300 306 303 
rect 303 303 306 306 
rect 303 306 306 309 
rect 303 309 306 312 
rect 303 312 306 315 
rect 303 315 306 318 
rect 303 318 306 321 
rect 303 321 306 324 
rect 303 324 306 327 
rect 303 327 306 330 
rect 303 330 306 333 
rect 303 333 306 336 
rect 303 336 306 339 
rect 303 339 306 342 
rect 303 342 306 345 
rect 303 345 306 348 
rect 303 348 306 351 
rect 303 351 306 354 
rect 303 354 306 357 
rect 303 357 306 360 
rect 303 360 306 363 
rect 303 363 306 366 
rect 303 366 306 369 
rect 303 369 306 372 
rect 303 372 306 375 
rect 303 375 306 378 
rect 303 378 306 381 
rect 303 381 306 384 
rect 303 384 306 387 
rect 303 387 306 390 
rect 303 390 306 393 
rect 303 393 306 396 
rect 303 396 306 399 
rect 303 399 306 402 
rect 303 402 306 405 
rect 303 405 306 408 
rect 303 408 306 411 
rect 303 411 306 414 
rect 303 414 306 417 
rect 303 417 306 420 
rect 303 420 306 423 
rect 303 423 306 426 
rect 303 426 306 429 
rect 303 429 306 432 
rect 303 432 306 435 
rect 303 435 306 438 
rect 303 438 306 441 
rect 303 441 306 444 
rect 303 444 306 447 
rect 303 447 306 450 
rect 303 450 306 453 
rect 303 453 306 456 
rect 303 456 306 459 
rect 303 459 306 462 
rect 303 462 306 465 
rect 303 465 306 468 
rect 303 468 306 471 
rect 303 471 306 474 
rect 303 474 306 477 
rect 303 477 306 480 
rect 303 480 306 483 
rect 303 483 306 486 
rect 303 486 306 489 
rect 303 489 306 492 
rect 303 492 306 495 
rect 303 495 306 498 
rect 303 498 306 501 
rect 303 501 306 504 
rect 303 504 306 507 
rect 303 507 306 510 
rect 306 0 309 3 
rect 306 3 309 6 
rect 306 6 309 9 
rect 306 9 309 12 
rect 306 12 309 15 
rect 306 15 309 18 
rect 306 18 309 21 
rect 306 21 309 24 
rect 306 24 309 27 
rect 306 27 309 30 
rect 306 30 309 33 
rect 306 33 309 36 
rect 306 36 309 39 
rect 306 39 309 42 
rect 306 42 309 45 
rect 306 45 309 48 
rect 306 48 309 51 
rect 306 51 309 54 
rect 306 54 309 57 
rect 306 57 309 60 
rect 306 60 309 63 
rect 306 63 309 66 
rect 306 66 309 69 
rect 306 69 309 72 
rect 306 72 309 75 
rect 306 75 309 78 
rect 306 78 309 81 
rect 306 81 309 84 
rect 306 84 309 87 
rect 306 87 309 90 
rect 306 90 309 93 
rect 306 93 309 96 
rect 306 96 309 99 
rect 306 99 309 102 
rect 306 102 309 105 
rect 306 105 309 108 
rect 306 108 309 111 
rect 306 111 309 114 
rect 306 114 309 117 
rect 306 117 309 120 
rect 306 120 309 123 
rect 306 123 309 126 
rect 306 126 309 129 
rect 306 129 309 132 
rect 306 132 309 135 
rect 306 135 309 138 
rect 306 138 309 141 
rect 306 141 309 144 
rect 306 144 309 147 
rect 306 147 309 150 
rect 306 150 309 153 
rect 306 153 309 156 
rect 306 156 309 159 
rect 306 159 309 162 
rect 306 162 309 165 
rect 306 165 309 168 
rect 306 168 309 171 
rect 306 171 309 174 
rect 306 174 309 177 
rect 306 177 309 180 
rect 306 180 309 183 
rect 306 183 309 186 
rect 306 186 309 189 
rect 306 189 309 192 
rect 306 192 309 195 
rect 306 195 309 198 
rect 306 198 309 201 
rect 306 201 309 204 
rect 306 204 309 207 
rect 306 207 309 210 
rect 306 210 309 213 
rect 306 213 309 216 
rect 306 216 309 219 
rect 306 219 309 222 
rect 306 222 309 225 
rect 306 225 309 228 
rect 306 228 309 231 
rect 306 231 309 234 
rect 306 234 309 237 
rect 306 237 309 240 
rect 306 240 309 243 
rect 306 243 309 246 
rect 306 246 309 249 
rect 306 249 309 252 
rect 306 252 309 255 
rect 306 255 309 258 
rect 306 258 309 261 
rect 306 261 309 264 
rect 306 264 309 267 
rect 306 267 309 270 
rect 306 270 309 273 
rect 306 273 309 276 
rect 306 276 309 279 
rect 306 279 309 282 
rect 306 282 309 285 
rect 306 285 309 288 
rect 306 288 309 291 
rect 306 291 309 294 
rect 306 294 309 297 
rect 306 297 309 300 
rect 306 300 309 303 
rect 306 303 309 306 
rect 306 306 309 309 
rect 306 309 309 312 
rect 306 312 309 315 
rect 306 315 309 318 
rect 306 318 309 321 
rect 306 321 309 324 
rect 306 324 309 327 
rect 306 327 309 330 
rect 306 330 309 333 
rect 306 333 309 336 
rect 306 336 309 339 
rect 306 339 309 342 
rect 306 342 309 345 
rect 306 345 309 348 
rect 306 348 309 351 
rect 306 351 309 354 
rect 306 354 309 357 
rect 306 357 309 360 
rect 306 360 309 363 
rect 306 363 309 366 
rect 306 366 309 369 
rect 306 369 309 372 
rect 306 372 309 375 
rect 306 375 309 378 
rect 306 378 309 381 
rect 306 381 309 384 
rect 306 384 309 387 
rect 306 387 309 390 
rect 306 390 309 393 
rect 306 393 309 396 
rect 306 396 309 399 
rect 306 399 309 402 
rect 306 402 309 405 
rect 306 405 309 408 
rect 306 408 309 411 
rect 306 411 309 414 
rect 306 414 309 417 
rect 306 417 309 420 
rect 306 420 309 423 
rect 306 423 309 426 
rect 306 426 309 429 
rect 306 429 309 432 
rect 306 432 309 435 
rect 306 435 309 438 
rect 306 438 309 441 
rect 306 441 309 444 
rect 306 444 309 447 
rect 306 447 309 450 
rect 306 450 309 453 
rect 306 453 309 456 
rect 306 456 309 459 
rect 306 459 309 462 
rect 306 462 309 465 
rect 306 465 309 468 
rect 306 468 309 471 
rect 306 471 309 474 
rect 306 474 309 477 
rect 306 477 309 480 
rect 306 480 309 483 
rect 306 483 309 486 
rect 306 486 309 489 
rect 306 489 309 492 
rect 306 492 309 495 
rect 306 495 309 498 
rect 306 498 309 501 
rect 306 501 309 504 
rect 306 504 309 507 
rect 306 507 309 510 
rect 309 0 312 3 
rect 309 3 312 6 
rect 309 6 312 9 
rect 309 9 312 12 
rect 309 12 312 15 
rect 309 15 312 18 
rect 309 18 312 21 
rect 309 21 312 24 
rect 309 24 312 27 
rect 309 27 312 30 
rect 309 30 312 33 
rect 309 33 312 36 
rect 309 36 312 39 
rect 309 39 312 42 
rect 309 42 312 45 
rect 309 45 312 48 
rect 309 48 312 51 
rect 309 51 312 54 
rect 309 54 312 57 
rect 309 57 312 60 
rect 309 60 312 63 
rect 309 63 312 66 
rect 309 66 312 69 
rect 309 69 312 72 
rect 309 72 312 75 
rect 309 75 312 78 
rect 309 78 312 81 
rect 309 81 312 84 
rect 309 84 312 87 
rect 309 87 312 90 
rect 309 90 312 93 
rect 309 93 312 96 
rect 309 96 312 99 
rect 309 99 312 102 
rect 309 102 312 105 
rect 309 105 312 108 
rect 309 108 312 111 
rect 309 111 312 114 
rect 309 114 312 117 
rect 309 117 312 120 
rect 309 120 312 123 
rect 309 123 312 126 
rect 309 126 312 129 
rect 309 129 312 132 
rect 309 132 312 135 
rect 309 135 312 138 
rect 309 138 312 141 
rect 309 141 312 144 
rect 309 144 312 147 
rect 309 147 312 150 
rect 309 150 312 153 
rect 309 153 312 156 
rect 309 156 312 159 
rect 309 159 312 162 
rect 309 162 312 165 
rect 309 165 312 168 
rect 309 168 312 171 
rect 309 171 312 174 
rect 309 174 312 177 
rect 309 177 312 180 
rect 309 180 312 183 
rect 309 183 312 186 
rect 309 186 312 189 
rect 309 189 312 192 
rect 309 192 312 195 
rect 309 195 312 198 
rect 309 198 312 201 
rect 309 201 312 204 
rect 309 204 312 207 
rect 309 207 312 210 
rect 309 210 312 213 
rect 309 213 312 216 
rect 309 216 312 219 
rect 309 219 312 222 
rect 309 222 312 225 
rect 309 225 312 228 
rect 309 228 312 231 
rect 309 231 312 234 
rect 309 234 312 237 
rect 309 237 312 240 
rect 309 240 312 243 
rect 309 243 312 246 
rect 309 246 312 249 
rect 309 249 312 252 
rect 309 252 312 255 
rect 309 255 312 258 
rect 309 258 312 261 
rect 309 261 312 264 
rect 309 264 312 267 
rect 309 267 312 270 
rect 309 270 312 273 
rect 309 273 312 276 
rect 309 276 312 279 
rect 309 279 312 282 
rect 309 282 312 285 
rect 309 285 312 288 
rect 309 288 312 291 
rect 309 291 312 294 
rect 309 294 312 297 
rect 309 297 312 300 
rect 309 300 312 303 
rect 309 303 312 306 
rect 309 306 312 309 
rect 309 309 312 312 
rect 309 312 312 315 
rect 309 315 312 318 
rect 309 318 312 321 
rect 309 321 312 324 
rect 309 324 312 327 
rect 309 327 312 330 
rect 309 330 312 333 
rect 309 333 312 336 
rect 309 336 312 339 
rect 309 339 312 342 
rect 309 342 312 345 
rect 309 345 312 348 
rect 309 348 312 351 
rect 309 351 312 354 
rect 309 354 312 357 
rect 309 357 312 360 
rect 309 360 312 363 
rect 309 363 312 366 
rect 309 366 312 369 
rect 309 369 312 372 
rect 309 372 312 375 
rect 309 375 312 378 
rect 309 378 312 381 
rect 309 381 312 384 
rect 309 384 312 387 
rect 309 387 312 390 
rect 309 390 312 393 
rect 309 393 312 396 
rect 309 396 312 399 
rect 309 399 312 402 
rect 309 402 312 405 
rect 309 405 312 408 
rect 309 408 312 411 
rect 309 411 312 414 
rect 309 414 312 417 
rect 309 417 312 420 
rect 309 420 312 423 
rect 309 423 312 426 
rect 309 426 312 429 
rect 309 429 312 432 
rect 309 432 312 435 
rect 309 435 312 438 
rect 309 438 312 441 
rect 309 441 312 444 
rect 309 444 312 447 
rect 309 447 312 450 
rect 309 450 312 453 
rect 309 453 312 456 
rect 309 456 312 459 
rect 309 459 312 462 
rect 309 462 312 465 
rect 309 465 312 468 
rect 309 468 312 471 
rect 309 471 312 474 
rect 309 474 312 477 
rect 309 477 312 480 
rect 309 480 312 483 
rect 309 483 312 486 
rect 309 486 312 489 
rect 309 489 312 492 
rect 309 492 312 495 
rect 309 495 312 498 
rect 309 498 312 501 
rect 309 501 312 504 
rect 309 504 312 507 
rect 309 507 312 510 
rect 312 0 315 3 
rect 312 3 315 6 
rect 312 6 315 9 
rect 312 9 315 12 
rect 312 12 315 15 
rect 312 15 315 18 
rect 312 18 315 21 
rect 312 21 315 24 
rect 312 24 315 27 
rect 312 27 315 30 
rect 312 30 315 33 
rect 312 33 315 36 
rect 312 36 315 39 
rect 312 39 315 42 
rect 312 42 315 45 
rect 312 45 315 48 
rect 312 48 315 51 
rect 312 51 315 54 
rect 312 54 315 57 
rect 312 57 315 60 
rect 312 60 315 63 
rect 312 63 315 66 
rect 312 66 315 69 
rect 312 69 315 72 
rect 312 72 315 75 
rect 312 75 315 78 
rect 312 78 315 81 
rect 312 81 315 84 
rect 312 84 315 87 
rect 312 87 315 90 
rect 312 90 315 93 
rect 312 93 315 96 
rect 312 96 315 99 
rect 312 99 315 102 
rect 312 102 315 105 
rect 312 105 315 108 
rect 312 108 315 111 
rect 312 111 315 114 
rect 312 114 315 117 
rect 312 117 315 120 
rect 312 120 315 123 
rect 312 123 315 126 
rect 312 126 315 129 
rect 312 129 315 132 
rect 312 132 315 135 
rect 312 135 315 138 
rect 312 138 315 141 
rect 312 141 315 144 
rect 312 144 315 147 
rect 312 147 315 150 
rect 312 150 315 153 
rect 312 153 315 156 
rect 312 156 315 159 
rect 312 159 315 162 
rect 312 162 315 165 
rect 312 165 315 168 
rect 312 168 315 171 
rect 312 171 315 174 
rect 312 174 315 177 
rect 312 177 315 180 
rect 312 180 315 183 
rect 312 183 315 186 
rect 312 186 315 189 
rect 312 189 315 192 
rect 312 192 315 195 
rect 312 195 315 198 
rect 312 198 315 201 
rect 312 201 315 204 
rect 312 204 315 207 
rect 312 207 315 210 
rect 312 210 315 213 
rect 312 213 315 216 
rect 312 216 315 219 
rect 312 219 315 222 
rect 312 222 315 225 
rect 312 225 315 228 
rect 312 228 315 231 
rect 312 231 315 234 
rect 312 234 315 237 
rect 312 237 315 240 
rect 312 240 315 243 
rect 312 243 315 246 
rect 312 246 315 249 
rect 312 249 315 252 
rect 312 252 315 255 
rect 312 255 315 258 
rect 312 258 315 261 
rect 312 261 315 264 
rect 312 264 315 267 
rect 312 267 315 270 
rect 312 270 315 273 
rect 312 273 315 276 
rect 312 276 315 279 
rect 312 279 315 282 
rect 312 282 315 285 
rect 312 285 315 288 
rect 312 288 315 291 
rect 312 291 315 294 
rect 312 294 315 297 
rect 312 297 315 300 
rect 312 300 315 303 
rect 312 303 315 306 
rect 312 306 315 309 
rect 312 309 315 312 
rect 312 312 315 315 
rect 312 315 315 318 
rect 312 318 315 321 
rect 312 321 315 324 
rect 312 324 315 327 
rect 312 327 315 330 
rect 312 330 315 333 
rect 312 333 315 336 
rect 312 336 315 339 
rect 312 339 315 342 
rect 312 342 315 345 
rect 312 345 315 348 
rect 312 348 315 351 
rect 312 351 315 354 
rect 312 354 315 357 
rect 312 357 315 360 
rect 312 360 315 363 
rect 312 363 315 366 
rect 312 366 315 369 
rect 312 369 315 372 
rect 312 372 315 375 
rect 312 375 315 378 
rect 312 378 315 381 
rect 312 381 315 384 
rect 312 384 315 387 
rect 312 387 315 390 
rect 312 390 315 393 
rect 312 393 315 396 
rect 312 396 315 399 
rect 312 399 315 402 
rect 312 402 315 405 
rect 312 405 315 408 
rect 312 408 315 411 
rect 312 411 315 414 
rect 312 414 315 417 
rect 312 417 315 420 
rect 312 420 315 423 
rect 312 423 315 426 
rect 312 426 315 429 
rect 312 429 315 432 
rect 312 432 315 435 
rect 312 435 315 438 
rect 312 438 315 441 
rect 312 441 315 444 
rect 312 444 315 447 
rect 312 447 315 450 
rect 312 450 315 453 
rect 312 453 315 456 
rect 312 456 315 459 
rect 312 459 315 462 
rect 312 462 315 465 
rect 312 465 315 468 
rect 312 468 315 471 
rect 312 471 315 474 
rect 312 474 315 477 
rect 312 477 315 480 
rect 312 480 315 483 
rect 312 483 315 486 
rect 312 486 315 489 
rect 312 489 315 492 
rect 312 492 315 495 
rect 312 495 315 498 
rect 312 498 315 501 
rect 312 501 315 504 
rect 312 504 315 507 
rect 312 507 315 510 
rect 315 0 318 3 
rect 315 3 318 6 
rect 315 6 318 9 
rect 315 9 318 12 
rect 315 12 318 15 
rect 315 15 318 18 
rect 315 18 318 21 
rect 315 21 318 24 
rect 315 24 318 27 
rect 315 27 318 30 
rect 315 30 318 33 
rect 315 33 318 36 
rect 315 36 318 39 
rect 315 39 318 42 
rect 315 42 318 45 
rect 315 45 318 48 
rect 315 48 318 51 
rect 315 51 318 54 
rect 315 54 318 57 
rect 315 57 318 60 
rect 315 60 318 63 
rect 315 63 318 66 
rect 315 66 318 69 
rect 315 69 318 72 
rect 315 72 318 75 
rect 315 75 318 78 
rect 315 78 318 81 
rect 315 81 318 84 
rect 315 84 318 87 
rect 315 87 318 90 
rect 315 90 318 93 
rect 315 93 318 96 
rect 315 96 318 99 
rect 315 99 318 102 
rect 315 102 318 105 
rect 315 105 318 108 
rect 315 108 318 111 
rect 315 111 318 114 
rect 315 114 318 117 
rect 315 117 318 120 
rect 315 120 318 123 
rect 315 123 318 126 
rect 315 126 318 129 
rect 315 129 318 132 
rect 315 132 318 135 
rect 315 135 318 138 
rect 315 138 318 141 
rect 315 141 318 144 
rect 315 144 318 147 
rect 315 147 318 150 
rect 315 150 318 153 
rect 315 153 318 156 
rect 315 156 318 159 
rect 315 159 318 162 
rect 315 162 318 165 
rect 315 165 318 168 
rect 315 168 318 171 
rect 315 171 318 174 
rect 315 174 318 177 
rect 315 177 318 180 
rect 315 180 318 183 
rect 315 183 318 186 
rect 315 186 318 189 
rect 315 189 318 192 
rect 315 192 318 195 
rect 315 195 318 198 
rect 315 198 318 201 
rect 315 201 318 204 
rect 315 204 318 207 
rect 315 207 318 210 
rect 315 210 318 213 
rect 315 213 318 216 
rect 315 216 318 219 
rect 315 219 318 222 
rect 315 222 318 225 
rect 315 225 318 228 
rect 315 228 318 231 
rect 315 231 318 234 
rect 315 234 318 237 
rect 315 237 318 240 
rect 315 240 318 243 
rect 315 243 318 246 
rect 315 246 318 249 
rect 315 249 318 252 
rect 315 252 318 255 
rect 315 255 318 258 
rect 315 258 318 261 
rect 315 261 318 264 
rect 315 264 318 267 
rect 315 267 318 270 
rect 315 270 318 273 
rect 315 273 318 276 
rect 315 276 318 279 
rect 315 279 318 282 
rect 315 282 318 285 
rect 315 285 318 288 
rect 315 288 318 291 
rect 315 291 318 294 
rect 315 294 318 297 
rect 315 297 318 300 
rect 315 300 318 303 
rect 315 303 318 306 
rect 315 306 318 309 
rect 315 309 318 312 
rect 315 312 318 315 
rect 315 315 318 318 
rect 315 318 318 321 
rect 315 321 318 324 
rect 315 324 318 327 
rect 315 327 318 330 
rect 315 330 318 333 
rect 315 333 318 336 
rect 315 336 318 339 
rect 315 339 318 342 
rect 315 342 318 345 
rect 315 345 318 348 
rect 315 348 318 351 
rect 315 351 318 354 
rect 315 354 318 357 
rect 315 357 318 360 
rect 315 360 318 363 
rect 315 363 318 366 
rect 315 366 318 369 
rect 315 369 318 372 
rect 315 372 318 375 
rect 315 375 318 378 
rect 315 378 318 381 
rect 315 381 318 384 
rect 315 384 318 387 
rect 315 387 318 390 
rect 315 390 318 393 
rect 315 393 318 396 
rect 315 396 318 399 
rect 315 399 318 402 
rect 315 402 318 405 
rect 315 405 318 408 
rect 315 408 318 411 
rect 315 411 318 414 
rect 315 414 318 417 
rect 315 417 318 420 
rect 315 420 318 423 
rect 315 423 318 426 
rect 315 426 318 429 
rect 315 429 318 432 
rect 315 432 318 435 
rect 315 435 318 438 
rect 315 438 318 441 
rect 315 441 318 444 
rect 315 444 318 447 
rect 315 447 318 450 
rect 315 450 318 453 
rect 315 453 318 456 
rect 315 456 318 459 
rect 315 459 318 462 
rect 315 462 318 465 
rect 315 465 318 468 
rect 315 468 318 471 
rect 315 471 318 474 
rect 315 474 318 477 
rect 315 477 318 480 
rect 315 480 318 483 
rect 315 483 318 486 
rect 315 486 318 489 
rect 315 489 318 492 
rect 315 492 318 495 
rect 315 495 318 498 
rect 315 498 318 501 
rect 315 501 318 504 
rect 315 504 318 507 
rect 315 507 318 510 
rect 318 0 321 3 
rect 318 3 321 6 
rect 318 6 321 9 
rect 318 9 321 12 
rect 318 12 321 15 
rect 318 15 321 18 
rect 318 18 321 21 
rect 318 21 321 24 
rect 318 24 321 27 
rect 318 27 321 30 
rect 318 30 321 33 
rect 318 33 321 36 
rect 318 36 321 39 
rect 318 39 321 42 
rect 318 42 321 45 
rect 318 45 321 48 
rect 318 48 321 51 
rect 318 51 321 54 
rect 318 54 321 57 
rect 318 57 321 60 
rect 318 60 321 63 
rect 318 63 321 66 
rect 318 66 321 69 
rect 318 69 321 72 
rect 318 72 321 75 
rect 318 75 321 78 
rect 318 78 321 81 
rect 318 81 321 84 
rect 318 84 321 87 
rect 318 87 321 90 
rect 318 90 321 93 
rect 318 93 321 96 
rect 318 96 321 99 
rect 318 99 321 102 
rect 318 102 321 105 
rect 318 105 321 108 
rect 318 108 321 111 
rect 318 111 321 114 
rect 318 114 321 117 
rect 318 117 321 120 
rect 318 120 321 123 
rect 318 123 321 126 
rect 318 126 321 129 
rect 318 129 321 132 
rect 318 132 321 135 
rect 318 135 321 138 
rect 318 138 321 141 
rect 318 141 321 144 
rect 318 144 321 147 
rect 318 147 321 150 
rect 318 150 321 153 
rect 318 153 321 156 
rect 318 156 321 159 
rect 318 159 321 162 
rect 318 162 321 165 
rect 318 165 321 168 
rect 318 168 321 171 
rect 318 171 321 174 
rect 318 174 321 177 
rect 318 177 321 180 
rect 318 180 321 183 
rect 318 183 321 186 
rect 318 186 321 189 
rect 318 189 321 192 
rect 318 192 321 195 
rect 318 195 321 198 
rect 318 198 321 201 
rect 318 201 321 204 
rect 318 204 321 207 
rect 318 207 321 210 
rect 318 210 321 213 
rect 318 213 321 216 
rect 318 216 321 219 
rect 318 219 321 222 
rect 318 222 321 225 
rect 318 225 321 228 
rect 318 228 321 231 
rect 318 231 321 234 
rect 318 234 321 237 
rect 318 237 321 240 
rect 318 240 321 243 
rect 318 243 321 246 
rect 318 246 321 249 
rect 318 249 321 252 
rect 318 252 321 255 
rect 318 255 321 258 
rect 318 258 321 261 
rect 318 261 321 264 
rect 318 264 321 267 
rect 318 267 321 270 
rect 318 270 321 273 
rect 318 273 321 276 
rect 318 276 321 279 
rect 318 279 321 282 
rect 318 282 321 285 
rect 318 285 321 288 
rect 318 288 321 291 
rect 318 291 321 294 
rect 318 294 321 297 
rect 318 297 321 300 
rect 318 300 321 303 
rect 318 303 321 306 
rect 318 306 321 309 
rect 318 309 321 312 
rect 318 312 321 315 
rect 318 315 321 318 
rect 318 318 321 321 
rect 318 321 321 324 
rect 318 324 321 327 
rect 318 327 321 330 
rect 318 330 321 333 
rect 318 333 321 336 
rect 318 336 321 339 
rect 318 339 321 342 
rect 318 342 321 345 
rect 318 345 321 348 
rect 318 348 321 351 
rect 318 351 321 354 
rect 318 354 321 357 
rect 318 357 321 360 
rect 318 360 321 363 
rect 318 363 321 366 
rect 318 366 321 369 
rect 318 369 321 372 
rect 318 372 321 375 
rect 318 375 321 378 
rect 318 378 321 381 
rect 318 381 321 384 
rect 318 384 321 387 
rect 318 387 321 390 
rect 318 390 321 393 
rect 318 393 321 396 
rect 318 396 321 399 
rect 318 399 321 402 
rect 318 402 321 405 
rect 318 405 321 408 
rect 318 408 321 411 
rect 318 411 321 414 
rect 318 414 321 417 
rect 318 417 321 420 
rect 318 420 321 423 
rect 318 423 321 426 
rect 318 426 321 429 
rect 318 429 321 432 
rect 318 432 321 435 
rect 318 435 321 438 
rect 318 438 321 441 
rect 318 441 321 444 
rect 318 444 321 447 
rect 318 447 321 450 
rect 318 450 321 453 
rect 318 453 321 456 
rect 318 456 321 459 
rect 318 459 321 462 
rect 318 462 321 465 
rect 318 465 321 468 
rect 318 468 321 471 
rect 318 471 321 474 
rect 318 474 321 477 
rect 318 477 321 480 
rect 318 480 321 483 
rect 318 483 321 486 
rect 318 486 321 489 
rect 318 489 321 492 
rect 318 492 321 495 
rect 318 495 321 498 
rect 318 498 321 501 
rect 318 501 321 504 
rect 318 504 321 507 
rect 318 507 321 510 
rect 321 0 324 3 
rect 321 3 324 6 
rect 321 6 324 9 
rect 321 9 324 12 
rect 321 12 324 15 
rect 321 15 324 18 
rect 321 18 324 21 
rect 321 21 324 24 
rect 321 24 324 27 
rect 321 27 324 30 
rect 321 30 324 33 
rect 321 33 324 36 
rect 321 36 324 39 
rect 321 39 324 42 
rect 321 42 324 45 
rect 321 45 324 48 
rect 321 48 324 51 
rect 321 51 324 54 
rect 321 54 324 57 
rect 321 57 324 60 
rect 321 60 324 63 
rect 321 63 324 66 
rect 321 66 324 69 
rect 321 69 324 72 
rect 321 72 324 75 
rect 321 75 324 78 
rect 321 78 324 81 
rect 321 81 324 84 
rect 321 84 324 87 
rect 321 87 324 90 
rect 321 90 324 93 
rect 321 93 324 96 
rect 321 96 324 99 
rect 321 99 324 102 
rect 321 102 324 105 
rect 321 105 324 108 
rect 321 108 324 111 
rect 321 111 324 114 
rect 321 114 324 117 
rect 321 117 324 120 
rect 321 120 324 123 
rect 321 123 324 126 
rect 321 126 324 129 
rect 321 129 324 132 
rect 321 132 324 135 
rect 321 135 324 138 
rect 321 138 324 141 
rect 321 141 324 144 
rect 321 144 324 147 
rect 321 147 324 150 
rect 321 150 324 153 
rect 321 153 324 156 
rect 321 156 324 159 
rect 321 159 324 162 
rect 321 162 324 165 
rect 321 165 324 168 
rect 321 168 324 171 
rect 321 171 324 174 
rect 321 174 324 177 
rect 321 177 324 180 
rect 321 180 324 183 
rect 321 183 324 186 
rect 321 186 324 189 
rect 321 189 324 192 
rect 321 192 324 195 
rect 321 195 324 198 
rect 321 198 324 201 
rect 321 201 324 204 
rect 321 204 324 207 
rect 321 207 324 210 
rect 321 210 324 213 
rect 321 213 324 216 
rect 321 216 324 219 
rect 321 219 324 222 
rect 321 222 324 225 
rect 321 225 324 228 
rect 321 228 324 231 
rect 321 231 324 234 
rect 321 234 324 237 
rect 321 237 324 240 
rect 321 240 324 243 
rect 321 243 324 246 
rect 321 246 324 249 
rect 321 249 324 252 
rect 321 252 324 255 
rect 321 255 324 258 
rect 321 258 324 261 
rect 321 261 324 264 
rect 321 264 324 267 
rect 321 267 324 270 
rect 321 270 324 273 
rect 321 273 324 276 
rect 321 276 324 279 
rect 321 279 324 282 
rect 321 282 324 285 
rect 321 285 324 288 
rect 321 288 324 291 
rect 321 291 324 294 
rect 321 294 324 297 
rect 321 297 324 300 
rect 321 300 324 303 
rect 321 303 324 306 
rect 321 306 324 309 
rect 321 309 324 312 
rect 321 312 324 315 
rect 321 315 324 318 
rect 321 318 324 321 
rect 321 321 324 324 
rect 321 324 324 327 
rect 321 327 324 330 
rect 321 330 324 333 
rect 321 333 324 336 
rect 321 336 324 339 
rect 321 339 324 342 
rect 321 342 324 345 
rect 321 345 324 348 
rect 321 348 324 351 
rect 321 351 324 354 
rect 321 354 324 357 
rect 321 357 324 360 
rect 321 360 324 363 
rect 321 363 324 366 
rect 321 366 324 369 
rect 321 369 324 372 
rect 321 372 324 375 
rect 321 375 324 378 
rect 321 378 324 381 
rect 321 381 324 384 
rect 321 384 324 387 
rect 321 387 324 390 
rect 321 390 324 393 
rect 321 393 324 396 
rect 321 396 324 399 
rect 321 399 324 402 
rect 321 402 324 405 
rect 321 405 324 408 
rect 321 408 324 411 
rect 321 411 324 414 
rect 321 414 324 417 
rect 321 417 324 420 
rect 321 420 324 423 
rect 321 423 324 426 
rect 321 426 324 429 
rect 321 429 324 432 
rect 321 432 324 435 
rect 321 435 324 438 
rect 321 438 324 441 
rect 321 441 324 444 
rect 321 444 324 447 
rect 321 447 324 450 
rect 321 450 324 453 
rect 321 453 324 456 
rect 321 456 324 459 
rect 321 459 324 462 
rect 321 462 324 465 
rect 321 465 324 468 
rect 321 468 324 471 
rect 321 471 324 474 
rect 321 474 324 477 
rect 321 477 324 480 
rect 321 480 324 483 
rect 321 483 324 486 
rect 321 486 324 489 
rect 321 489 324 492 
rect 321 492 324 495 
rect 321 495 324 498 
rect 321 498 324 501 
rect 321 501 324 504 
rect 321 504 324 507 
rect 321 507 324 510 
rect 324 0 327 3 
rect 324 3 327 6 
rect 324 6 327 9 
rect 324 9 327 12 
rect 324 12 327 15 
rect 324 15 327 18 
rect 324 18 327 21 
rect 324 21 327 24 
rect 324 24 327 27 
rect 324 27 327 30 
rect 324 30 327 33 
rect 324 33 327 36 
rect 324 36 327 39 
rect 324 39 327 42 
rect 324 42 327 45 
rect 324 45 327 48 
rect 324 48 327 51 
rect 324 51 327 54 
rect 324 54 327 57 
rect 324 57 327 60 
rect 324 60 327 63 
rect 324 63 327 66 
rect 324 66 327 69 
rect 324 69 327 72 
rect 324 72 327 75 
rect 324 75 327 78 
rect 324 78 327 81 
rect 324 81 327 84 
rect 324 84 327 87 
rect 324 87 327 90 
rect 324 90 327 93 
rect 324 93 327 96 
rect 324 96 327 99 
rect 324 99 327 102 
rect 324 102 327 105 
rect 324 105 327 108 
rect 324 108 327 111 
rect 324 111 327 114 
rect 324 114 327 117 
rect 324 117 327 120 
rect 324 120 327 123 
rect 324 123 327 126 
rect 324 126 327 129 
rect 324 129 327 132 
rect 324 132 327 135 
rect 324 135 327 138 
rect 324 138 327 141 
rect 324 141 327 144 
rect 324 144 327 147 
rect 324 147 327 150 
rect 324 150 327 153 
rect 324 153 327 156 
rect 324 156 327 159 
rect 324 159 327 162 
rect 324 162 327 165 
rect 324 165 327 168 
rect 324 168 327 171 
rect 324 171 327 174 
rect 324 174 327 177 
rect 324 177 327 180 
rect 324 180 327 183 
rect 324 183 327 186 
rect 324 186 327 189 
rect 324 189 327 192 
rect 324 192 327 195 
rect 324 195 327 198 
rect 324 198 327 201 
rect 324 201 327 204 
rect 324 204 327 207 
rect 324 207 327 210 
rect 324 210 327 213 
rect 324 213 327 216 
rect 324 216 327 219 
rect 324 219 327 222 
rect 324 222 327 225 
rect 324 225 327 228 
rect 324 228 327 231 
rect 324 231 327 234 
rect 324 234 327 237 
rect 324 237 327 240 
rect 324 240 327 243 
rect 324 243 327 246 
rect 324 246 327 249 
rect 324 249 327 252 
rect 324 252 327 255 
rect 324 255 327 258 
rect 324 258 327 261 
rect 324 261 327 264 
rect 324 264 327 267 
rect 324 267 327 270 
rect 324 270 327 273 
rect 324 273 327 276 
rect 324 276 327 279 
rect 324 279 327 282 
rect 324 282 327 285 
rect 324 285 327 288 
rect 324 288 327 291 
rect 324 291 327 294 
rect 324 294 327 297 
rect 324 297 327 300 
rect 324 300 327 303 
rect 324 303 327 306 
rect 324 306 327 309 
rect 324 309 327 312 
rect 324 312 327 315 
rect 324 315 327 318 
rect 324 318 327 321 
rect 324 321 327 324 
rect 324 324 327 327 
rect 324 327 327 330 
rect 324 330 327 333 
rect 324 333 327 336 
rect 324 336 327 339 
rect 324 339 327 342 
rect 324 342 327 345 
rect 324 345 327 348 
rect 324 348 327 351 
rect 324 351 327 354 
rect 324 354 327 357 
rect 324 357 327 360 
rect 324 360 327 363 
rect 324 363 327 366 
rect 324 366 327 369 
rect 324 369 327 372 
rect 324 372 327 375 
rect 324 375 327 378 
rect 324 378 327 381 
rect 324 381 327 384 
rect 324 384 327 387 
rect 324 387 327 390 
rect 324 390 327 393 
rect 324 393 327 396 
rect 324 396 327 399 
rect 324 399 327 402 
rect 324 402 327 405 
rect 324 405 327 408 
rect 324 408 327 411 
rect 324 411 327 414 
rect 324 414 327 417 
rect 324 417 327 420 
rect 324 420 327 423 
rect 324 423 327 426 
rect 324 426 327 429 
rect 324 429 327 432 
rect 324 432 327 435 
rect 324 435 327 438 
rect 324 438 327 441 
rect 324 441 327 444 
rect 324 444 327 447 
rect 324 447 327 450 
rect 324 450 327 453 
rect 324 453 327 456 
rect 324 456 327 459 
rect 324 459 327 462 
rect 324 462 327 465 
rect 324 465 327 468 
rect 324 468 327 471 
rect 324 471 327 474 
rect 324 474 327 477 
rect 324 477 327 480 
rect 324 480 327 483 
rect 324 483 327 486 
rect 324 486 327 489 
rect 324 489 327 492 
rect 324 492 327 495 
rect 324 495 327 498 
rect 324 498 327 501 
rect 324 501 327 504 
rect 324 504 327 507 
rect 324 507 327 510 
rect 327 0 330 3 
rect 327 3 330 6 
rect 327 6 330 9 
rect 327 9 330 12 
rect 327 12 330 15 
rect 327 15 330 18 
rect 327 18 330 21 
rect 327 21 330 24 
rect 327 24 330 27 
rect 327 27 330 30 
rect 327 30 330 33 
rect 327 33 330 36 
rect 327 36 330 39 
rect 327 39 330 42 
rect 327 42 330 45 
rect 327 45 330 48 
rect 327 48 330 51 
rect 327 51 330 54 
rect 327 54 330 57 
rect 327 57 330 60 
rect 327 60 330 63 
rect 327 63 330 66 
rect 327 66 330 69 
rect 327 69 330 72 
rect 327 72 330 75 
rect 327 75 330 78 
rect 327 78 330 81 
rect 327 81 330 84 
rect 327 84 330 87 
rect 327 87 330 90 
rect 327 90 330 93 
rect 327 93 330 96 
rect 327 96 330 99 
rect 327 99 330 102 
rect 327 102 330 105 
rect 327 105 330 108 
rect 327 108 330 111 
rect 327 111 330 114 
rect 327 114 330 117 
rect 327 117 330 120 
rect 327 120 330 123 
rect 327 123 330 126 
rect 327 126 330 129 
rect 327 129 330 132 
rect 327 132 330 135 
rect 327 135 330 138 
rect 327 138 330 141 
rect 327 141 330 144 
rect 327 144 330 147 
rect 327 147 330 150 
rect 327 150 330 153 
rect 327 153 330 156 
rect 327 156 330 159 
rect 327 159 330 162 
rect 327 162 330 165 
rect 327 165 330 168 
rect 327 168 330 171 
rect 327 171 330 174 
rect 327 174 330 177 
rect 327 177 330 180 
rect 327 180 330 183 
rect 327 183 330 186 
rect 327 186 330 189 
rect 327 189 330 192 
rect 327 192 330 195 
rect 327 195 330 198 
rect 327 198 330 201 
rect 327 201 330 204 
rect 327 204 330 207 
rect 327 207 330 210 
rect 327 210 330 213 
rect 327 213 330 216 
rect 327 216 330 219 
rect 327 219 330 222 
rect 327 222 330 225 
rect 327 225 330 228 
rect 327 228 330 231 
rect 327 231 330 234 
rect 327 234 330 237 
rect 327 237 330 240 
rect 327 240 330 243 
rect 327 243 330 246 
rect 327 246 330 249 
rect 327 249 330 252 
rect 327 252 330 255 
rect 327 255 330 258 
rect 327 258 330 261 
rect 327 261 330 264 
rect 327 264 330 267 
rect 327 267 330 270 
rect 327 270 330 273 
rect 327 273 330 276 
rect 327 276 330 279 
rect 327 279 330 282 
rect 327 282 330 285 
rect 327 285 330 288 
rect 327 288 330 291 
rect 327 291 330 294 
rect 327 294 330 297 
rect 327 297 330 300 
rect 327 300 330 303 
rect 327 303 330 306 
rect 327 306 330 309 
rect 327 309 330 312 
rect 327 312 330 315 
rect 327 315 330 318 
rect 327 318 330 321 
rect 327 321 330 324 
rect 327 324 330 327 
rect 327 327 330 330 
rect 327 330 330 333 
rect 327 333 330 336 
rect 327 336 330 339 
rect 327 339 330 342 
rect 327 342 330 345 
rect 327 345 330 348 
rect 327 348 330 351 
rect 327 351 330 354 
rect 327 354 330 357 
rect 327 357 330 360 
rect 327 360 330 363 
rect 327 363 330 366 
rect 327 366 330 369 
rect 327 369 330 372 
rect 327 372 330 375 
rect 327 375 330 378 
rect 327 378 330 381 
rect 327 381 330 384 
rect 327 384 330 387 
rect 327 387 330 390 
rect 327 390 330 393 
rect 327 393 330 396 
rect 327 396 330 399 
rect 327 399 330 402 
rect 327 402 330 405 
rect 327 405 330 408 
rect 327 408 330 411 
rect 327 411 330 414 
rect 327 414 330 417 
rect 327 417 330 420 
rect 327 420 330 423 
rect 327 423 330 426 
rect 327 426 330 429 
rect 327 429 330 432 
rect 327 432 330 435 
rect 327 435 330 438 
rect 327 438 330 441 
rect 327 441 330 444 
rect 327 444 330 447 
rect 327 447 330 450 
rect 327 450 330 453 
rect 327 453 330 456 
rect 327 456 330 459 
rect 327 459 330 462 
rect 327 462 330 465 
rect 327 465 330 468 
rect 327 468 330 471 
rect 327 471 330 474 
rect 327 474 330 477 
rect 327 477 330 480 
rect 327 480 330 483 
rect 327 483 330 486 
rect 327 486 330 489 
rect 327 489 330 492 
rect 327 492 330 495 
rect 327 495 330 498 
rect 327 498 330 501 
rect 327 501 330 504 
rect 327 504 330 507 
rect 327 507 330 510 
rect 330 0 333 3 
rect 330 3 333 6 
rect 330 6 333 9 
rect 330 9 333 12 
rect 330 12 333 15 
rect 330 15 333 18 
rect 330 18 333 21 
rect 330 21 333 24 
rect 330 24 333 27 
rect 330 27 333 30 
rect 330 30 333 33 
rect 330 33 333 36 
rect 330 36 333 39 
rect 330 39 333 42 
rect 330 42 333 45 
rect 330 45 333 48 
rect 330 48 333 51 
rect 330 51 333 54 
rect 330 54 333 57 
rect 330 57 333 60 
rect 330 60 333 63 
rect 330 63 333 66 
rect 330 66 333 69 
rect 330 69 333 72 
rect 330 72 333 75 
rect 330 75 333 78 
rect 330 78 333 81 
rect 330 81 333 84 
rect 330 84 333 87 
rect 330 87 333 90 
rect 330 90 333 93 
rect 330 93 333 96 
rect 330 96 333 99 
rect 330 99 333 102 
rect 330 102 333 105 
rect 330 105 333 108 
rect 330 108 333 111 
rect 330 111 333 114 
rect 330 114 333 117 
rect 330 117 333 120 
rect 330 120 333 123 
rect 330 123 333 126 
rect 330 126 333 129 
rect 330 129 333 132 
rect 330 132 333 135 
rect 330 135 333 138 
rect 330 138 333 141 
rect 330 141 333 144 
rect 330 144 333 147 
rect 330 147 333 150 
rect 330 150 333 153 
rect 330 153 333 156 
rect 330 156 333 159 
rect 330 159 333 162 
rect 330 162 333 165 
rect 330 165 333 168 
rect 330 168 333 171 
rect 330 171 333 174 
rect 330 174 333 177 
rect 330 177 333 180 
rect 330 180 333 183 
rect 330 183 333 186 
rect 330 186 333 189 
rect 330 189 333 192 
rect 330 192 333 195 
rect 330 195 333 198 
rect 330 198 333 201 
rect 330 201 333 204 
rect 330 204 333 207 
rect 330 207 333 210 
rect 330 210 333 213 
rect 330 213 333 216 
rect 330 216 333 219 
rect 330 219 333 222 
rect 330 222 333 225 
rect 330 225 333 228 
rect 330 228 333 231 
rect 330 231 333 234 
rect 330 234 333 237 
rect 330 237 333 240 
rect 330 240 333 243 
rect 330 243 333 246 
rect 330 246 333 249 
rect 330 249 333 252 
rect 330 252 333 255 
rect 330 255 333 258 
rect 330 258 333 261 
rect 330 261 333 264 
rect 330 264 333 267 
rect 330 267 333 270 
rect 330 270 333 273 
rect 330 273 333 276 
rect 330 276 333 279 
rect 330 279 333 282 
rect 330 282 333 285 
rect 330 285 333 288 
rect 330 288 333 291 
rect 330 291 333 294 
rect 330 294 333 297 
rect 330 297 333 300 
rect 330 300 333 303 
rect 330 303 333 306 
rect 330 306 333 309 
rect 330 309 333 312 
rect 330 312 333 315 
rect 330 315 333 318 
rect 330 318 333 321 
rect 330 321 333 324 
rect 330 324 333 327 
rect 330 327 333 330 
rect 330 330 333 333 
rect 330 333 333 336 
rect 330 336 333 339 
rect 330 339 333 342 
rect 330 342 333 345 
rect 330 345 333 348 
rect 330 348 333 351 
rect 330 351 333 354 
rect 330 354 333 357 
rect 330 357 333 360 
rect 330 360 333 363 
rect 330 363 333 366 
rect 330 366 333 369 
rect 330 369 333 372 
rect 330 372 333 375 
rect 330 375 333 378 
rect 330 378 333 381 
rect 330 381 333 384 
rect 330 384 333 387 
rect 330 387 333 390 
rect 330 390 333 393 
rect 330 393 333 396 
rect 330 396 333 399 
rect 330 399 333 402 
rect 330 402 333 405 
rect 330 405 333 408 
rect 330 408 333 411 
rect 330 411 333 414 
rect 330 414 333 417 
rect 330 417 333 420 
rect 330 420 333 423 
rect 330 423 333 426 
rect 330 426 333 429 
rect 330 429 333 432 
rect 330 432 333 435 
rect 330 435 333 438 
rect 330 438 333 441 
rect 330 441 333 444 
rect 330 444 333 447 
rect 330 447 333 450 
rect 330 450 333 453 
rect 330 453 333 456 
rect 330 456 333 459 
rect 330 459 333 462 
rect 330 462 333 465 
rect 330 465 333 468 
rect 330 468 333 471 
rect 330 471 333 474 
rect 330 474 333 477 
rect 330 477 333 480 
rect 330 480 333 483 
rect 330 483 333 486 
rect 330 486 333 489 
rect 330 489 333 492 
rect 330 492 333 495 
rect 330 495 333 498 
rect 330 498 333 501 
rect 330 501 333 504 
rect 330 504 333 507 
rect 330 507 333 510 
rect 333 0 336 3 
rect 333 3 336 6 
rect 333 6 336 9 
rect 333 9 336 12 
rect 333 12 336 15 
rect 333 15 336 18 
rect 333 18 336 21 
rect 333 21 336 24 
rect 333 24 336 27 
rect 333 27 336 30 
rect 333 30 336 33 
rect 333 33 336 36 
rect 333 36 336 39 
rect 333 39 336 42 
rect 333 42 336 45 
rect 333 45 336 48 
rect 333 48 336 51 
rect 333 51 336 54 
rect 333 54 336 57 
rect 333 57 336 60 
rect 333 60 336 63 
rect 333 63 336 66 
rect 333 66 336 69 
rect 333 69 336 72 
rect 333 72 336 75 
rect 333 75 336 78 
rect 333 78 336 81 
rect 333 81 336 84 
rect 333 84 336 87 
rect 333 87 336 90 
rect 333 90 336 93 
rect 333 93 336 96 
rect 333 96 336 99 
rect 333 99 336 102 
rect 333 102 336 105 
rect 333 105 336 108 
rect 333 108 336 111 
rect 333 111 336 114 
rect 333 114 336 117 
rect 333 117 336 120 
rect 333 120 336 123 
rect 333 123 336 126 
rect 333 126 336 129 
rect 333 129 336 132 
rect 333 132 336 135 
rect 333 135 336 138 
rect 333 138 336 141 
rect 333 141 336 144 
rect 333 144 336 147 
rect 333 147 336 150 
rect 333 150 336 153 
rect 333 153 336 156 
rect 333 156 336 159 
rect 333 159 336 162 
rect 333 162 336 165 
rect 333 165 336 168 
rect 333 168 336 171 
rect 333 171 336 174 
rect 333 174 336 177 
rect 333 177 336 180 
rect 333 180 336 183 
rect 333 183 336 186 
rect 333 186 336 189 
rect 333 189 336 192 
rect 333 192 336 195 
rect 333 195 336 198 
rect 333 198 336 201 
rect 333 201 336 204 
rect 333 204 336 207 
rect 333 207 336 210 
rect 333 210 336 213 
rect 333 213 336 216 
rect 333 216 336 219 
rect 333 219 336 222 
rect 333 222 336 225 
rect 333 225 336 228 
rect 333 228 336 231 
rect 333 231 336 234 
rect 333 234 336 237 
rect 333 237 336 240 
rect 333 240 336 243 
rect 333 243 336 246 
rect 333 246 336 249 
rect 333 249 336 252 
rect 333 252 336 255 
rect 333 255 336 258 
rect 333 258 336 261 
rect 333 261 336 264 
rect 333 264 336 267 
rect 333 267 336 270 
rect 333 270 336 273 
rect 333 273 336 276 
rect 333 276 336 279 
rect 333 279 336 282 
rect 333 282 336 285 
rect 333 285 336 288 
rect 333 288 336 291 
rect 333 291 336 294 
rect 333 294 336 297 
rect 333 297 336 300 
rect 333 300 336 303 
rect 333 303 336 306 
rect 333 306 336 309 
rect 333 309 336 312 
rect 333 312 336 315 
rect 333 315 336 318 
rect 333 318 336 321 
rect 333 321 336 324 
rect 333 324 336 327 
rect 333 327 336 330 
rect 333 330 336 333 
rect 333 333 336 336 
rect 333 336 336 339 
rect 333 339 336 342 
rect 333 342 336 345 
rect 333 345 336 348 
rect 333 348 336 351 
rect 333 351 336 354 
rect 333 354 336 357 
rect 333 357 336 360 
rect 333 360 336 363 
rect 333 363 336 366 
rect 333 366 336 369 
rect 333 369 336 372 
rect 333 372 336 375 
rect 333 375 336 378 
rect 333 378 336 381 
rect 333 381 336 384 
rect 333 384 336 387 
rect 333 387 336 390 
rect 333 390 336 393 
rect 333 393 336 396 
rect 333 396 336 399 
rect 333 399 336 402 
rect 333 402 336 405 
rect 333 405 336 408 
rect 333 408 336 411 
rect 333 411 336 414 
rect 333 414 336 417 
rect 333 417 336 420 
rect 333 420 336 423 
rect 333 423 336 426 
rect 333 426 336 429 
rect 333 429 336 432 
rect 333 432 336 435 
rect 333 435 336 438 
rect 333 438 336 441 
rect 333 441 336 444 
rect 333 444 336 447 
rect 333 447 336 450 
rect 333 450 336 453 
rect 333 453 336 456 
rect 333 456 336 459 
rect 333 459 336 462 
rect 333 462 336 465 
rect 333 465 336 468 
rect 333 468 336 471 
rect 333 471 336 474 
rect 333 474 336 477 
rect 333 477 336 480 
rect 333 480 336 483 
rect 333 483 336 486 
rect 333 486 336 489 
rect 333 489 336 492 
rect 333 492 336 495 
rect 333 495 336 498 
rect 333 498 336 501 
rect 333 501 336 504 
rect 333 504 336 507 
rect 333 507 336 510 
rect 336 0 339 3 
rect 336 3 339 6 
rect 336 6 339 9 
rect 336 9 339 12 
rect 336 12 339 15 
rect 336 15 339 18 
rect 336 18 339 21 
rect 336 21 339 24 
rect 336 24 339 27 
rect 336 27 339 30 
rect 336 30 339 33 
rect 336 33 339 36 
rect 336 36 339 39 
rect 336 39 339 42 
rect 336 42 339 45 
rect 336 45 339 48 
rect 336 48 339 51 
rect 336 51 339 54 
rect 336 54 339 57 
rect 336 57 339 60 
rect 336 60 339 63 
rect 336 63 339 66 
rect 336 66 339 69 
rect 336 69 339 72 
rect 336 72 339 75 
rect 336 75 339 78 
rect 336 78 339 81 
rect 336 81 339 84 
rect 336 84 339 87 
rect 336 87 339 90 
rect 336 90 339 93 
rect 336 93 339 96 
rect 336 96 339 99 
rect 336 99 339 102 
rect 336 102 339 105 
rect 336 105 339 108 
rect 336 108 339 111 
rect 336 111 339 114 
rect 336 114 339 117 
rect 336 117 339 120 
rect 336 120 339 123 
rect 336 123 339 126 
rect 336 126 339 129 
rect 336 129 339 132 
rect 336 132 339 135 
rect 336 135 339 138 
rect 336 138 339 141 
rect 336 141 339 144 
rect 336 144 339 147 
rect 336 147 339 150 
rect 336 150 339 153 
rect 336 153 339 156 
rect 336 156 339 159 
rect 336 159 339 162 
rect 336 162 339 165 
rect 336 165 339 168 
rect 336 168 339 171 
rect 336 171 339 174 
rect 336 174 339 177 
rect 336 177 339 180 
rect 336 180 339 183 
rect 336 183 339 186 
rect 336 186 339 189 
rect 336 189 339 192 
rect 336 192 339 195 
rect 336 195 339 198 
rect 336 198 339 201 
rect 336 201 339 204 
rect 336 204 339 207 
rect 336 207 339 210 
rect 336 210 339 213 
rect 336 213 339 216 
rect 336 216 339 219 
rect 336 219 339 222 
rect 336 222 339 225 
rect 336 225 339 228 
rect 336 228 339 231 
rect 336 231 339 234 
rect 336 234 339 237 
rect 336 237 339 240 
rect 336 240 339 243 
rect 336 243 339 246 
rect 336 246 339 249 
rect 336 249 339 252 
rect 336 252 339 255 
rect 336 255 339 258 
rect 336 258 339 261 
rect 336 261 339 264 
rect 336 264 339 267 
rect 336 267 339 270 
rect 336 270 339 273 
rect 336 273 339 276 
rect 336 276 339 279 
rect 336 279 339 282 
rect 336 282 339 285 
rect 336 285 339 288 
rect 336 288 339 291 
rect 336 291 339 294 
rect 336 294 339 297 
rect 336 297 339 300 
rect 336 300 339 303 
rect 336 303 339 306 
rect 336 306 339 309 
rect 336 309 339 312 
rect 336 312 339 315 
rect 336 315 339 318 
rect 336 318 339 321 
rect 336 321 339 324 
rect 336 324 339 327 
rect 336 327 339 330 
rect 336 330 339 333 
rect 336 333 339 336 
rect 336 336 339 339 
rect 336 339 339 342 
rect 336 342 339 345 
rect 336 345 339 348 
rect 336 348 339 351 
rect 336 351 339 354 
rect 336 354 339 357 
rect 336 357 339 360 
rect 336 360 339 363 
rect 336 363 339 366 
rect 336 366 339 369 
rect 336 369 339 372 
rect 336 372 339 375 
rect 336 375 339 378 
rect 336 378 339 381 
rect 336 381 339 384 
rect 336 384 339 387 
rect 336 387 339 390 
rect 336 390 339 393 
rect 336 393 339 396 
rect 336 396 339 399 
rect 336 399 339 402 
rect 336 402 339 405 
rect 336 405 339 408 
rect 336 408 339 411 
rect 336 411 339 414 
rect 336 414 339 417 
rect 336 417 339 420 
rect 336 420 339 423 
rect 336 423 339 426 
rect 336 426 339 429 
rect 336 429 339 432 
rect 336 432 339 435 
rect 336 435 339 438 
rect 336 438 339 441 
rect 336 441 339 444 
rect 336 444 339 447 
rect 336 447 339 450 
rect 336 450 339 453 
rect 336 453 339 456 
rect 336 456 339 459 
rect 336 459 339 462 
rect 336 462 339 465 
rect 336 465 339 468 
rect 336 468 339 471 
rect 336 471 339 474 
rect 336 474 339 477 
rect 336 477 339 480 
rect 336 480 339 483 
rect 336 483 339 486 
rect 336 486 339 489 
rect 336 489 339 492 
rect 336 492 339 495 
rect 336 495 339 498 
rect 336 498 339 501 
rect 336 501 339 504 
rect 336 504 339 507 
rect 336 507 339 510 
rect 339 0 342 3 
rect 339 3 342 6 
rect 339 6 342 9 
rect 339 9 342 12 
rect 339 12 342 15 
rect 339 15 342 18 
rect 339 18 342 21 
rect 339 21 342 24 
rect 339 24 342 27 
rect 339 27 342 30 
rect 339 30 342 33 
rect 339 33 342 36 
rect 339 36 342 39 
rect 339 39 342 42 
rect 339 42 342 45 
rect 339 45 342 48 
rect 339 48 342 51 
rect 339 51 342 54 
rect 339 54 342 57 
rect 339 57 342 60 
rect 339 60 342 63 
rect 339 63 342 66 
rect 339 66 342 69 
rect 339 69 342 72 
rect 339 72 342 75 
rect 339 75 342 78 
rect 339 78 342 81 
rect 339 81 342 84 
rect 339 84 342 87 
rect 339 87 342 90 
rect 339 90 342 93 
rect 339 93 342 96 
rect 339 96 342 99 
rect 339 99 342 102 
rect 339 102 342 105 
rect 339 105 342 108 
rect 339 108 342 111 
rect 339 111 342 114 
rect 339 114 342 117 
rect 339 117 342 120 
rect 339 120 342 123 
rect 339 123 342 126 
rect 339 126 342 129 
rect 339 129 342 132 
rect 339 132 342 135 
rect 339 135 342 138 
rect 339 138 342 141 
rect 339 141 342 144 
rect 339 144 342 147 
rect 339 147 342 150 
rect 339 150 342 153 
rect 339 153 342 156 
rect 339 156 342 159 
rect 339 159 342 162 
rect 339 162 342 165 
rect 339 165 342 168 
rect 339 168 342 171 
rect 339 171 342 174 
rect 339 174 342 177 
rect 339 177 342 180 
rect 339 180 342 183 
rect 339 183 342 186 
rect 339 186 342 189 
rect 339 189 342 192 
rect 339 192 342 195 
rect 339 195 342 198 
rect 339 198 342 201 
rect 339 201 342 204 
rect 339 204 342 207 
rect 339 207 342 210 
rect 339 210 342 213 
rect 339 213 342 216 
rect 339 216 342 219 
rect 339 219 342 222 
rect 339 222 342 225 
rect 339 225 342 228 
rect 339 228 342 231 
rect 339 231 342 234 
rect 339 234 342 237 
rect 339 237 342 240 
rect 339 240 342 243 
rect 339 243 342 246 
rect 339 246 342 249 
rect 339 249 342 252 
rect 339 252 342 255 
rect 339 255 342 258 
rect 339 258 342 261 
rect 339 261 342 264 
rect 339 264 342 267 
rect 339 267 342 270 
rect 339 270 342 273 
rect 339 273 342 276 
rect 339 276 342 279 
rect 339 279 342 282 
rect 339 282 342 285 
rect 339 285 342 288 
rect 339 288 342 291 
rect 339 291 342 294 
rect 339 294 342 297 
rect 339 297 342 300 
rect 339 300 342 303 
rect 339 303 342 306 
rect 339 306 342 309 
rect 339 309 342 312 
rect 339 312 342 315 
rect 339 315 342 318 
rect 339 318 342 321 
rect 339 321 342 324 
rect 339 324 342 327 
rect 339 327 342 330 
rect 339 330 342 333 
rect 339 333 342 336 
rect 339 336 342 339 
rect 339 339 342 342 
rect 339 342 342 345 
rect 339 345 342 348 
rect 339 348 342 351 
rect 339 351 342 354 
rect 339 354 342 357 
rect 339 357 342 360 
rect 339 360 342 363 
rect 339 363 342 366 
rect 339 366 342 369 
rect 339 369 342 372 
rect 339 372 342 375 
rect 339 375 342 378 
rect 339 378 342 381 
rect 339 381 342 384 
rect 339 384 342 387 
rect 339 387 342 390 
rect 339 390 342 393 
rect 339 393 342 396 
rect 339 396 342 399 
rect 339 399 342 402 
rect 339 402 342 405 
rect 339 405 342 408 
rect 339 408 342 411 
rect 339 411 342 414 
rect 339 414 342 417 
rect 339 417 342 420 
rect 339 420 342 423 
rect 339 423 342 426 
rect 339 426 342 429 
rect 339 429 342 432 
rect 339 432 342 435 
rect 339 435 342 438 
rect 339 438 342 441 
rect 339 441 342 444 
rect 339 444 342 447 
rect 339 447 342 450 
rect 339 450 342 453 
rect 339 453 342 456 
rect 339 456 342 459 
rect 339 459 342 462 
rect 339 462 342 465 
rect 339 465 342 468 
rect 339 468 342 471 
rect 339 471 342 474 
rect 339 474 342 477 
rect 339 477 342 480 
rect 339 480 342 483 
rect 339 483 342 486 
rect 339 486 342 489 
rect 339 489 342 492 
rect 339 492 342 495 
rect 339 495 342 498 
rect 339 498 342 501 
rect 339 501 342 504 
rect 339 504 342 507 
rect 339 507 342 510 
rect 342 0 345 3 
rect 342 3 345 6 
rect 342 6 345 9 
rect 342 9 345 12 
rect 342 12 345 15 
rect 342 15 345 18 
rect 342 18 345 21 
rect 342 21 345 24 
rect 342 24 345 27 
rect 342 27 345 30 
rect 342 30 345 33 
rect 342 33 345 36 
rect 342 36 345 39 
rect 342 39 345 42 
rect 342 42 345 45 
rect 342 45 345 48 
rect 342 48 345 51 
rect 342 51 345 54 
rect 342 54 345 57 
rect 342 57 345 60 
rect 342 60 345 63 
rect 342 63 345 66 
rect 342 66 345 69 
rect 342 69 345 72 
rect 342 72 345 75 
rect 342 75 345 78 
rect 342 78 345 81 
rect 342 81 345 84 
rect 342 84 345 87 
rect 342 87 345 90 
rect 342 90 345 93 
rect 342 93 345 96 
rect 342 96 345 99 
rect 342 99 345 102 
rect 342 102 345 105 
rect 342 105 345 108 
rect 342 108 345 111 
rect 342 111 345 114 
rect 342 114 345 117 
rect 342 117 345 120 
rect 342 120 345 123 
rect 342 123 345 126 
rect 342 126 345 129 
rect 342 129 345 132 
rect 342 132 345 135 
rect 342 135 345 138 
rect 342 138 345 141 
rect 342 141 345 144 
rect 342 144 345 147 
rect 342 147 345 150 
rect 342 150 345 153 
rect 342 153 345 156 
rect 342 156 345 159 
rect 342 159 345 162 
rect 342 162 345 165 
rect 342 165 345 168 
rect 342 168 345 171 
rect 342 171 345 174 
rect 342 174 345 177 
rect 342 177 345 180 
rect 342 180 345 183 
rect 342 183 345 186 
rect 342 186 345 189 
rect 342 189 345 192 
rect 342 192 345 195 
rect 342 195 345 198 
rect 342 198 345 201 
rect 342 201 345 204 
rect 342 204 345 207 
rect 342 207 345 210 
rect 342 210 345 213 
rect 342 213 345 216 
rect 342 216 345 219 
rect 342 219 345 222 
rect 342 222 345 225 
rect 342 225 345 228 
rect 342 228 345 231 
rect 342 231 345 234 
rect 342 234 345 237 
rect 342 237 345 240 
rect 342 240 345 243 
rect 342 243 345 246 
rect 342 246 345 249 
rect 342 249 345 252 
rect 342 252 345 255 
rect 342 255 345 258 
rect 342 258 345 261 
rect 342 261 345 264 
rect 342 264 345 267 
rect 342 267 345 270 
rect 342 270 345 273 
rect 342 273 345 276 
rect 342 276 345 279 
rect 342 279 345 282 
rect 342 282 345 285 
rect 342 285 345 288 
rect 342 288 345 291 
rect 342 291 345 294 
rect 342 294 345 297 
rect 342 297 345 300 
rect 342 300 345 303 
rect 342 303 345 306 
rect 342 306 345 309 
rect 342 309 345 312 
rect 342 312 345 315 
rect 342 315 345 318 
rect 342 318 345 321 
rect 342 321 345 324 
rect 342 324 345 327 
rect 342 327 345 330 
rect 342 330 345 333 
rect 342 333 345 336 
rect 342 336 345 339 
rect 342 339 345 342 
rect 342 342 345 345 
rect 342 345 345 348 
rect 342 348 345 351 
rect 342 351 345 354 
rect 342 354 345 357 
rect 342 357 345 360 
rect 342 360 345 363 
rect 342 363 345 366 
rect 342 366 345 369 
rect 342 369 345 372 
rect 342 372 345 375 
rect 342 375 345 378 
rect 342 378 345 381 
rect 342 381 345 384 
rect 342 384 345 387 
rect 342 387 345 390 
rect 342 390 345 393 
rect 342 393 345 396 
rect 342 396 345 399 
rect 342 399 345 402 
rect 342 402 345 405 
rect 342 405 345 408 
rect 342 408 345 411 
rect 342 411 345 414 
rect 342 414 345 417 
rect 342 417 345 420 
rect 342 420 345 423 
rect 342 423 345 426 
rect 342 426 345 429 
rect 342 429 345 432 
rect 342 432 345 435 
rect 342 435 345 438 
rect 342 438 345 441 
rect 342 441 345 444 
rect 342 444 345 447 
rect 342 447 345 450 
rect 342 450 345 453 
rect 342 453 345 456 
rect 342 456 345 459 
rect 342 459 345 462 
rect 342 462 345 465 
rect 342 465 345 468 
rect 342 468 345 471 
rect 342 471 345 474 
rect 342 474 345 477 
rect 342 477 345 480 
rect 342 480 345 483 
rect 342 483 345 486 
rect 342 486 345 489 
rect 342 489 345 492 
rect 342 492 345 495 
rect 342 495 345 498 
rect 342 498 345 501 
rect 342 501 345 504 
rect 342 504 345 507 
rect 342 507 345 510 
rect 345 0 348 3 
rect 345 3 348 6 
rect 345 6 348 9 
rect 345 9 348 12 
rect 345 12 348 15 
rect 345 15 348 18 
rect 345 18 348 21 
rect 345 21 348 24 
rect 345 24 348 27 
rect 345 27 348 30 
rect 345 30 348 33 
rect 345 33 348 36 
rect 345 36 348 39 
rect 345 39 348 42 
rect 345 42 348 45 
rect 345 45 348 48 
rect 345 48 348 51 
rect 345 51 348 54 
rect 345 54 348 57 
rect 345 57 348 60 
rect 345 60 348 63 
rect 345 63 348 66 
rect 345 66 348 69 
rect 345 69 348 72 
rect 345 72 348 75 
rect 345 75 348 78 
rect 345 78 348 81 
rect 345 81 348 84 
rect 345 84 348 87 
rect 345 87 348 90 
rect 345 90 348 93 
rect 345 93 348 96 
rect 345 96 348 99 
rect 345 99 348 102 
rect 345 102 348 105 
rect 345 105 348 108 
rect 345 108 348 111 
rect 345 111 348 114 
rect 345 114 348 117 
rect 345 117 348 120 
rect 345 120 348 123 
rect 345 123 348 126 
rect 345 126 348 129 
rect 345 129 348 132 
rect 345 132 348 135 
rect 345 135 348 138 
rect 345 138 348 141 
rect 345 141 348 144 
rect 345 144 348 147 
rect 345 147 348 150 
rect 345 150 348 153 
rect 345 153 348 156 
rect 345 156 348 159 
rect 345 159 348 162 
rect 345 162 348 165 
rect 345 165 348 168 
rect 345 168 348 171 
rect 345 171 348 174 
rect 345 174 348 177 
rect 345 177 348 180 
rect 345 180 348 183 
rect 345 183 348 186 
rect 345 186 348 189 
rect 345 189 348 192 
rect 345 192 348 195 
rect 345 195 348 198 
rect 345 198 348 201 
rect 345 201 348 204 
rect 345 204 348 207 
rect 345 207 348 210 
rect 345 210 348 213 
rect 345 213 348 216 
rect 345 216 348 219 
rect 345 219 348 222 
rect 345 222 348 225 
rect 345 225 348 228 
rect 345 228 348 231 
rect 345 231 348 234 
rect 345 234 348 237 
rect 345 237 348 240 
rect 345 240 348 243 
rect 345 243 348 246 
rect 345 246 348 249 
rect 345 249 348 252 
rect 345 252 348 255 
rect 345 255 348 258 
rect 345 258 348 261 
rect 345 261 348 264 
rect 345 264 348 267 
rect 345 267 348 270 
rect 345 270 348 273 
rect 345 273 348 276 
rect 345 276 348 279 
rect 345 279 348 282 
rect 345 282 348 285 
rect 345 285 348 288 
rect 345 288 348 291 
rect 345 291 348 294 
rect 345 294 348 297 
rect 345 297 348 300 
rect 345 300 348 303 
rect 345 303 348 306 
rect 345 306 348 309 
rect 345 309 348 312 
rect 345 312 348 315 
rect 345 315 348 318 
rect 345 318 348 321 
rect 345 321 348 324 
rect 345 324 348 327 
rect 345 327 348 330 
rect 345 330 348 333 
rect 345 333 348 336 
rect 345 336 348 339 
rect 345 339 348 342 
rect 345 342 348 345 
rect 345 345 348 348 
rect 345 348 348 351 
rect 345 351 348 354 
rect 345 354 348 357 
rect 345 357 348 360 
rect 345 360 348 363 
rect 345 363 348 366 
rect 345 366 348 369 
rect 345 369 348 372 
rect 345 372 348 375 
rect 345 375 348 378 
rect 345 378 348 381 
rect 345 381 348 384 
rect 345 384 348 387 
rect 345 387 348 390 
rect 345 390 348 393 
rect 345 393 348 396 
rect 345 396 348 399 
rect 345 399 348 402 
rect 345 402 348 405 
rect 345 405 348 408 
rect 345 408 348 411 
rect 345 411 348 414 
rect 345 414 348 417 
rect 345 417 348 420 
rect 345 420 348 423 
rect 345 423 348 426 
rect 345 426 348 429 
rect 345 429 348 432 
rect 345 432 348 435 
rect 345 435 348 438 
rect 345 438 348 441 
rect 345 441 348 444 
rect 345 444 348 447 
rect 345 447 348 450 
rect 345 450 348 453 
rect 345 453 348 456 
rect 345 456 348 459 
rect 345 459 348 462 
rect 345 462 348 465 
rect 345 465 348 468 
rect 345 468 348 471 
rect 345 471 348 474 
rect 345 474 348 477 
rect 345 477 348 480 
rect 345 480 348 483 
rect 345 483 348 486 
rect 345 486 348 489 
rect 345 489 348 492 
rect 345 492 348 495 
rect 345 495 348 498 
rect 345 498 348 501 
rect 345 501 348 504 
rect 345 504 348 507 
rect 345 507 348 510 
rect 348 0 351 3 
rect 348 3 351 6 
rect 348 6 351 9 
rect 348 9 351 12 
rect 348 12 351 15 
rect 348 15 351 18 
rect 348 18 351 21 
rect 348 21 351 24 
rect 348 24 351 27 
rect 348 27 351 30 
rect 348 30 351 33 
rect 348 33 351 36 
rect 348 36 351 39 
rect 348 39 351 42 
rect 348 42 351 45 
rect 348 45 351 48 
rect 348 48 351 51 
rect 348 51 351 54 
rect 348 54 351 57 
rect 348 57 351 60 
rect 348 60 351 63 
rect 348 63 351 66 
rect 348 66 351 69 
rect 348 69 351 72 
rect 348 72 351 75 
rect 348 75 351 78 
rect 348 78 351 81 
rect 348 81 351 84 
rect 348 84 351 87 
rect 348 87 351 90 
rect 348 90 351 93 
rect 348 93 351 96 
rect 348 96 351 99 
rect 348 99 351 102 
rect 348 102 351 105 
rect 348 105 351 108 
rect 348 108 351 111 
rect 348 111 351 114 
rect 348 114 351 117 
rect 348 117 351 120 
rect 348 120 351 123 
rect 348 123 351 126 
rect 348 126 351 129 
rect 348 129 351 132 
rect 348 132 351 135 
rect 348 135 351 138 
rect 348 138 351 141 
rect 348 141 351 144 
rect 348 144 351 147 
rect 348 147 351 150 
rect 348 150 351 153 
rect 348 153 351 156 
rect 348 156 351 159 
rect 348 159 351 162 
rect 348 162 351 165 
rect 348 165 351 168 
rect 348 168 351 171 
rect 348 171 351 174 
rect 348 174 351 177 
rect 348 177 351 180 
rect 348 180 351 183 
rect 348 183 351 186 
rect 348 186 351 189 
rect 348 189 351 192 
rect 348 192 351 195 
rect 348 195 351 198 
rect 348 198 351 201 
rect 348 201 351 204 
rect 348 204 351 207 
rect 348 207 351 210 
rect 348 210 351 213 
rect 348 213 351 216 
rect 348 216 351 219 
rect 348 219 351 222 
rect 348 222 351 225 
rect 348 225 351 228 
rect 348 228 351 231 
rect 348 231 351 234 
rect 348 234 351 237 
rect 348 237 351 240 
rect 348 240 351 243 
rect 348 243 351 246 
rect 348 246 351 249 
rect 348 249 351 252 
rect 348 252 351 255 
rect 348 255 351 258 
rect 348 258 351 261 
rect 348 261 351 264 
rect 348 264 351 267 
rect 348 267 351 270 
rect 348 270 351 273 
rect 348 273 351 276 
rect 348 276 351 279 
rect 348 279 351 282 
rect 348 282 351 285 
rect 348 285 351 288 
rect 348 288 351 291 
rect 348 291 351 294 
rect 348 294 351 297 
rect 348 297 351 300 
rect 348 300 351 303 
rect 348 303 351 306 
rect 348 306 351 309 
rect 348 309 351 312 
rect 348 312 351 315 
rect 348 315 351 318 
rect 348 318 351 321 
rect 348 321 351 324 
rect 348 324 351 327 
rect 348 327 351 330 
rect 348 330 351 333 
rect 348 333 351 336 
rect 348 336 351 339 
rect 348 339 351 342 
rect 348 342 351 345 
rect 348 345 351 348 
rect 348 348 351 351 
rect 348 351 351 354 
rect 348 354 351 357 
rect 348 357 351 360 
rect 348 360 351 363 
rect 348 363 351 366 
rect 348 366 351 369 
rect 348 369 351 372 
rect 348 372 351 375 
rect 348 375 351 378 
rect 348 378 351 381 
rect 348 381 351 384 
rect 348 384 351 387 
rect 348 387 351 390 
rect 348 390 351 393 
rect 348 393 351 396 
rect 348 396 351 399 
rect 348 399 351 402 
rect 348 402 351 405 
rect 348 405 351 408 
rect 348 408 351 411 
rect 348 411 351 414 
rect 348 414 351 417 
rect 348 417 351 420 
rect 348 420 351 423 
rect 348 423 351 426 
rect 348 426 351 429 
rect 348 429 351 432 
rect 348 432 351 435 
rect 348 435 351 438 
rect 348 438 351 441 
rect 348 441 351 444 
rect 348 444 351 447 
rect 348 447 351 450 
rect 348 450 351 453 
rect 348 453 351 456 
rect 348 456 351 459 
rect 348 459 351 462 
rect 348 462 351 465 
rect 348 465 351 468 
rect 348 468 351 471 
rect 348 471 351 474 
rect 348 474 351 477 
rect 348 477 351 480 
rect 348 480 351 483 
rect 348 483 351 486 
rect 348 486 351 489 
rect 348 489 351 492 
rect 348 492 351 495 
rect 348 495 351 498 
rect 348 498 351 501 
rect 348 501 351 504 
rect 348 504 351 507 
rect 348 507 351 510 
rect 351 0 354 3 
rect 351 3 354 6 
rect 351 6 354 9 
rect 351 9 354 12 
rect 351 12 354 15 
rect 351 15 354 18 
rect 351 18 354 21 
rect 351 21 354 24 
rect 351 24 354 27 
rect 351 27 354 30 
rect 351 30 354 33 
rect 351 33 354 36 
rect 351 36 354 39 
rect 351 39 354 42 
rect 351 42 354 45 
rect 351 45 354 48 
rect 351 48 354 51 
rect 351 51 354 54 
rect 351 54 354 57 
rect 351 57 354 60 
rect 351 60 354 63 
rect 351 63 354 66 
rect 351 66 354 69 
rect 351 69 354 72 
rect 351 72 354 75 
rect 351 75 354 78 
rect 351 78 354 81 
rect 351 81 354 84 
rect 351 84 354 87 
rect 351 87 354 90 
rect 351 90 354 93 
rect 351 93 354 96 
rect 351 96 354 99 
rect 351 99 354 102 
rect 351 102 354 105 
rect 351 105 354 108 
rect 351 108 354 111 
rect 351 111 354 114 
rect 351 114 354 117 
rect 351 117 354 120 
rect 351 120 354 123 
rect 351 123 354 126 
rect 351 126 354 129 
rect 351 129 354 132 
rect 351 132 354 135 
rect 351 135 354 138 
rect 351 138 354 141 
rect 351 141 354 144 
rect 351 144 354 147 
rect 351 147 354 150 
rect 351 150 354 153 
rect 351 153 354 156 
rect 351 156 354 159 
rect 351 159 354 162 
rect 351 162 354 165 
rect 351 165 354 168 
rect 351 168 354 171 
rect 351 171 354 174 
rect 351 174 354 177 
rect 351 177 354 180 
rect 351 180 354 183 
rect 351 183 354 186 
rect 351 186 354 189 
rect 351 189 354 192 
rect 351 192 354 195 
rect 351 195 354 198 
rect 351 198 354 201 
rect 351 201 354 204 
rect 351 204 354 207 
rect 351 207 354 210 
rect 351 210 354 213 
rect 351 213 354 216 
rect 351 216 354 219 
rect 351 219 354 222 
rect 351 222 354 225 
rect 351 225 354 228 
rect 351 228 354 231 
rect 351 231 354 234 
rect 351 234 354 237 
rect 351 237 354 240 
rect 351 240 354 243 
rect 351 243 354 246 
rect 351 246 354 249 
rect 351 249 354 252 
rect 351 252 354 255 
rect 351 255 354 258 
rect 351 258 354 261 
rect 351 261 354 264 
rect 351 264 354 267 
rect 351 267 354 270 
rect 351 270 354 273 
rect 351 273 354 276 
rect 351 276 354 279 
rect 351 279 354 282 
rect 351 282 354 285 
rect 351 285 354 288 
rect 351 288 354 291 
rect 351 291 354 294 
rect 351 294 354 297 
rect 351 297 354 300 
rect 351 300 354 303 
rect 351 303 354 306 
rect 351 306 354 309 
rect 351 309 354 312 
rect 351 312 354 315 
rect 351 315 354 318 
rect 351 318 354 321 
rect 351 321 354 324 
rect 351 324 354 327 
rect 351 327 354 330 
rect 351 330 354 333 
rect 351 333 354 336 
rect 351 336 354 339 
rect 351 339 354 342 
rect 351 342 354 345 
rect 351 345 354 348 
rect 351 348 354 351 
rect 351 351 354 354 
rect 351 354 354 357 
rect 351 357 354 360 
rect 351 360 354 363 
rect 351 363 354 366 
rect 351 366 354 369 
rect 351 369 354 372 
rect 351 372 354 375 
rect 351 375 354 378 
rect 351 378 354 381 
rect 351 381 354 384 
rect 351 384 354 387 
rect 351 387 354 390 
rect 351 390 354 393 
rect 351 393 354 396 
rect 351 396 354 399 
rect 351 399 354 402 
rect 351 402 354 405 
rect 351 405 354 408 
rect 351 408 354 411 
rect 351 411 354 414 
rect 351 414 354 417 
rect 351 417 354 420 
rect 351 420 354 423 
rect 351 423 354 426 
rect 351 426 354 429 
rect 351 429 354 432 
rect 351 432 354 435 
rect 351 435 354 438 
rect 351 438 354 441 
rect 351 441 354 444 
rect 351 444 354 447 
rect 351 447 354 450 
rect 351 450 354 453 
rect 351 453 354 456 
rect 351 456 354 459 
rect 351 459 354 462 
rect 351 462 354 465 
rect 351 465 354 468 
rect 351 468 354 471 
rect 351 471 354 474 
rect 351 474 354 477 
rect 351 477 354 480 
rect 351 480 354 483 
rect 351 483 354 486 
rect 351 486 354 489 
rect 351 489 354 492 
rect 351 492 354 495 
rect 351 495 354 498 
rect 351 498 354 501 
rect 351 501 354 504 
rect 351 504 354 507 
rect 351 507 354 510 
rect 354 0 357 3 
rect 354 3 357 6 
rect 354 6 357 9 
rect 354 9 357 12 
rect 354 12 357 15 
rect 354 15 357 18 
rect 354 18 357 21 
rect 354 21 357 24 
rect 354 24 357 27 
rect 354 27 357 30 
rect 354 30 357 33 
rect 354 33 357 36 
rect 354 36 357 39 
rect 354 39 357 42 
rect 354 42 357 45 
rect 354 45 357 48 
rect 354 48 357 51 
rect 354 51 357 54 
rect 354 54 357 57 
rect 354 57 357 60 
rect 354 60 357 63 
rect 354 63 357 66 
rect 354 66 357 69 
rect 354 69 357 72 
rect 354 72 357 75 
rect 354 75 357 78 
rect 354 78 357 81 
rect 354 81 357 84 
rect 354 84 357 87 
rect 354 87 357 90 
rect 354 90 357 93 
rect 354 93 357 96 
rect 354 96 357 99 
rect 354 99 357 102 
rect 354 102 357 105 
rect 354 105 357 108 
rect 354 108 357 111 
rect 354 111 357 114 
rect 354 114 357 117 
rect 354 117 357 120 
rect 354 120 357 123 
rect 354 123 357 126 
rect 354 126 357 129 
rect 354 129 357 132 
rect 354 132 357 135 
rect 354 135 357 138 
rect 354 138 357 141 
rect 354 141 357 144 
rect 354 144 357 147 
rect 354 147 357 150 
rect 354 150 357 153 
rect 354 153 357 156 
rect 354 156 357 159 
rect 354 159 357 162 
rect 354 162 357 165 
rect 354 165 357 168 
rect 354 168 357 171 
rect 354 171 357 174 
rect 354 174 357 177 
rect 354 177 357 180 
rect 354 180 357 183 
rect 354 183 357 186 
rect 354 186 357 189 
rect 354 189 357 192 
rect 354 192 357 195 
rect 354 195 357 198 
rect 354 198 357 201 
rect 354 201 357 204 
rect 354 204 357 207 
rect 354 207 357 210 
rect 354 210 357 213 
rect 354 213 357 216 
rect 354 216 357 219 
rect 354 219 357 222 
rect 354 222 357 225 
rect 354 225 357 228 
rect 354 228 357 231 
rect 354 231 357 234 
rect 354 234 357 237 
rect 354 237 357 240 
rect 354 240 357 243 
rect 354 243 357 246 
rect 354 246 357 249 
rect 354 249 357 252 
rect 354 252 357 255 
rect 354 255 357 258 
rect 354 258 357 261 
rect 354 261 357 264 
rect 354 264 357 267 
rect 354 267 357 270 
rect 354 270 357 273 
rect 354 273 357 276 
rect 354 276 357 279 
rect 354 279 357 282 
rect 354 282 357 285 
rect 354 285 357 288 
rect 354 288 357 291 
rect 354 291 357 294 
rect 354 294 357 297 
rect 354 297 357 300 
rect 354 300 357 303 
rect 354 303 357 306 
rect 354 306 357 309 
rect 354 309 357 312 
rect 354 312 357 315 
rect 354 315 357 318 
rect 354 318 357 321 
rect 354 321 357 324 
rect 354 324 357 327 
rect 354 327 357 330 
rect 354 330 357 333 
rect 354 333 357 336 
rect 354 336 357 339 
rect 354 339 357 342 
rect 354 342 357 345 
rect 354 345 357 348 
rect 354 348 357 351 
rect 354 351 357 354 
rect 354 354 357 357 
rect 354 357 357 360 
rect 354 360 357 363 
rect 354 363 357 366 
rect 354 366 357 369 
rect 354 369 357 372 
rect 354 372 357 375 
rect 354 375 357 378 
rect 354 378 357 381 
rect 354 381 357 384 
rect 354 384 357 387 
rect 354 387 357 390 
rect 354 390 357 393 
rect 354 393 357 396 
rect 354 396 357 399 
rect 354 399 357 402 
rect 354 402 357 405 
rect 354 405 357 408 
rect 354 408 357 411 
rect 354 411 357 414 
rect 354 414 357 417 
rect 354 417 357 420 
rect 354 420 357 423 
rect 354 423 357 426 
rect 354 426 357 429 
rect 354 429 357 432 
rect 354 432 357 435 
rect 354 435 357 438 
rect 354 438 357 441 
rect 354 441 357 444 
rect 354 444 357 447 
rect 354 447 357 450 
rect 354 450 357 453 
rect 354 453 357 456 
rect 354 456 357 459 
rect 354 459 357 462 
rect 354 462 357 465 
rect 354 465 357 468 
rect 354 468 357 471 
rect 354 471 357 474 
rect 354 474 357 477 
rect 354 477 357 480 
rect 354 480 357 483 
rect 354 483 357 486 
rect 354 486 357 489 
rect 354 489 357 492 
rect 354 492 357 495 
rect 354 495 357 498 
rect 354 498 357 501 
rect 354 501 357 504 
rect 354 504 357 507 
rect 354 507 357 510 
rect 357 0 360 3 
rect 357 3 360 6 
rect 357 6 360 9 
rect 357 9 360 12 
rect 357 12 360 15 
rect 357 15 360 18 
rect 357 18 360 21 
rect 357 21 360 24 
rect 357 24 360 27 
rect 357 27 360 30 
rect 357 30 360 33 
rect 357 33 360 36 
rect 357 36 360 39 
rect 357 39 360 42 
rect 357 42 360 45 
rect 357 45 360 48 
rect 357 48 360 51 
rect 357 51 360 54 
rect 357 54 360 57 
rect 357 57 360 60 
rect 357 60 360 63 
rect 357 63 360 66 
rect 357 66 360 69 
rect 357 69 360 72 
rect 357 72 360 75 
rect 357 75 360 78 
rect 357 78 360 81 
rect 357 81 360 84 
rect 357 84 360 87 
rect 357 87 360 90 
rect 357 90 360 93 
rect 357 93 360 96 
rect 357 96 360 99 
rect 357 99 360 102 
rect 357 102 360 105 
rect 357 105 360 108 
rect 357 108 360 111 
rect 357 111 360 114 
rect 357 114 360 117 
rect 357 117 360 120 
rect 357 120 360 123 
rect 357 123 360 126 
rect 357 126 360 129 
rect 357 129 360 132 
rect 357 132 360 135 
rect 357 135 360 138 
rect 357 138 360 141 
rect 357 141 360 144 
rect 357 144 360 147 
rect 357 147 360 150 
rect 357 150 360 153 
rect 357 153 360 156 
rect 357 156 360 159 
rect 357 159 360 162 
rect 357 162 360 165 
rect 357 165 360 168 
rect 357 168 360 171 
rect 357 171 360 174 
rect 357 174 360 177 
rect 357 177 360 180 
rect 357 180 360 183 
rect 357 183 360 186 
rect 357 186 360 189 
rect 357 189 360 192 
rect 357 192 360 195 
rect 357 195 360 198 
rect 357 198 360 201 
rect 357 201 360 204 
rect 357 204 360 207 
rect 357 207 360 210 
rect 357 210 360 213 
rect 357 213 360 216 
rect 357 216 360 219 
rect 357 219 360 222 
rect 357 222 360 225 
rect 357 225 360 228 
rect 357 228 360 231 
rect 357 231 360 234 
rect 357 234 360 237 
rect 357 237 360 240 
rect 357 240 360 243 
rect 357 243 360 246 
rect 357 246 360 249 
rect 357 249 360 252 
rect 357 252 360 255 
rect 357 255 360 258 
rect 357 258 360 261 
rect 357 261 360 264 
rect 357 264 360 267 
rect 357 267 360 270 
rect 357 270 360 273 
rect 357 273 360 276 
rect 357 276 360 279 
rect 357 279 360 282 
rect 357 282 360 285 
rect 357 285 360 288 
rect 357 288 360 291 
rect 357 291 360 294 
rect 357 294 360 297 
rect 357 297 360 300 
rect 357 300 360 303 
rect 357 303 360 306 
rect 357 306 360 309 
rect 357 309 360 312 
rect 357 312 360 315 
rect 357 315 360 318 
rect 357 318 360 321 
rect 357 321 360 324 
rect 357 324 360 327 
rect 357 327 360 330 
rect 357 330 360 333 
rect 357 333 360 336 
rect 357 336 360 339 
rect 357 339 360 342 
rect 357 342 360 345 
rect 357 345 360 348 
rect 357 348 360 351 
rect 357 351 360 354 
rect 357 354 360 357 
rect 357 357 360 360 
rect 357 360 360 363 
rect 357 363 360 366 
rect 357 366 360 369 
rect 357 369 360 372 
rect 357 372 360 375 
rect 357 375 360 378 
rect 357 378 360 381 
rect 357 381 360 384 
rect 357 384 360 387 
rect 357 387 360 390 
rect 357 390 360 393 
rect 357 393 360 396 
rect 357 396 360 399 
rect 357 399 360 402 
rect 357 402 360 405 
rect 357 405 360 408 
rect 357 408 360 411 
rect 357 411 360 414 
rect 357 414 360 417 
rect 357 417 360 420 
rect 357 420 360 423 
rect 357 423 360 426 
rect 357 426 360 429 
rect 357 429 360 432 
rect 357 432 360 435 
rect 357 435 360 438 
rect 357 438 360 441 
rect 357 441 360 444 
rect 357 444 360 447 
rect 357 447 360 450 
rect 357 450 360 453 
rect 357 453 360 456 
rect 357 456 360 459 
rect 357 459 360 462 
rect 357 462 360 465 
rect 357 465 360 468 
rect 357 468 360 471 
rect 357 471 360 474 
rect 357 474 360 477 
rect 357 477 360 480 
rect 357 480 360 483 
rect 357 483 360 486 
rect 357 486 360 489 
rect 357 489 360 492 
rect 357 492 360 495 
rect 357 495 360 498 
rect 357 498 360 501 
rect 357 501 360 504 
rect 357 504 360 507 
rect 357 507 360 510 
rect 360 0 363 3 
rect 360 3 363 6 
rect 360 6 363 9 
rect 360 9 363 12 
rect 360 12 363 15 
rect 360 15 363 18 
rect 360 18 363 21 
rect 360 21 363 24 
rect 360 24 363 27 
rect 360 27 363 30 
rect 360 30 363 33 
rect 360 33 363 36 
rect 360 36 363 39 
rect 360 39 363 42 
rect 360 42 363 45 
rect 360 45 363 48 
rect 360 48 363 51 
rect 360 51 363 54 
rect 360 54 363 57 
rect 360 57 363 60 
rect 360 60 363 63 
rect 360 63 363 66 
rect 360 66 363 69 
rect 360 69 363 72 
rect 360 72 363 75 
rect 360 75 363 78 
rect 360 78 363 81 
rect 360 81 363 84 
rect 360 84 363 87 
rect 360 87 363 90 
rect 360 90 363 93 
rect 360 93 363 96 
rect 360 96 363 99 
rect 360 99 363 102 
rect 360 102 363 105 
rect 360 105 363 108 
rect 360 108 363 111 
rect 360 111 363 114 
rect 360 114 363 117 
rect 360 117 363 120 
rect 360 120 363 123 
rect 360 123 363 126 
rect 360 126 363 129 
rect 360 129 363 132 
rect 360 132 363 135 
rect 360 135 363 138 
rect 360 138 363 141 
rect 360 141 363 144 
rect 360 144 363 147 
rect 360 147 363 150 
rect 360 150 363 153 
rect 360 153 363 156 
rect 360 156 363 159 
rect 360 159 363 162 
rect 360 162 363 165 
rect 360 165 363 168 
rect 360 168 363 171 
rect 360 171 363 174 
rect 360 174 363 177 
rect 360 177 363 180 
rect 360 180 363 183 
rect 360 183 363 186 
rect 360 186 363 189 
rect 360 189 363 192 
rect 360 192 363 195 
rect 360 195 363 198 
rect 360 198 363 201 
rect 360 201 363 204 
rect 360 204 363 207 
rect 360 207 363 210 
rect 360 210 363 213 
rect 360 213 363 216 
rect 360 216 363 219 
rect 360 219 363 222 
rect 360 222 363 225 
rect 360 225 363 228 
rect 360 228 363 231 
rect 360 231 363 234 
rect 360 234 363 237 
rect 360 237 363 240 
rect 360 240 363 243 
rect 360 243 363 246 
rect 360 246 363 249 
rect 360 249 363 252 
rect 360 252 363 255 
rect 360 255 363 258 
rect 360 258 363 261 
rect 360 261 363 264 
rect 360 264 363 267 
rect 360 267 363 270 
rect 360 270 363 273 
rect 360 273 363 276 
rect 360 276 363 279 
rect 360 279 363 282 
rect 360 282 363 285 
rect 360 285 363 288 
rect 360 288 363 291 
rect 360 291 363 294 
rect 360 294 363 297 
rect 360 297 363 300 
rect 360 300 363 303 
rect 360 303 363 306 
rect 360 306 363 309 
rect 360 309 363 312 
rect 360 312 363 315 
rect 360 315 363 318 
rect 360 318 363 321 
rect 360 321 363 324 
rect 360 324 363 327 
rect 360 327 363 330 
rect 360 330 363 333 
rect 360 333 363 336 
rect 360 336 363 339 
rect 360 339 363 342 
rect 360 342 363 345 
rect 360 345 363 348 
rect 360 348 363 351 
rect 360 351 363 354 
rect 360 354 363 357 
rect 360 357 363 360 
rect 360 360 363 363 
rect 360 363 363 366 
rect 360 366 363 369 
rect 360 369 363 372 
rect 360 372 363 375 
rect 360 375 363 378 
rect 360 378 363 381 
rect 360 381 363 384 
rect 360 384 363 387 
rect 360 387 363 390 
rect 360 390 363 393 
rect 360 393 363 396 
rect 360 396 363 399 
rect 360 399 363 402 
rect 360 402 363 405 
rect 360 405 363 408 
rect 360 408 363 411 
rect 360 411 363 414 
rect 360 414 363 417 
rect 360 417 363 420 
rect 360 420 363 423 
rect 360 423 363 426 
rect 360 426 363 429 
rect 360 429 363 432 
rect 360 432 363 435 
rect 360 435 363 438 
rect 360 438 363 441 
rect 360 441 363 444 
rect 360 444 363 447 
rect 360 447 363 450 
rect 360 450 363 453 
rect 360 453 363 456 
rect 360 456 363 459 
rect 360 459 363 462 
rect 360 462 363 465 
rect 360 465 363 468 
rect 360 468 363 471 
rect 360 471 363 474 
rect 360 474 363 477 
rect 360 477 363 480 
rect 360 480 363 483 
rect 360 483 363 486 
rect 360 486 363 489 
rect 360 489 363 492 
rect 360 492 363 495 
rect 360 495 363 498 
rect 360 498 363 501 
rect 360 501 363 504 
rect 360 504 363 507 
rect 360 507 363 510 
rect 363 0 366 3 
rect 363 3 366 6 
rect 363 6 366 9 
rect 363 9 366 12 
rect 363 12 366 15 
rect 363 15 366 18 
rect 363 18 366 21 
rect 363 21 366 24 
rect 363 24 366 27 
rect 363 27 366 30 
rect 363 30 366 33 
rect 363 33 366 36 
rect 363 36 366 39 
rect 363 39 366 42 
rect 363 42 366 45 
rect 363 45 366 48 
rect 363 48 366 51 
rect 363 51 366 54 
rect 363 54 366 57 
rect 363 57 366 60 
rect 363 60 366 63 
rect 363 63 366 66 
rect 363 66 366 69 
rect 363 69 366 72 
rect 363 72 366 75 
rect 363 75 366 78 
rect 363 78 366 81 
rect 363 81 366 84 
rect 363 84 366 87 
rect 363 87 366 90 
rect 363 90 366 93 
rect 363 93 366 96 
rect 363 96 366 99 
rect 363 99 366 102 
rect 363 102 366 105 
rect 363 105 366 108 
rect 363 108 366 111 
rect 363 111 366 114 
rect 363 114 366 117 
rect 363 117 366 120 
rect 363 120 366 123 
rect 363 123 366 126 
rect 363 126 366 129 
rect 363 129 366 132 
rect 363 132 366 135 
rect 363 135 366 138 
rect 363 138 366 141 
rect 363 141 366 144 
rect 363 144 366 147 
rect 363 147 366 150 
rect 363 150 366 153 
rect 363 153 366 156 
rect 363 156 366 159 
rect 363 159 366 162 
rect 363 162 366 165 
rect 363 165 366 168 
rect 363 168 366 171 
rect 363 171 366 174 
rect 363 174 366 177 
rect 363 177 366 180 
rect 363 180 366 183 
rect 363 183 366 186 
rect 363 186 366 189 
rect 363 189 366 192 
rect 363 192 366 195 
rect 363 195 366 198 
rect 363 198 366 201 
rect 363 201 366 204 
rect 363 204 366 207 
rect 363 207 366 210 
rect 363 210 366 213 
rect 363 213 366 216 
rect 363 216 366 219 
rect 363 219 366 222 
rect 363 222 366 225 
rect 363 225 366 228 
rect 363 228 366 231 
rect 363 231 366 234 
rect 363 234 366 237 
rect 363 237 366 240 
rect 363 240 366 243 
rect 363 243 366 246 
rect 363 246 366 249 
rect 363 249 366 252 
rect 363 252 366 255 
rect 363 255 366 258 
rect 363 258 366 261 
rect 363 261 366 264 
rect 363 264 366 267 
rect 363 267 366 270 
rect 363 270 366 273 
rect 363 273 366 276 
rect 363 276 366 279 
rect 363 279 366 282 
rect 363 282 366 285 
rect 363 285 366 288 
rect 363 288 366 291 
rect 363 291 366 294 
rect 363 294 366 297 
rect 363 297 366 300 
rect 363 300 366 303 
rect 363 303 366 306 
rect 363 306 366 309 
rect 363 309 366 312 
rect 363 312 366 315 
rect 363 315 366 318 
rect 363 318 366 321 
rect 363 321 366 324 
rect 363 324 366 327 
rect 363 327 366 330 
rect 363 330 366 333 
rect 363 333 366 336 
rect 363 336 366 339 
rect 363 339 366 342 
rect 363 342 366 345 
rect 363 345 366 348 
rect 363 348 366 351 
rect 363 351 366 354 
rect 363 354 366 357 
rect 363 357 366 360 
rect 363 360 366 363 
rect 363 363 366 366 
rect 363 366 366 369 
rect 363 369 366 372 
rect 363 372 366 375 
rect 363 375 366 378 
rect 363 378 366 381 
rect 363 381 366 384 
rect 363 384 366 387 
rect 363 387 366 390 
rect 363 390 366 393 
rect 363 393 366 396 
rect 363 396 366 399 
rect 363 399 366 402 
rect 363 402 366 405 
rect 363 405 366 408 
rect 363 408 366 411 
rect 363 411 366 414 
rect 363 414 366 417 
rect 363 417 366 420 
rect 363 420 366 423 
rect 363 423 366 426 
rect 363 426 366 429 
rect 363 429 366 432 
rect 363 432 366 435 
rect 363 435 366 438 
rect 363 438 366 441 
rect 363 441 366 444 
rect 363 444 366 447 
rect 363 447 366 450 
rect 363 450 366 453 
rect 363 453 366 456 
rect 363 456 366 459 
rect 363 459 366 462 
rect 363 462 366 465 
rect 363 465 366 468 
rect 363 468 366 471 
rect 363 471 366 474 
rect 363 474 366 477 
rect 363 477 366 480 
rect 363 480 366 483 
rect 363 483 366 486 
rect 363 486 366 489 
rect 363 489 366 492 
rect 363 492 366 495 
rect 363 495 366 498 
rect 363 498 366 501 
rect 363 501 366 504 
rect 363 504 366 507 
rect 363 507 366 510 
rect 366 0 369 3 
rect 366 3 369 6 
rect 366 6 369 9 
rect 366 9 369 12 
rect 366 12 369 15 
rect 366 15 369 18 
rect 366 18 369 21 
rect 366 21 369 24 
rect 366 24 369 27 
rect 366 27 369 30 
rect 366 30 369 33 
rect 366 33 369 36 
rect 366 36 369 39 
rect 366 39 369 42 
rect 366 42 369 45 
rect 366 45 369 48 
rect 366 48 369 51 
rect 366 51 369 54 
rect 366 54 369 57 
rect 366 57 369 60 
rect 366 60 369 63 
rect 366 63 369 66 
rect 366 66 369 69 
rect 366 69 369 72 
rect 366 72 369 75 
rect 366 75 369 78 
rect 366 78 369 81 
rect 366 81 369 84 
rect 366 84 369 87 
rect 366 87 369 90 
rect 366 90 369 93 
rect 366 93 369 96 
rect 366 96 369 99 
rect 366 99 369 102 
rect 366 102 369 105 
rect 366 105 369 108 
rect 366 108 369 111 
rect 366 111 369 114 
rect 366 114 369 117 
rect 366 117 369 120 
rect 366 120 369 123 
rect 366 123 369 126 
rect 366 126 369 129 
rect 366 129 369 132 
rect 366 132 369 135 
rect 366 135 369 138 
rect 366 138 369 141 
rect 366 141 369 144 
rect 366 144 369 147 
rect 366 147 369 150 
rect 366 150 369 153 
rect 366 153 369 156 
rect 366 156 369 159 
rect 366 159 369 162 
rect 366 162 369 165 
rect 366 165 369 168 
rect 366 168 369 171 
rect 366 171 369 174 
rect 366 174 369 177 
rect 366 177 369 180 
rect 366 180 369 183 
rect 366 183 369 186 
rect 366 186 369 189 
rect 366 189 369 192 
rect 366 192 369 195 
rect 366 195 369 198 
rect 366 198 369 201 
rect 366 201 369 204 
rect 366 204 369 207 
rect 366 207 369 210 
rect 366 210 369 213 
rect 366 213 369 216 
rect 366 216 369 219 
rect 366 219 369 222 
rect 366 222 369 225 
rect 366 225 369 228 
rect 366 228 369 231 
rect 366 231 369 234 
rect 366 234 369 237 
rect 366 237 369 240 
rect 366 240 369 243 
rect 366 243 369 246 
rect 366 246 369 249 
rect 366 249 369 252 
rect 366 252 369 255 
rect 366 255 369 258 
rect 366 258 369 261 
rect 366 261 369 264 
rect 366 264 369 267 
rect 366 267 369 270 
rect 366 270 369 273 
rect 366 273 369 276 
rect 366 276 369 279 
rect 366 279 369 282 
rect 366 282 369 285 
rect 366 285 369 288 
rect 366 288 369 291 
rect 366 291 369 294 
rect 366 294 369 297 
rect 366 297 369 300 
rect 366 300 369 303 
rect 366 303 369 306 
rect 366 306 369 309 
rect 366 309 369 312 
rect 366 312 369 315 
rect 366 315 369 318 
rect 366 318 369 321 
rect 366 321 369 324 
rect 366 324 369 327 
rect 366 327 369 330 
rect 366 330 369 333 
rect 366 333 369 336 
rect 366 336 369 339 
rect 366 339 369 342 
rect 366 342 369 345 
rect 366 345 369 348 
rect 366 348 369 351 
rect 366 351 369 354 
rect 366 354 369 357 
rect 366 357 369 360 
rect 366 360 369 363 
rect 366 363 369 366 
rect 366 366 369 369 
rect 366 369 369 372 
rect 366 372 369 375 
rect 366 375 369 378 
rect 366 378 369 381 
rect 366 381 369 384 
rect 366 384 369 387 
rect 366 387 369 390 
rect 366 390 369 393 
rect 366 393 369 396 
rect 366 396 369 399 
rect 366 399 369 402 
rect 366 402 369 405 
rect 366 405 369 408 
rect 366 408 369 411 
rect 366 411 369 414 
rect 366 414 369 417 
rect 366 417 369 420 
rect 366 420 369 423 
rect 366 423 369 426 
rect 366 426 369 429 
rect 366 429 369 432 
rect 366 432 369 435 
rect 366 435 369 438 
rect 366 438 369 441 
rect 366 441 369 444 
rect 366 444 369 447 
rect 366 447 369 450 
rect 366 450 369 453 
rect 366 453 369 456 
rect 366 456 369 459 
rect 366 459 369 462 
rect 366 462 369 465 
rect 366 465 369 468 
rect 366 468 369 471 
rect 366 471 369 474 
rect 366 474 369 477 
rect 366 477 369 480 
rect 366 480 369 483 
rect 366 483 369 486 
rect 366 486 369 489 
rect 366 489 369 492 
rect 366 492 369 495 
rect 366 495 369 498 
rect 366 498 369 501 
rect 366 501 369 504 
rect 366 504 369 507 
rect 366 507 369 510 
rect 369 0 372 3 
rect 369 3 372 6 
rect 369 6 372 9 
rect 369 9 372 12 
rect 369 12 372 15 
rect 369 15 372 18 
rect 369 18 372 21 
rect 369 21 372 24 
rect 369 24 372 27 
rect 369 27 372 30 
rect 369 30 372 33 
rect 369 33 372 36 
rect 369 36 372 39 
rect 369 39 372 42 
rect 369 42 372 45 
rect 369 45 372 48 
rect 369 48 372 51 
rect 369 51 372 54 
rect 369 54 372 57 
rect 369 57 372 60 
rect 369 60 372 63 
rect 369 63 372 66 
rect 369 66 372 69 
rect 369 69 372 72 
rect 369 72 372 75 
rect 369 75 372 78 
rect 369 78 372 81 
rect 369 81 372 84 
rect 369 84 372 87 
rect 369 87 372 90 
rect 369 90 372 93 
rect 369 93 372 96 
rect 369 96 372 99 
rect 369 99 372 102 
rect 369 102 372 105 
rect 369 105 372 108 
rect 369 108 372 111 
rect 369 111 372 114 
rect 369 114 372 117 
rect 369 117 372 120 
rect 369 120 372 123 
rect 369 123 372 126 
rect 369 126 372 129 
rect 369 129 372 132 
rect 369 132 372 135 
rect 369 135 372 138 
rect 369 138 372 141 
rect 369 141 372 144 
rect 369 144 372 147 
rect 369 147 372 150 
rect 369 150 372 153 
rect 369 153 372 156 
rect 369 156 372 159 
rect 369 159 372 162 
rect 369 162 372 165 
rect 369 165 372 168 
rect 369 168 372 171 
rect 369 171 372 174 
rect 369 174 372 177 
rect 369 177 372 180 
rect 369 180 372 183 
rect 369 183 372 186 
rect 369 186 372 189 
rect 369 189 372 192 
rect 369 192 372 195 
rect 369 195 372 198 
rect 369 198 372 201 
rect 369 201 372 204 
rect 369 204 372 207 
rect 369 207 372 210 
rect 369 210 372 213 
rect 369 213 372 216 
rect 369 216 372 219 
rect 369 219 372 222 
rect 369 222 372 225 
rect 369 225 372 228 
rect 369 228 372 231 
rect 369 231 372 234 
rect 369 234 372 237 
rect 369 237 372 240 
rect 369 240 372 243 
rect 369 243 372 246 
rect 369 246 372 249 
rect 369 249 372 252 
rect 369 252 372 255 
rect 369 255 372 258 
rect 369 258 372 261 
rect 369 261 372 264 
rect 369 264 372 267 
rect 369 267 372 270 
rect 369 270 372 273 
rect 369 273 372 276 
rect 369 276 372 279 
rect 369 279 372 282 
rect 369 282 372 285 
rect 369 285 372 288 
rect 369 288 372 291 
rect 369 291 372 294 
rect 369 294 372 297 
rect 369 297 372 300 
rect 369 300 372 303 
rect 369 303 372 306 
rect 369 306 372 309 
rect 369 309 372 312 
rect 369 312 372 315 
rect 369 315 372 318 
rect 369 318 372 321 
rect 369 321 372 324 
rect 369 324 372 327 
rect 369 327 372 330 
rect 369 330 372 333 
rect 369 333 372 336 
rect 369 336 372 339 
rect 369 339 372 342 
rect 369 342 372 345 
rect 369 345 372 348 
rect 369 348 372 351 
rect 369 351 372 354 
rect 369 354 372 357 
rect 369 357 372 360 
rect 369 360 372 363 
rect 369 363 372 366 
rect 369 366 372 369 
rect 369 369 372 372 
rect 369 372 372 375 
rect 369 375 372 378 
rect 369 378 372 381 
rect 369 381 372 384 
rect 369 384 372 387 
rect 369 387 372 390 
rect 369 390 372 393 
rect 369 393 372 396 
rect 369 396 372 399 
rect 369 399 372 402 
rect 369 402 372 405 
rect 369 405 372 408 
rect 369 408 372 411 
rect 369 411 372 414 
rect 369 414 372 417 
rect 369 417 372 420 
rect 369 420 372 423 
rect 369 423 372 426 
rect 369 426 372 429 
rect 369 429 372 432 
rect 369 432 372 435 
rect 369 435 372 438 
rect 369 438 372 441 
rect 369 441 372 444 
rect 369 444 372 447 
rect 369 447 372 450 
rect 369 450 372 453 
rect 369 453 372 456 
rect 369 456 372 459 
rect 369 459 372 462 
rect 369 462 372 465 
rect 369 465 372 468 
rect 369 468 372 471 
rect 369 471 372 474 
rect 369 474 372 477 
rect 369 477 372 480 
rect 369 480 372 483 
rect 369 483 372 486 
rect 369 486 372 489 
rect 369 489 372 492 
rect 369 492 372 495 
rect 369 495 372 498 
rect 369 498 372 501 
rect 369 501 372 504 
rect 369 504 372 507 
rect 369 507 372 510 
rect 372 0 375 3 
rect 372 3 375 6 
rect 372 6 375 9 
rect 372 9 375 12 
rect 372 12 375 15 
rect 372 15 375 18 
rect 372 18 375 21 
rect 372 21 375 24 
rect 372 24 375 27 
rect 372 27 375 30 
rect 372 30 375 33 
rect 372 33 375 36 
rect 372 36 375 39 
rect 372 39 375 42 
rect 372 42 375 45 
rect 372 45 375 48 
rect 372 48 375 51 
rect 372 51 375 54 
rect 372 54 375 57 
rect 372 57 375 60 
rect 372 60 375 63 
rect 372 63 375 66 
rect 372 66 375 69 
rect 372 69 375 72 
rect 372 72 375 75 
rect 372 75 375 78 
rect 372 78 375 81 
rect 372 81 375 84 
rect 372 84 375 87 
rect 372 87 375 90 
rect 372 90 375 93 
rect 372 93 375 96 
rect 372 96 375 99 
rect 372 99 375 102 
rect 372 102 375 105 
rect 372 105 375 108 
rect 372 108 375 111 
rect 372 111 375 114 
rect 372 114 375 117 
rect 372 117 375 120 
rect 372 120 375 123 
rect 372 123 375 126 
rect 372 126 375 129 
rect 372 129 375 132 
rect 372 132 375 135 
rect 372 135 375 138 
rect 372 138 375 141 
rect 372 141 375 144 
rect 372 144 375 147 
rect 372 147 375 150 
rect 372 150 375 153 
rect 372 153 375 156 
rect 372 156 375 159 
rect 372 159 375 162 
rect 372 162 375 165 
rect 372 165 375 168 
rect 372 168 375 171 
rect 372 171 375 174 
rect 372 174 375 177 
rect 372 177 375 180 
rect 372 180 375 183 
rect 372 183 375 186 
rect 372 186 375 189 
rect 372 189 375 192 
rect 372 192 375 195 
rect 372 195 375 198 
rect 372 198 375 201 
rect 372 201 375 204 
rect 372 204 375 207 
rect 372 207 375 210 
rect 372 210 375 213 
rect 372 213 375 216 
rect 372 216 375 219 
rect 372 219 375 222 
rect 372 222 375 225 
rect 372 225 375 228 
rect 372 228 375 231 
rect 372 231 375 234 
rect 372 234 375 237 
rect 372 237 375 240 
rect 372 240 375 243 
rect 372 243 375 246 
rect 372 246 375 249 
rect 372 249 375 252 
rect 372 252 375 255 
rect 372 255 375 258 
rect 372 258 375 261 
rect 372 261 375 264 
rect 372 264 375 267 
rect 372 267 375 270 
rect 372 270 375 273 
rect 372 273 375 276 
rect 372 276 375 279 
rect 372 279 375 282 
rect 372 282 375 285 
rect 372 285 375 288 
rect 372 288 375 291 
rect 372 291 375 294 
rect 372 294 375 297 
rect 372 297 375 300 
rect 372 300 375 303 
rect 372 303 375 306 
rect 372 306 375 309 
rect 372 309 375 312 
rect 372 312 375 315 
rect 372 315 375 318 
rect 372 318 375 321 
rect 372 321 375 324 
rect 372 324 375 327 
rect 372 327 375 330 
rect 372 330 375 333 
rect 372 333 375 336 
rect 372 336 375 339 
rect 372 339 375 342 
rect 372 342 375 345 
rect 372 345 375 348 
rect 372 348 375 351 
rect 372 351 375 354 
rect 372 354 375 357 
rect 372 357 375 360 
rect 372 360 375 363 
rect 372 363 375 366 
rect 372 366 375 369 
rect 372 369 375 372 
rect 372 372 375 375 
rect 372 375 375 378 
rect 372 378 375 381 
rect 372 381 375 384 
rect 372 384 375 387 
rect 372 387 375 390 
rect 372 390 375 393 
rect 372 393 375 396 
rect 372 396 375 399 
rect 372 399 375 402 
rect 372 402 375 405 
rect 372 405 375 408 
rect 372 408 375 411 
rect 372 411 375 414 
rect 372 414 375 417 
rect 372 417 375 420 
rect 372 420 375 423 
rect 372 423 375 426 
rect 372 426 375 429 
rect 372 429 375 432 
rect 372 432 375 435 
rect 372 435 375 438 
rect 372 438 375 441 
rect 372 441 375 444 
rect 372 444 375 447 
rect 372 447 375 450 
rect 372 450 375 453 
rect 372 453 375 456 
rect 372 456 375 459 
rect 372 459 375 462 
rect 372 462 375 465 
rect 372 465 375 468 
rect 372 468 375 471 
rect 372 471 375 474 
rect 372 474 375 477 
rect 372 477 375 480 
rect 372 480 375 483 
rect 372 483 375 486 
rect 372 486 375 489 
rect 372 489 375 492 
rect 372 492 375 495 
rect 372 495 375 498 
rect 372 498 375 501 
rect 372 501 375 504 
rect 372 504 375 507 
rect 372 507 375 510 
rect 375 0 378 3 
rect 375 3 378 6 
rect 375 6 378 9 
rect 375 9 378 12 
rect 375 12 378 15 
rect 375 15 378 18 
rect 375 18 378 21 
rect 375 21 378 24 
rect 375 24 378 27 
rect 375 27 378 30 
rect 375 30 378 33 
rect 375 33 378 36 
rect 375 36 378 39 
rect 375 39 378 42 
rect 375 42 378 45 
rect 375 45 378 48 
rect 375 48 378 51 
rect 375 51 378 54 
rect 375 54 378 57 
rect 375 57 378 60 
rect 375 60 378 63 
rect 375 63 378 66 
rect 375 66 378 69 
rect 375 69 378 72 
rect 375 72 378 75 
rect 375 75 378 78 
rect 375 78 378 81 
rect 375 81 378 84 
rect 375 84 378 87 
rect 375 87 378 90 
rect 375 90 378 93 
rect 375 93 378 96 
rect 375 96 378 99 
rect 375 99 378 102 
rect 375 102 378 105 
rect 375 105 378 108 
rect 375 108 378 111 
rect 375 111 378 114 
rect 375 114 378 117 
rect 375 117 378 120 
rect 375 120 378 123 
rect 375 123 378 126 
rect 375 126 378 129 
rect 375 129 378 132 
rect 375 132 378 135 
rect 375 135 378 138 
rect 375 138 378 141 
rect 375 141 378 144 
rect 375 144 378 147 
rect 375 147 378 150 
rect 375 150 378 153 
rect 375 153 378 156 
rect 375 156 378 159 
rect 375 159 378 162 
rect 375 162 378 165 
rect 375 165 378 168 
rect 375 168 378 171 
rect 375 171 378 174 
rect 375 174 378 177 
rect 375 177 378 180 
rect 375 180 378 183 
rect 375 183 378 186 
rect 375 186 378 189 
rect 375 189 378 192 
rect 375 192 378 195 
rect 375 195 378 198 
rect 375 198 378 201 
rect 375 201 378 204 
rect 375 204 378 207 
rect 375 207 378 210 
rect 375 210 378 213 
rect 375 213 378 216 
rect 375 216 378 219 
rect 375 219 378 222 
rect 375 222 378 225 
rect 375 225 378 228 
rect 375 228 378 231 
rect 375 231 378 234 
rect 375 234 378 237 
rect 375 237 378 240 
rect 375 240 378 243 
rect 375 243 378 246 
rect 375 246 378 249 
rect 375 249 378 252 
rect 375 252 378 255 
rect 375 255 378 258 
rect 375 258 378 261 
rect 375 261 378 264 
rect 375 264 378 267 
rect 375 267 378 270 
rect 375 270 378 273 
rect 375 273 378 276 
rect 375 276 378 279 
rect 375 279 378 282 
rect 375 282 378 285 
rect 375 285 378 288 
rect 375 288 378 291 
rect 375 291 378 294 
rect 375 294 378 297 
rect 375 297 378 300 
rect 375 300 378 303 
rect 375 303 378 306 
rect 375 306 378 309 
rect 375 309 378 312 
rect 375 312 378 315 
rect 375 315 378 318 
rect 375 318 378 321 
rect 375 321 378 324 
rect 375 324 378 327 
rect 375 327 378 330 
rect 375 330 378 333 
rect 375 333 378 336 
rect 375 336 378 339 
rect 375 339 378 342 
rect 375 342 378 345 
rect 375 345 378 348 
rect 375 348 378 351 
rect 375 351 378 354 
rect 375 354 378 357 
rect 375 357 378 360 
rect 375 360 378 363 
rect 375 363 378 366 
rect 375 366 378 369 
rect 375 369 378 372 
rect 375 372 378 375 
rect 375 375 378 378 
rect 375 378 378 381 
rect 375 381 378 384 
rect 375 384 378 387 
rect 375 387 378 390 
rect 375 390 378 393 
rect 375 393 378 396 
rect 375 396 378 399 
rect 375 399 378 402 
rect 375 402 378 405 
rect 375 405 378 408 
rect 375 408 378 411 
rect 375 411 378 414 
rect 375 414 378 417 
rect 375 417 378 420 
rect 375 420 378 423 
rect 375 423 378 426 
rect 375 426 378 429 
rect 375 429 378 432 
rect 375 432 378 435 
rect 375 435 378 438 
rect 375 438 378 441 
rect 375 441 378 444 
rect 375 444 378 447 
rect 375 447 378 450 
rect 375 450 378 453 
rect 375 453 378 456 
rect 375 456 378 459 
rect 375 459 378 462 
rect 375 462 378 465 
rect 375 465 378 468 
rect 375 468 378 471 
rect 375 471 378 474 
rect 375 474 378 477 
rect 375 477 378 480 
rect 375 480 378 483 
rect 375 483 378 486 
rect 375 486 378 489 
rect 375 489 378 492 
rect 375 492 378 495 
rect 375 495 378 498 
rect 375 498 378 501 
rect 375 501 378 504 
rect 375 504 378 507 
rect 375 507 378 510 
rect 378 0 381 3 
rect 378 3 381 6 
rect 378 6 381 9 
rect 378 9 381 12 
rect 378 12 381 15 
rect 378 15 381 18 
rect 378 18 381 21 
rect 378 21 381 24 
rect 378 24 381 27 
rect 378 27 381 30 
rect 378 30 381 33 
rect 378 33 381 36 
rect 378 36 381 39 
rect 378 39 381 42 
rect 378 42 381 45 
rect 378 45 381 48 
rect 378 48 381 51 
rect 378 51 381 54 
rect 378 54 381 57 
rect 378 57 381 60 
rect 378 60 381 63 
rect 378 63 381 66 
rect 378 66 381 69 
rect 378 69 381 72 
rect 378 72 381 75 
rect 378 75 381 78 
rect 378 78 381 81 
rect 378 81 381 84 
rect 378 84 381 87 
rect 378 87 381 90 
rect 378 90 381 93 
rect 378 93 381 96 
rect 378 96 381 99 
rect 378 99 381 102 
rect 378 102 381 105 
rect 378 105 381 108 
rect 378 108 381 111 
rect 378 111 381 114 
rect 378 114 381 117 
rect 378 117 381 120 
rect 378 120 381 123 
rect 378 123 381 126 
rect 378 126 381 129 
rect 378 129 381 132 
rect 378 132 381 135 
rect 378 135 381 138 
rect 378 138 381 141 
rect 378 141 381 144 
rect 378 144 381 147 
rect 378 147 381 150 
rect 378 150 381 153 
rect 378 153 381 156 
rect 378 156 381 159 
rect 378 159 381 162 
rect 378 162 381 165 
rect 378 165 381 168 
rect 378 168 381 171 
rect 378 171 381 174 
rect 378 174 381 177 
rect 378 177 381 180 
rect 378 180 381 183 
rect 378 183 381 186 
rect 378 186 381 189 
rect 378 189 381 192 
rect 378 192 381 195 
rect 378 195 381 198 
rect 378 198 381 201 
rect 378 201 381 204 
rect 378 204 381 207 
rect 378 207 381 210 
rect 378 210 381 213 
rect 378 213 381 216 
rect 378 216 381 219 
rect 378 219 381 222 
rect 378 222 381 225 
rect 378 225 381 228 
rect 378 228 381 231 
rect 378 231 381 234 
rect 378 234 381 237 
rect 378 237 381 240 
rect 378 240 381 243 
rect 378 243 381 246 
rect 378 246 381 249 
rect 378 249 381 252 
rect 378 252 381 255 
rect 378 255 381 258 
rect 378 258 381 261 
rect 378 261 381 264 
rect 378 264 381 267 
rect 378 267 381 270 
rect 378 270 381 273 
rect 378 273 381 276 
rect 378 276 381 279 
rect 378 279 381 282 
rect 378 282 381 285 
rect 378 285 381 288 
rect 378 288 381 291 
rect 378 291 381 294 
rect 378 294 381 297 
rect 378 297 381 300 
rect 378 300 381 303 
rect 378 303 381 306 
rect 378 306 381 309 
rect 378 309 381 312 
rect 378 312 381 315 
rect 378 315 381 318 
rect 378 318 381 321 
rect 378 321 381 324 
rect 378 324 381 327 
rect 378 327 381 330 
rect 378 330 381 333 
rect 378 333 381 336 
rect 378 336 381 339 
rect 378 339 381 342 
rect 378 342 381 345 
rect 378 345 381 348 
rect 378 348 381 351 
rect 378 351 381 354 
rect 378 354 381 357 
rect 378 357 381 360 
rect 378 360 381 363 
rect 378 363 381 366 
rect 378 366 381 369 
rect 378 369 381 372 
rect 378 372 381 375 
rect 378 375 381 378 
rect 378 378 381 381 
rect 378 381 381 384 
rect 378 384 381 387 
rect 378 387 381 390 
rect 378 390 381 393 
rect 378 393 381 396 
rect 378 396 381 399 
rect 378 399 381 402 
rect 378 402 381 405 
rect 378 405 381 408 
rect 378 408 381 411 
rect 378 411 381 414 
rect 378 414 381 417 
rect 378 417 381 420 
rect 378 420 381 423 
rect 378 423 381 426 
rect 378 426 381 429 
rect 378 429 381 432 
rect 378 432 381 435 
rect 378 435 381 438 
rect 378 438 381 441 
rect 378 441 381 444 
rect 378 444 381 447 
rect 378 447 381 450 
rect 378 450 381 453 
rect 378 453 381 456 
rect 378 456 381 459 
rect 378 459 381 462 
rect 378 462 381 465 
rect 378 465 381 468 
rect 378 468 381 471 
rect 378 471 381 474 
rect 378 474 381 477 
rect 378 477 381 480 
rect 378 480 381 483 
rect 378 483 381 486 
rect 378 486 381 489 
rect 378 489 381 492 
rect 378 492 381 495 
rect 378 495 381 498 
rect 378 498 381 501 
rect 378 501 381 504 
rect 378 504 381 507 
rect 378 507 381 510 
rect 381 0 384 3 
rect 381 3 384 6 
rect 381 6 384 9 
rect 381 9 384 12 
rect 381 12 384 15 
rect 381 15 384 18 
rect 381 18 384 21 
rect 381 21 384 24 
rect 381 24 384 27 
rect 381 27 384 30 
rect 381 30 384 33 
rect 381 33 384 36 
rect 381 36 384 39 
rect 381 39 384 42 
rect 381 42 384 45 
rect 381 45 384 48 
rect 381 48 384 51 
rect 381 51 384 54 
rect 381 54 384 57 
rect 381 57 384 60 
rect 381 60 384 63 
rect 381 63 384 66 
rect 381 66 384 69 
rect 381 69 384 72 
rect 381 72 384 75 
rect 381 75 384 78 
rect 381 78 384 81 
rect 381 81 384 84 
rect 381 84 384 87 
rect 381 87 384 90 
rect 381 90 384 93 
rect 381 93 384 96 
rect 381 96 384 99 
rect 381 99 384 102 
rect 381 102 384 105 
rect 381 105 384 108 
rect 381 108 384 111 
rect 381 111 384 114 
rect 381 114 384 117 
rect 381 117 384 120 
rect 381 120 384 123 
rect 381 123 384 126 
rect 381 126 384 129 
rect 381 129 384 132 
rect 381 132 384 135 
rect 381 135 384 138 
rect 381 138 384 141 
rect 381 141 384 144 
rect 381 144 384 147 
rect 381 147 384 150 
rect 381 150 384 153 
rect 381 153 384 156 
rect 381 156 384 159 
rect 381 159 384 162 
rect 381 162 384 165 
rect 381 165 384 168 
rect 381 168 384 171 
rect 381 171 384 174 
rect 381 174 384 177 
rect 381 177 384 180 
rect 381 180 384 183 
rect 381 183 384 186 
rect 381 186 384 189 
rect 381 189 384 192 
rect 381 192 384 195 
rect 381 195 384 198 
rect 381 198 384 201 
rect 381 201 384 204 
rect 381 204 384 207 
rect 381 207 384 210 
rect 381 210 384 213 
rect 381 213 384 216 
rect 381 216 384 219 
rect 381 219 384 222 
rect 381 222 384 225 
rect 381 225 384 228 
rect 381 228 384 231 
rect 381 231 384 234 
rect 381 234 384 237 
rect 381 237 384 240 
rect 381 240 384 243 
rect 381 243 384 246 
rect 381 246 384 249 
rect 381 249 384 252 
rect 381 252 384 255 
rect 381 255 384 258 
rect 381 258 384 261 
rect 381 261 384 264 
rect 381 264 384 267 
rect 381 267 384 270 
rect 381 270 384 273 
rect 381 273 384 276 
rect 381 276 384 279 
rect 381 279 384 282 
rect 381 282 384 285 
rect 381 285 384 288 
rect 381 288 384 291 
rect 381 291 384 294 
rect 381 294 384 297 
rect 381 297 384 300 
rect 381 300 384 303 
rect 381 303 384 306 
rect 381 306 384 309 
rect 381 309 384 312 
rect 381 312 384 315 
rect 381 315 384 318 
rect 381 318 384 321 
rect 381 321 384 324 
rect 381 324 384 327 
rect 381 327 384 330 
rect 381 330 384 333 
rect 381 333 384 336 
rect 381 336 384 339 
rect 381 339 384 342 
rect 381 342 384 345 
rect 381 345 384 348 
rect 381 348 384 351 
rect 381 351 384 354 
rect 381 354 384 357 
rect 381 357 384 360 
rect 381 360 384 363 
rect 381 363 384 366 
rect 381 366 384 369 
rect 381 369 384 372 
rect 381 372 384 375 
rect 381 375 384 378 
rect 381 378 384 381 
rect 381 381 384 384 
rect 381 384 384 387 
rect 381 387 384 390 
rect 381 390 384 393 
rect 381 393 384 396 
rect 381 396 384 399 
rect 381 399 384 402 
rect 381 402 384 405 
rect 381 405 384 408 
rect 381 408 384 411 
rect 381 411 384 414 
rect 381 414 384 417 
rect 381 417 384 420 
rect 381 420 384 423 
rect 381 423 384 426 
rect 381 426 384 429 
rect 381 429 384 432 
rect 381 432 384 435 
rect 381 435 384 438 
rect 381 438 384 441 
rect 381 441 384 444 
rect 381 444 384 447 
rect 381 447 384 450 
rect 381 450 384 453 
rect 381 453 384 456 
rect 381 456 384 459 
rect 381 459 384 462 
rect 381 462 384 465 
rect 381 465 384 468 
rect 381 468 384 471 
rect 381 471 384 474 
rect 381 474 384 477 
rect 381 477 384 480 
rect 381 480 384 483 
rect 381 483 384 486 
rect 381 486 384 489 
rect 381 489 384 492 
rect 381 492 384 495 
rect 381 495 384 498 
rect 381 498 384 501 
rect 381 501 384 504 
rect 381 504 384 507 
rect 381 507 384 510 
rect 384 0 387 3 
rect 384 3 387 6 
rect 384 6 387 9 
rect 384 9 387 12 
rect 384 12 387 15 
rect 384 15 387 18 
rect 384 18 387 21 
rect 384 21 387 24 
rect 384 24 387 27 
rect 384 27 387 30 
rect 384 30 387 33 
rect 384 33 387 36 
rect 384 36 387 39 
rect 384 39 387 42 
rect 384 42 387 45 
rect 384 45 387 48 
rect 384 48 387 51 
rect 384 51 387 54 
rect 384 54 387 57 
rect 384 57 387 60 
rect 384 60 387 63 
rect 384 63 387 66 
rect 384 66 387 69 
rect 384 69 387 72 
rect 384 72 387 75 
rect 384 75 387 78 
rect 384 78 387 81 
rect 384 81 387 84 
rect 384 84 387 87 
rect 384 87 387 90 
rect 384 90 387 93 
rect 384 93 387 96 
rect 384 96 387 99 
rect 384 99 387 102 
rect 384 102 387 105 
rect 384 105 387 108 
rect 384 108 387 111 
rect 384 111 387 114 
rect 384 114 387 117 
rect 384 117 387 120 
rect 384 120 387 123 
rect 384 123 387 126 
rect 384 126 387 129 
rect 384 129 387 132 
rect 384 132 387 135 
rect 384 135 387 138 
rect 384 138 387 141 
rect 384 141 387 144 
rect 384 144 387 147 
rect 384 147 387 150 
rect 384 150 387 153 
rect 384 153 387 156 
rect 384 156 387 159 
rect 384 159 387 162 
rect 384 162 387 165 
rect 384 165 387 168 
rect 384 168 387 171 
rect 384 171 387 174 
rect 384 174 387 177 
rect 384 177 387 180 
rect 384 180 387 183 
rect 384 183 387 186 
rect 384 186 387 189 
rect 384 189 387 192 
rect 384 192 387 195 
rect 384 195 387 198 
rect 384 198 387 201 
rect 384 201 387 204 
rect 384 204 387 207 
rect 384 207 387 210 
rect 384 210 387 213 
rect 384 213 387 216 
rect 384 216 387 219 
rect 384 219 387 222 
rect 384 222 387 225 
rect 384 225 387 228 
rect 384 228 387 231 
rect 384 231 387 234 
rect 384 234 387 237 
rect 384 237 387 240 
rect 384 240 387 243 
rect 384 243 387 246 
rect 384 246 387 249 
rect 384 249 387 252 
rect 384 252 387 255 
rect 384 255 387 258 
rect 384 258 387 261 
rect 384 261 387 264 
rect 384 264 387 267 
rect 384 267 387 270 
rect 384 270 387 273 
rect 384 273 387 276 
rect 384 276 387 279 
rect 384 279 387 282 
rect 384 282 387 285 
rect 384 285 387 288 
rect 384 288 387 291 
rect 384 291 387 294 
rect 384 294 387 297 
rect 384 297 387 300 
rect 384 300 387 303 
rect 384 303 387 306 
rect 384 306 387 309 
rect 384 309 387 312 
rect 384 312 387 315 
rect 384 315 387 318 
rect 384 318 387 321 
rect 384 321 387 324 
rect 384 324 387 327 
rect 384 327 387 330 
rect 384 330 387 333 
rect 384 333 387 336 
rect 384 336 387 339 
rect 384 339 387 342 
rect 384 342 387 345 
rect 384 345 387 348 
rect 384 348 387 351 
rect 384 351 387 354 
rect 384 354 387 357 
rect 384 357 387 360 
rect 384 360 387 363 
rect 384 363 387 366 
rect 384 366 387 369 
rect 384 369 387 372 
rect 384 372 387 375 
rect 384 375 387 378 
rect 384 378 387 381 
rect 384 381 387 384 
rect 384 384 387 387 
rect 384 387 387 390 
rect 384 390 387 393 
rect 384 393 387 396 
rect 384 396 387 399 
rect 384 399 387 402 
rect 384 402 387 405 
rect 384 405 387 408 
rect 384 408 387 411 
rect 384 411 387 414 
rect 384 414 387 417 
rect 384 417 387 420 
rect 384 420 387 423 
rect 384 423 387 426 
rect 384 426 387 429 
rect 384 429 387 432 
rect 384 432 387 435 
rect 384 435 387 438 
rect 384 438 387 441 
rect 384 441 387 444 
rect 384 444 387 447 
rect 384 447 387 450 
rect 384 450 387 453 
rect 384 453 387 456 
rect 384 456 387 459 
rect 384 459 387 462 
rect 384 462 387 465 
rect 384 465 387 468 
rect 384 468 387 471 
rect 384 471 387 474 
rect 384 474 387 477 
rect 384 477 387 480 
rect 384 480 387 483 
rect 384 483 387 486 
rect 384 486 387 489 
rect 384 489 387 492 
rect 384 492 387 495 
rect 384 495 387 498 
rect 384 498 387 501 
rect 384 501 387 504 
rect 384 504 387 507 
rect 384 507 387 510 
rect 387 0 390 3 
rect 387 3 390 6 
rect 387 6 390 9 
rect 387 9 390 12 
rect 387 12 390 15 
rect 387 15 390 18 
rect 387 18 390 21 
rect 387 21 390 24 
rect 387 24 390 27 
rect 387 27 390 30 
rect 387 30 390 33 
rect 387 33 390 36 
rect 387 36 390 39 
rect 387 39 390 42 
rect 387 42 390 45 
rect 387 45 390 48 
rect 387 48 390 51 
rect 387 51 390 54 
rect 387 54 390 57 
rect 387 57 390 60 
rect 387 60 390 63 
rect 387 63 390 66 
rect 387 66 390 69 
rect 387 69 390 72 
rect 387 72 390 75 
rect 387 75 390 78 
rect 387 78 390 81 
rect 387 81 390 84 
rect 387 84 390 87 
rect 387 87 390 90 
rect 387 90 390 93 
rect 387 93 390 96 
rect 387 96 390 99 
rect 387 99 390 102 
rect 387 102 390 105 
rect 387 105 390 108 
rect 387 108 390 111 
rect 387 111 390 114 
rect 387 114 390 117 
rect 387 117 390 120 
rect 387 120 390 123 
rect 387 123 390 126 
rect 387 126 390 129 
rect 387 129 390 132 
rect 387 132 390 135 
rect 387 135 390 138 
rect 387 138 390 141 
rect 387 141 390 144 
rect 387 144 390 147 
rect 387 147 390 150 
rect 387 150 390 153 
rect 387 153 390 156 
rect 387 156 390 159 
rect 387 159 390 162 
rect 387 162 390 165 
rect 387 165 390 168 
rect 387 168 390 171 
rect 387 171 390 174 
rect 387 174 390 177 
rect 387 177 390 180 
rect 387 180 390 183 
rect 387 183 390 186 
rect 387 186 390 189 
rect 387 189 390 192 
rect 387 192 390 195 
rect 387 195 390 198 
rect 387 198 390 201 
rect 387 201 390 204 
rect 387 204 390 207 
rect 387 207 390 210 
rect 387 210 390 213 
rect 387 213 390 216 
rect 387 216 390 219 
rect 387 219 390 222 
rect 387 222 390 225 
rect 387 225 390 228 
rect 387 228 390 231 
rect 387 231 390 234 
rect 387 234 390 237 
rect 387 237 390 240 
rect 387 240 390 243 
rect 387 243 390 246 
rect 387 246 390 249 
rect 387 249 390 252 
rect 387 252 390 255 
rect 387 255 390 258 
rect 387 258 390 261 
rect 387 261 390 264 
rect 387 264 390 267 
rect 387 267 390 270 
rect 387 270 390 273 
rect 387 273 390 276 
rect 387 276 390 279 
rect 387 279 390 282 
rect 387 282 390 285 
rect 387 285 390 288 
rect 387 288 390 291 
rect 387 291 390 294 
rect 387 294 390 297 
rect 387 297 390 300 
rect 387 300 390 303 
rect 387 303 390 306 
rect 387 306 390 309 
rect 387 309 390 312 
rect 387 312 390 315 
rect 387 315 390 318 
rect 387 318 390 321 
rect 387 321 390 324 
rect 387 324 390 327 
rect 387 327 390 330 
rect 387 330 390 333 
rect 387 333 390 336 
rect 387 336 390 339 
rect 387 339 390 342 
rect 387 342 390 345 
rect 387 345 390 348 
rect 387 348 390 351 
rect 387 351 390 354 
rect 387 354 390 357 
rect 387 357 390 360 
rect 387 360 390 363 
rect 387 363 390 366 
rect 387 366 390 369 
rect 387 369 390 372 
rect 387 372 390 375 
rect 387 375 390 378 
rect 387 378 390 381 
rect 387 381 390 384 
rect 387 384 390 387 
rect 387 387 390 390 
rect 387 390 390 393 
rect 387 393 390 396 
rect 387 396 390 399 
rect 387 399 390 402 
rect 387 402 390 405 
rect 387 405 390 408 
rect 387 408 390 411 
rect 387 411 390 414 
rect 387 414 390 417 
rect 387 417 390 420 
rect 387 420 390 423 
rect 387 423 390 426 
rect 387 426 390 429 
rect 387 429 390 432 
rect 387 432 390 435 
rect 387 435 390 438 
rect 387 438 390 441 
rect 387 441 390 444 
rect 387 444 390 447 
rect 387 447 390 450 
rect 387 450 390 453 
rect 387 453 390 456 
rect 387 456 390 459 
rect 387 459 390 462 
rect 387 462 390 465 
rect 387 465 390 468 
rect 387 468 390 471 
rect 387 471 390 474 
rect 387 474 390 477 
rect 387 477 390 480 
rect 387 480 390 483 
rect 387 483 390 486 
rect 387 486 390 489 
rect 387 489 390 492 
rect 387 492 390 495 
rect 387 495 390 498 
rect 387 498 390 501 
rect 387 501 390 504 
rect 387 504 390 507 
rect 387 507 390 510 
rect 390 0 393 3 
rect 390 3 393 6 
rect 390 6 393 9 
rect 390 9 393 12 
rect 390 12 393 15 
rect 390 15 393 18 
rect 390 18 393 21 
rect 390 21 393 24 
rect 390 24 393 27 
rect 390 27 393 30 
rect 390 30 393 33 
rect 390 33 393 36 
rect 390 36 393 39 
rect 390 39 393 42 
rect 390 42 393 45 
rect 390 45 393 48 
rect 390 48 393 51 
rect 390 51 393 54 
rect 390 54 393 57 
rect 390 57 393 60 
rect 390 60 393 63 
rect 390 63 393 66 
rect 390 66 393 69 
rect 390 69 393 72 
rect 390 72 393 75 
rect 390 75 393 78 
rect 390 78 393 81 
rect 390 81 393 84 
rect 390 84 393 87 
rect 390 87 393 90 
rect 390 90 393 93 
rect 390 93 393 96 
rect 390 96 393 99 
rect 390 99 393 102 
rect 390 102 393 105 
rect 390 105 393 108 
rect 390 108 393 111 
rect 390 111 393 114 
rect 390 114 393 117 
rect 390 117 393 120 
rect 390 120 393 123 
rect 390 123 393 126 
rect 390 126 393 129 
rect 390 129 393 132 
rect 390 132 393 135 
rect 390 135 393 138 
rect 390 138 393 141 
rect 390 141 393 144 
rect 390 144 393 147 
rect 390 147 393 150 
rect 390 150 393 153 
rect 390 153 393 156 
rect 390 156 393 159 
rect 390 159 393 162 
rect 390 162 393 165 
rect 390 165 393 168 
rect 390 168 393 171 
rect 390 171 393 174 
rect 390 174 393 177 
rect 390 177 393 180 
rect 390 180 393 183 
rect 390 183 393 186 
rect 390 186 393 189 
rect 390 189 393 192 
rect 390 192 393 195 
rect 390 195 393 198 
rect 390 198 393 201 
rect 390 201 393 204 
rect 390 204 393 207 
rect 390 207 393 210 
rect 390 210 393 213 
rect 390 213 393 216 
rect 390 216 393 219 
rect 390 219 393 222 
rect 390 222 393 225 
rect 390 225 393 228 
rect 390 228 393 231 
rect 390 231 393 234 
rect 390 234 393 237 
rect 390 237 393 240 
rect 390 240 393 243 
rect 390 243 393 246 
rect 390 246 393 249 
rect 390 249 393 252 
rect 390 252 393 255 
rect 390 255 393 258 
rect 390 258 393 261 
rect 390 261 393 264 
rect 390 264 393 267 
rect 390 267 393 270 
rect 390 270 393 273 
rect 390 273 393 276 
rect 390 276 393 279 
rect 390 279 393 282 
rect 390 282 393 285 
rect 390 285 393 288 
rect 390 288 393 291 
rect 390 291 393 294 
rect 390 294 393 297 
rect 390 297 393 300 
rect 390 300 393 303 
rect 390 303 393 306 
rect 390 306 393 309 
rect 390 309 393 312 
rect 390 312 393 315 
rect 390 315 393 318 
rect 390 318 393 321 
rect 390 321 393 324 
rect 390 324 393 327 
rect 390 327 393 330 
rect 390 330 393 333 
rect 390 333 393 336 
rect 390 336 393 339 
rect 390 339 393 342 
rect 390 342 393 345 
rect 390 345 393 348 
rect 390 348 393 351 
rect 390 351 393 354 
rect 390 354 393 357 
rect 390 357 393 360 
rect 390 360 393 363 
rect 390 363 393 366 
rect 390 366 393 369 
rect 390 369 393 372 
rect 390 372 393 375 
rect 390 375 393 378 
rect 390 378 393 381 
rect 390 381 393 384 
rect 390 384 393 387 
rect 390 387 393 390 
rect 390 390 393 393 
rect 390 393 393 396 
rect 390 396 393 399 
rect 390 399 393 402 
rect 390 402 393 405 
rect 390 405 393 408 
rect 390 408 393 411 
rect 390 411 393 414 
rect 390 414 393 417 
rect 390 417 393 420 
rect 390 420 393 423 
rect 390 423 393 426 
rect 390 426 393 429 
rect 390 429 393 432 
rect 390 432 393 435 
rect 390 435 393 438 
rect 390 438 393 441 
rect 390 441 393 444 
rect 390 444 393 447 
rect 390 447 393 450 
rect 390 450 393 453 
rect 390 453 393 456 
rect 390 456 393 459 
rect 390 459 393 462 
rect 390 462 393 465 
rect 390 465 393 468 
rect 390 468 393 471 
rect 390 471 393 474 
rect 390 474 393 477 
rect 390 477 393 480 
rect 390 480 393 483 
rect 390 483 393 486 
rect 390 486 393 489 
rect 390 489 393 492 
rect 390 492 393 495 
rect 390 495 393 498 
rect 390 498 393 501 
rect 390 501 393 504 
rect 390 504 393 507 
rect 390 507 393 510 
rect 393 0 396 3 
rect 393 3 396 6 
rect 393 6 396 9 
rect 393 9 396 12 
rect 393 12 396 15 
rect 393 15 396 18 
rect 393 18 396 21 
rect 393 21 396 24 
rect 393 24 396 27 
rect 393 27 396 30 
rect 393 30 396 33 
rect 393 33 396 36 
rect 393 36 396 39 
rect 393 39 396 42 
rect 393 42 396 45 
rect 393 45 396 48 
rect 393 48 396 51 
rect 393 51 396 54 
rect 393 54 396 57 
rect 393 57 396 60 
rect 393 60 396 63 
rect 393 63 396 66 
rect 393 66 396 69 
rect 393 69 396 72 
rect 393 72 396 75 
rect 393 75 396 78 
rect 393 78 396 81 
rect 393 81 396 84 
rect 393 84 396 87 
rect 393 87 396 90 
rect 393 90 396 93 
rect 393 93 396 96 
rect 393 96 396 99 
rect 393 99 396 102 
rect 393 102 396 105 
rect 393 105 396 108 
rect 393 108 396 111 
rect 393 111 396 114 
rect 393 114 396 117 
rect 393 117 396 120 
rect 393 120 396 123 
rect 393 123 396 126 
rect 393 126 396 129 
rect 393 129 396 132 
rect 393 132 396 135 
rect 393 135 396 138 
rect 393 138 396 141 
rect 393 141 396 144 
rect 393 144 396 147 
rect 393 147 396 150 
rect 393 150 396 153 
rect 393 153 396 156 
rect 393 156 396 159 
rect 393 159 396 162 
rect 393 162 396 165 
rect 393 165 396 168 
rect 393 168 396 171 
rect 393 171 396 174 
rect 393 174 396 177 
rect 393 177 396 180 
rect 393 180 396 183 
rect 393 183 396 186 
rect 393 186 396 189 
rect 393 189 396 192 
rect 393 192 396 195 
rect 393 195 396 198 
rect 393 198 396 201 
rect 393 201 396 204 
rect 393 204 396 207 
rect 393 207 396 210 
rect 393 210 396 213 
rect 393 213 396 216 
rect 393 216 396 219 
rect 393 219 396 222 
rect 393 222 396 225 
rect 393 225 396 228 
rect 393 228 396 231 
rect 393 231 396 234 
rect 393 234 396 237 
rect 393 237 396 240 
rect 393 240 396 243 
rect 393 243 396 246 
rect 393 246 396 249 
rect 393 249 396 252 
rect 393 252 396 255 
rect 393 255 396 258 
rect 393 258 396 261 
rect 393 261 396 264 
rect 393 264 396 267 
rect 393 267 396 270 
rect 393 270 396 273 
rect 393 273 396 276 
rect 393 276 396 279 
rect 393 279 396 282 
rect 393 282 396 285 
rect 393 285 396 288 
rect 393 288 396 291 
rect 393 291 396 294 
rect 393 294 396 297 
rect 393 297 396 300 
rect 393 300 396 303 
rect 393 303 396 306 
rect 393 306 396 309 
rect 393 309 396 312 
rect 393 312 396 315 
rect 393 315 396 318 
rect 393 318 396 321 
rect 393 321 396 324 
rect 393 324 396 327 
rect 393 327 396 330 
rect 393 330 396 333 
rect 393 333 396 336 
rect 393 336 396 339 
rect 393 339 396 342 
rect 393 342 396 345 
rect 393 345 396 348 
rect 393 348 396 351 
rect 393 351 396 354 
rect 393 354 396 357 
rect 393 357 396 360 
rect 393 360 396 363 
rect 393 363 396 366 
rect 393 366 396 369 
rect 393 369 396 372 
rect 393 372 396 375 
rect 393 375 396 378 
rect 393 378 396 381 
rect 393 381 396 384 
rect 393 384 396 387 
rect 393 387 396 390 
rect 393 390 396 393 
rect 393 393 396 396 
rect 393 396 396 399 
rect 393 399 396 402 
rect 393 402 396 405 
rect 393 405 396 408 
rect 393 408 396 411 
rect 393 411 396 414 
rect 393 414 396 417 
rect 393 417 396 420 
rect 393 420 396 423 
rect 393 423 396 426 
rect 393 426 396 429 
rect 393 429 396 432 
rect 393 432 396 435 
rect 393 435 396 438 
rect 393 438 396 441 
rect 393 441 396 444 
rect 393 444 396 447 
rect 393 447 396 450 
rect 393 450 396 453 
rect 393 453 396 456 
rect 393 456 396 459 
rect 393 459 396 462 
rect 393 462 396 465 
rect 393 465 396 468 
rect 393 468 396 471 
rect 393 471 396 474 
rect 393 474 396 477 
rect 393 477 396 480 
rect 393 480 396 483 
rect 393 483 396 486 
rect 393 486 396 489 
rect 393 489 396 492 
rect 393 492 396 495 
rect 393 495 396 498 
rect 393 498 396 501 
rect 393 501 396 504 
rect 393 504 396 507 
rect 393 507 396 510 
rect 396 0 399 3 
rect 396 3 399 6 
rect 396 6 399 9 
rect 396 9 399 12 
rect 396 12 399 15 
rect 396 15 399 18 
rect 396 18 399 21 
rect 396 21 399 24 
rect 396 24 399 27 
rect 396 27 399 30 
rect 396 30 399 33 
rect 396 33 399 36 
rect 396 36 399 39 
rect 396 39 399 42 
rect 396 42 399 45 
rect 396 45 399 48 
rect 396 48 399 51 
rect 396 51 399 54 
rect 396 54 399 57 
rect 396 57 399 60 
rect 396 60 399 63 
rect 396 63 399 66 
rect 396 66 399 69 
rect 396 69 399 72 
rect 396 72 399 75 
rect 396 75 399 78 
rect 396 78 399 81 
rect 396 81 399 84 
rect 396 84 399 87 
rect 396 87 399 90 
rect 396 90 399 93 
rect 396 93 399 96 
rect 396 96 399 99 
rect 396 99 399 102 
rect 396 102 399 105 
rect 396 105 399 108 
rect 396 108 399 111 
rect 396 111 399 114 
rect 396 114 399 117 
rect 396 117 399 120 
rect 396 120 399 123 
rect 396 123 399 126 
rect 396 126 399 129 
rect 396 129 399 132 
rect 396 132 399 135 
rect 396 135 399 138 
rect 396 138 399 141 
rect 396 141 399 144 
rect 396 144 399 147 
rect 396 147 399 150 
rect 396 150 399 153 
rect 396 153 399 156 
rect 396 156 399 159 
rect 396 159 399 162 
rect 396 162 399 165 
rect 396 165 399 168 
rect 396 168 399 171 
rect 396 171 399 174 
rect 396 174 399 177 
rect 396 177 399 180 
rect 396 180 399 183 
rect 396 183 399 186 
rect 396 186 399 189 
rect 396 189 399 192 
rect 396 192 399 195 
rect 396 195 399 198 
rect 396 198 399 201 
rect 396 201 399 204 
rect 396 204 399 207 
rect 396 207 399 210 
rect 396 210 399 213 
rect 396 213 399 216 
rect 396 216 399 219 
rect 396 219 399 222 
rect 396 222 399 225 
rect 396 225 399 228 
rect 396 228 399 231 
rect 396 231 399 234 
rect 396 234 399 237 
rect 396 237 399 240 
rect 396 240 399 243 
rect 396 243 399 246 
rect 396 246 399 249 
rect 396 249 399 252 
rect 396 252 399 255 
rect 396 255 399 258 
rect 396 258 399 261 
rect 396 261 399 264 
rect 396 264 399 267 
rect 396 267 399 270 
rect 396 270 399 273 
rect 396 273 399 276 
rect 396 276 399 279 
rect 396 279 399 282 
rect 396 282 399 285 
rect 396 285 399 288 
rect 396 288 399 291 
rect 396 291 399 294 
rect 396 294 399 297 
rect 396 297 399 300 
rect 396 300 399 303 
rect 396 303 399 306 
rect 396 306 399 309 
rect 396 309 399 312 
rect 396 312 399 315 
rect 396 315 399 318 
rect 396 318 399 321 
rect 396 321 399 324 
rect 396 324 399 327 
rect 396 327 399 330 
rect 396 330 399 333 
rect 396 333 399 336 
rect 396 336 399 339 
rect 396 339 399 342 
rect 396 342 399 345 
rect 396 345 399 348 
rect 396 348 399 351 
rect 396 351 399 354 
rect 396 354 399 357 
rect 396 357 399 360 
rect 396 360 399 363 
rect 396 363 399 366 
rect 396 366 399 369 
rect 396 369 399 372 
rect 396 372 399 375 
rect 396 375 399 378 
rect 396 378 399 381 
rect 396 381 399 384 
rect 396 384 399 387 
rect 396 387 399 390 
rect 396 390 399 393 
rect 396 393 399 396 
rect 396 396 399 399 
rect 396 399 399 402 
rect 396 402 399 405 
rect 396 405 399 408 
rect 396 408 399 411 
rect 396 411 399 414 
rect 396 414 399 417 
rect 396 417 399 420 
rect 396 420 399 423 
rect 396 423 399 426 
rect 396 426 399 429 
rect 396 429 399 432 
rect 396 432 399 435 
rect 396 435 399 438 
rect 396 438 399 441 
rect 396 441 399 444 
rect 396 444 399 447 
rect 396 447 399 450 
rect 396 450 399 453 
rect 396 453 399 456 
rect 396 456 399 459 
rect 396 459 399 462 
rect 396 462 399 465 
rect 396 465 399 468 
rect 396 468 399 471 
rect 396 471 399 474 
rect 396 474 399 477 
rect 396 477 399 480 
rect 396 480 399 483 
rect 396 483 399 486 
rect 396 486 399 489 
rect 396 489 399 492 
rect 396 492 399 495 
rect 396 495 399 498 
rect 396 498 399 501 
rect 396 501 399 504 
rect 396 504 399 507 
rect 396 507 399 510 
rect 399 0 402 3 
rect 399 3 402 6 
rect 399 6 402 9 
rect 399 9 402 12 
rect 399 12 402 15 
rect 399 15 402 18 
rect 399 18 402 21 
rect 399 21 402 24 
rect 399 24 402 27 
rect 399 27 402 30 
rect 399 30 402 33 
rect 399 33 402 36 
rect 399 36 402 39 
rect 399 39 402 42 
rect 399 42 402 45 
rect 399 45 402 48 
rect 399 48 402 51 
rect 399 51 402 54 
rect 399 54 402 57 
rect 399 57 402 60 
rect 399 60 402 63 
rect 399 63 402 66 
rect 399 66 402 69 
rect 399 69 402 72 
rect 399 72 402 75 
rect 399 75 402 78 
rect 399 78 402 81 
rect 399 81 402 84 
rect 399 84 402 87 
rect 399 87 402 90 
rect 399 90 402 93 
rect 399 93 402 96 
rect 399 96 402 99 
rect 399 99 402 102 
rect 399 102 402 105 
rect 399 105 402 108 
rect 399 108 402 111 
rect 399 111 402 114 
rect 399 114 402 117 
rect 399 117 402 120 
rect 399 120 402 123 
rect 399 123 402 126 
rect 399 126 402 129 
rect 399 129 402 132 
rect 399 132 402 135 
rect 399 135 402 138 
rect 399 138 402 141 
rect 399 141 402 144 
rect 399 144 402 147 
rect 399 147 402 150 
rect 399 150 402 153 
rect 399 153 402 156 
rect 399 156 402 159 
rect 399 159 402 162 
rect 399 162 402 165 
rect 399 165 402 168 
rect 399 168 402 171 
rect 399 171 402 174 
rect 399 174 402 177 
rect 399 177 402 180 
rect 399 180 402 183 
rect 399 183 402 186 
rect 399 186 402 189 
rect 399 189 402 192 
rect 399 192 402 195 
rect 399 195 402 198 
rect 399 198 402 201 
rect 399 201 402 204 
rect 399 204 402 207 
rect 399 207 402 210 
rect 399 210 402 213 
rect 399 213 402 216 
rect 399 216 402 219 
rect 399 219 402 222 
rect 399 222 402 225 
rect 399 225 402 228 
rect 399 228 402 231 
rect 399 231 402 234 
rect 399 234 402 237 
rect 399 237 402 240 
rect 399 240 402 243 
rect 399 243 402 246 
rect 399 246 402 249 
rect 399 249 402 252 
rect 399 252 402 255 
rect 399 255 402 258 
rect 399 258 402 261 
rect 399 261 402 264 
rect 399 264 402 267 
rect 399 267 402 270 
rect 399 270 402 273 
rect 399 273 402 276 
rect 399 276 402 279 
rect 399 279 402 282 
rect 399 282 402 285 
rect 399 285 402 288 
rect 399 288 402 291 
rect 399 291 402 294 
rect 399 294 402 297 
rect 399 297 402 300 
rect 399 300 402 303 
rect 399 303 402 306 
rect 399 306 402 309 
rect 399 309 402 312 
rect 399 312 402 315 
rect 399 315 402 318 
rect 399 318 402 321 
rect 399 321 402 324 
rect 399 324 402 327 
rect 399 327 402 330 
rect 399 330 402 333 
rect 399 333 402 336 
rect 399 336 402 339 
rect 399 339 402 342 
rect 399 342 402 345 
rect 399 345 402 348 
rect 399 348 402 351 
rect 399 351 402 354 
rect 399 354 402 357 
rect 399 357 402 360 
rect 399 360 402 363 
rect 399 363 402 366 
rect 399 366 402 369 
rect 399 369 402 372 
rect 399 372 402 375 
rect 399 375 402 378 
rect 399 378 402 381 
rect 399 381 402 384 
rect 399 384 402 387 
rect 399 387 402 390 
rect 399 390 402 393 
rect 399 393 402 396 
rect 399 396 402 399 
rect 399 399 402 402 
rect 399 402 402 405 
rect 399 405 402 408 
rect 399 408 402 411 
rect 399 411 402 414 
rect 399 414 402 417 
rect 399 417 402 420 
rect 399 420 402 423 
rect 399 423 402 426 
rect 399 426 402 429 
rect 399 429 402 432 
rect 399 432 402 435 
rect 399 435 402 438 
rect 399 438 402 441 
rect 399 441 402 444 
rect 399 444 402 447 
rect 399 447 402 450 
rect 399 450 402 453 
rect 399 453 402 456 
rect 399 456 402 459 
rect 399 459 402 462 
rect 399 462 402 465 
rect 399 465 402 468 
rect 399 468 402 471 
rect 399 471 402 474 
rect 399 474 402 477 
rect 399 477 402 480 
rect 399 480 402 483 
rect 399 483 402 486 
rect 399 486 402 489 
rect 399 489 402 492 
rect 399 492 402 495 
rect 399 495 402 498 
rect 399 498 402 501 
rect 399 501 402 504 
rect 399 504 402 507 
rect 399 507 402 510 
rect 402 0 405 3 
rect 402 3 405 6 
rect 402 6 405 9 
rect 402 9 405 12 
rect 402 12 405 15 
rect 402 15 405 18 
rect 402 18 405 21 
rect 402 21 405 24 
rect 402 24 405 27 
rect 402 27 405 30 
rect 402 30 405 33 
rect 402 33 405 36 
rect 402 36 405 39 
rect 402 39 405 42 
rect 402 42 405 45 
rect 402 45 405 48 
rect 402 48 405 51 
rect 402 51 405 54 
rect 402 54 405 57 
rect 402 57 405 60 
rect 402 60 405 63 
rect 402 63 405 66 
rect 402 66 405 69 
rect 402 69 405 72 
rect 402 72 405 75 
rect 402 75 405 78 
rect 402 78 405 81 
rect 402 81 405 84 
rect 402 84 405 87 
rect 402 87 405 90 
rect 402 90 405 93 
rect 402 93 405 96 
rect 402 96 405 99 
rect 402 99 405 102 
rect 402 102 405 105 
rect 402 105 405 108 
rect 402 108 405 111 
rect 402 111 405 114 
rect 402 114 405 117 
rect 402 117 405 120 
rect 402 120 405 123 
rect 402 123 405 126 
rect 402 126 405 129 
rect 402 129 405 132 
rect 402 132 405 135 
rect 402 135 405 138 
rect 402 138 405 141 
rect 402 141 405 144 
rect 402 144 405 147 
rect 402 147 405 150 
rect 402 150 405 153 
rect 402 153 405 156 
rect 402 156 405 159 
rect 402 159 405 162 
rect 402 162 405 165 
rect 402 165 405 168 
rect 402 168 405 171 
rect 402 171 405 174 
rect 402 174 405 177 
rect 402 177 405 180 
rect 402 180 405 183 
rect 402 183 405 186 
rect 402 186 405 189 
rect 402 189 405 192 
rect 402 192 405 195 
rect 402 195 405 198 
rect 402 198 405 201 
rect 402 201 405 204 
rect 402 204 405 207 
rect 402 207 405 210 
rect 402 210 405 213 
rect 402 213 405 216 
rect 402 216 405 219 
rect 402 219 405 222 
rect 402 222 405 225 
rect 402 225 405 228 
rect 402 228 405 231 
rect 402 231 405 234 
rect 402 234 405 237 
rect 402 237 405 240 
rect 402 240 405 243 
rect 402 243 405 246 
rect 402 246 405 249 
rect 402 249 405 252 
rect 402 252 405 255 
rect 402 255 405 258 
rect 402 258 405 261 
rect 402 261 405 264 
rect 402 264 405 267 
rect 402 267 405 270 
rect 402 270 405 273 
rect 402 273 405 276 
rect 402 276 405 279 
rect 402 279 405 282 
rect 402 282 405 285 
rect 402 285 405 288 
rect 402 288 405 291 
rect 402 291 405 294 
rect 402 294 405 297 
rect 402 297 405 300 
rect 402 300 405 303 
rect 402 303 405 306 
rect 402 306 405 309 
rect 402 309 405 312 
rect 402 312 405 315 
rect 402 315 405 318 
rect 402 318 405 321 
rect 402 321 405 324 
rect 402 324 405 327 
rect 402 327 405 330 
rect 402 330 405 333 
rect 402 333 405 336 
rect 402 336 405 339 
rect 402 339 405 342 
rect 402 342 405 345 
rect 402 345 405 348 
rect 402 348 405 351 
rect 402 351 405 354 
rect 402 354 405 357 
rect 402 357 405 360 
rect 402 360 405 363 
rect 402 363 405 366 
rect 402 366 405 369 
rect 402 369 405 372 
rect 402 372 405 375 
rect 402 375 405 378 
rect 402 378 405 381 
rect 402 381 405 384 
rect 402 384 405 387 
rect 402 387 405 390 
rect 402 390 405 393 
rect 402 393 405 396 
rect 402 396 405 399 
rect 402 399 405 402 
rect 402 402 405 405 
rect 402 405 405 408 
rect 402 408 405 411 
rect 402 411 405 414 
rect 402 414 405 417 
rect 402 417 405 420 
rect 402 420 405 423 
rect 402 423 405 426 
rect 402 426 405 429 
rect 402 429 405 432 
rect 402 432 405 435 
rect 402 435 405 438 
rect 402 438 405 441 
rect 402 441 405 444 
rect 402 444 405 447 
rect 402 447 405 450 
rect 402 450 405 453 
rect 402 453 405 456 
rect 402 456 405 459 
rect 402 459 405 462 
rect 402 462 405 465 
rect 402 465 405 468 
rect 402 468 405 471 
rect 402 471 405 474 
rect 402 474 405 477 
rect 402 477 405 480 
rect 402 480 405 483 
rect 402 483 405 486 
rect 402 486 405 489 
rect 402 489 405 492 
rect 402 492 405 495 
rect 402 495 405 498 
rect 402 498 405 501 
rect 402 501 405 504 
rect 402 504 405 507 
rect 402 507 405 510 
rect 405 0 408 3 
rect 405 3 408 6 
rect 405 6 408 9 
rect 405 9 408 12 
rect 405 12 408 15 
rect 405 15 408 18 
rect 405 18 408 21 
rect 405 21 408 24 
rect 405 24 408 27 
rect 405 27 408 30 
rect 405 30 408 33 
rect 405 33 408 36 
rect 405 36 408 39 
rect 405 39 408 42 
rect 405 42 408 45 
rect 405 45 408 48 
rect 405 48 408 51 
rect 405 51 408 54 
rect 405 54 408 57 
rect 405 57 408 60 
rect 405 60 408 63 
rect 405 63 408 66 
rect 405 66 408 69 
rect 405 69 408 72 
rect 405 72 408 75 
rect 405 75 408 78 
rect 405 78 408 81 
rect 405 81 408 84 
rect 405 84 408 87 
rect 405 87 408 90 
rect 405 90 408 93 
rect 405 93 408 96 
rect 405 96 408 99 
rect 405 99 408 102 
rect 405 102 408 105 
rect 405 105 408 108 
rect 405 108 408 111 
rect 405 111 408 114 
rect 405 114 408 117 
rect 405 117 408 120 
rect 405 120 408 123 
rect 405 123 408 126 
rect 405 126 408 129 
rect 405 129 408 132 
rect 405 132 408 135 
rect 405 135 408 138 
rect 405 138 408 141 
rect 405 141 408 144 
rect 405 144 408 147 
rect 405 147 408 150 
rect 405 150 408 153 
rect 405 153 408 156 
rect 405 156 408 159 
rect 405 159 408 162 
rect 405 162 408 165 
rect 405 165 408 168 
rect 405 168 408 171 
rect 405 171 408 174 
rect 405 174 408 177 
rect 405 177 408 180 
rect 405 180 408 183 
rect 405 183 408 186 
rect 405 186 408 189 
rect 405 189 408 192 
rect 405 192 408 195 
rect 405 195 408 198 
rect 405 198 408 201 
rect 405 201 408 204 
rect 405 204 408 207 
rect 405 207 408 210 
rect 405 210 408 213 
rect 405 213 408 216 
rect 405 216 408 219 
rect 405 219 408 222 
rect 405 222 408 225 
rect 405 225 408 228 
rect 405 228 408 231 
rect 405 231 408 234 
rect 405 234 408 237 
rect 405 237 408 240 
rect 405 240 408 243 
rect 405 243 408 246 
rect 405 246 408 249 
rect 405 249 408 252 
rect 405 252 408 255 
rect 405 255 408 258 
rect 405 258 408 261 
rect 405 261 408 264 
rect 405 264 408 267 
rect 405 267 408 270 
rect 405 270 408 273 
rect 405 273 408 276 
rect 405 276 408 279 
rect 405 279 408 282 
rect 405 282 408 285 
rect 405 285 408 288 
rect 405 288 408 291 
rect 405 291 408 294 
rect 405 294 408 297 
rect 405 297 408 300 
rect 405 300 408 303 
rect 405 303 408 306 
rect 405 306 408 309 
rect 405 309 408 312 
rect 405 312 408 315 
rect 405 315 408 318 
rect 405 318 408 321 
rect 405 321 408 324 
rect 405 324 408 327 
rect 405 327 408 330 
rect 405 330 408 333 
rect 405 333 408 336 
rect 405 336 408 339 
rect 405 339 408 342 
rect 405 342 408 345 
rect 405 345 408 348 
rect 405 348 408 351 
rect 405 351 408 354 
rect 405 354 408 357 
rect 405 357 408 360 
rect 405 360 408 363 
rect 405 363 408 366 
rect 405 366 408 369 
rect 405 369 408 372 
rect 405 372 408 375 
rect 405 375 408 378 
rect 405 378 408 381 
rect 405 381 408 384 
rect 405 384 408 387 
rect 405 387 408 390 
rect 405 390 408 393 
rect 405 393 408 396 
rect 405 396 408 399 
rect 405 399 408 402 
rect 405 402 408 405 
rect 405 405 408 408 
rect 405 408 408 411 
rect 405 411 408 414 
rect 405 414 408 417 
rect 405 417 408 420 
rect 405 420 408 423 
rect 405 423 408 426 
rect 405 426 408 429 
rect 405 429 408 432 
rect 405 432 408 435 
rect 405 435 408 438 
rect 405 438 408 441 
rect 405 441 408 444 
rect 405 444 408 447 
rect 405 447 408 450 
rect 405 450 408 453 
rect 405 453 408 456 
rect 405 456 408 459 
rect 405 459 408 462 
rect 405 462 408 465 
rect 405 465 408 468 
rect 405 468 408 471 
rect 405 471 408 474 
rect 405 474 408 477 
rect 405 477 408 480 
rect 405 480 408 483 
rect 405 483 408 486 
rect 405 486 408 489 
rect 405 489 408 492 
rect 405 492 408 495 
rect 405 495 408 498 
rect 405 498 408 501 
rect 405 501 408 504 
rect 405 504 408 507 
rect 405 507 408 510 
rect 408 0 411 3 
rect 408 3 411 6 
rect 408 6 411 9 
rect 408 9 411 12 
rect 408 12 411 15 
rect 408 15 411 18 
rect 408 18 411 21 
rect 408 21 411 24 
rect 408 24 411 27 
rect 408 27 411 30 
rect 408 30 411 33 
rect 408 33 411 36 
rect 408 36 411 39 
rect 408 39 411 42 
rect 408 42 411 45 
rect 408 45 411 48 
rect 408 48 411 51 
rect 408 51 411 54 
rect 408 54 411 57 
rect 408 57 411 60 
rect 408 60 411 63 
rect 408 63 411 66 
rect 408 66 411 69 
rect 408 69 411 72 
rect 408 72 411 75 
rect 408 75 411 78 
rect 408 78 411 81 
rect 408 81 411 84 
rect 408 84 411 87 
rect 408 87 411 90 
rect 408 90 411 93 
rect 408 93 411 96 
rect 408 96 411 99 
rect 408 99 411 102 
rect 408 102 411 105 
rect 408 105 411 108 
rect 408 108 411 111 
rect 408 111 411 114 
rect 408 114 411 117 
rect 408 117 411 120 
rect 408 120 411 123 
rect 408 123 411 126 
rect 408 126 411 129 
rect 408 129 411 132 
rect 408 132 411 135 
rect 408 135 411 138 
rect 408 138 411 141 
rect 408 141 411 144 
rect 408 144 411 147 
rect 408 147 411 150 
rect 408 150 411 153 
rect 408 153 411 156 
rect 408 156 411 159 
rect 408 159 411 162 
rect 408 162 411 165 
rect 408 165 411 168 
rect 408 168 411 171 
rect 408 171 411 174 
rect 408 174 411 177 
rect 408 177 411 180 
rect 408 180 411 183 
rect 408 183 411 186 
rect 408 186 411 189 
rect 408 189 411 192 
rect 408 192 411 195 
rect 408 195 411 198 
rect 408 198 411 201 
rect 408 201 411 204 
rect 408 204 411 207 
rect 408 207 411 210 
rect 408 210 411 213 
rect 408 213 411 216 
rect 408 216 411 219 
rect 408 219 411 222 
rect 408 222 411 225 
rect 408 225 411 228 
rect 408 228 411 231 
rect 408 231 411 234 
rect 408 234 411 237 
rect 408 237 411 240 
rect 408 240 411 243 
rect 408 243 411 246 
rect 408 246 411 249 
rect 408 249 411 252 
rect 408 252 411 255 
rect 408 255 411 258 
rect 408 258 411 261 
rect 408 261 411 264 
rect 408 264 411 267 
rect 408 267 411 270 
rect 408 270 411 273 
rect 408 273 411 276 
rect 408 276 411 279 
rect 408 279 411 282 
rect 408 282 411 285 
rect 408 285 411 288 
rect 408 288 411 291 
rect 408 291 411 294 
rect 408 294 411 297 
rect 408 297 411 300 
rect 408 300 411 303 
rect 408 303 411 306 
rect 408 306 411 309 
rect 408 309 411 312 
rect 408 312 411 315 
rect 408 315 411 318 
rect 408 318 411 321 
rect 408 321 411 324 
rect 408 324 411 327 
rect 408 327 411 330 
rect 408 330 411 333 
rect 408 333 411 336 
rect 408 336 411 339 
rect 408 339 411 342 
rect 408 342 411 345 
rect 408 345 411 348 
rect 408 348 411 351 
rect 408 351 411 354 
rect 408 354 411 357 
rect 408 357 411 360 
rect 408 360 411 363 
rect 408 363 411 366 
rect 408 366 411 369 
rect 408 369 411 372 
rect 408 372 411 375 
rect 408 375 411 378 
rect 408 378 411 381 
rect 408 381 411 384 
rect 408 384 411 387 
rect 408 387 411 390 
rect 408 390 411 393 
rect 408 393 411 396 
rect 408 396 411 399 
rect 408 399 411 402 
rect 408 402 411 405 
rect 408 405 411 408 
rect 408 408 411 411 
rect 408 411 411 414 
rect 408 414 411 417 
rect 408 417 411 420 
rect 408 420 411 423 
rect 408 423 411 426 
rect 408 426 411 429 
rect 408 429 411 432 
rect 408 432 411 435 
rect 408 435 411 438 
rect 408 438 411 441 
rect 408 441 411 444 
rect 408 444 411 447 
rect 408 447 411 450 
rect 408 450 411 453 
rect 408 453 411 456 
rect 408 456 411 459 
rect 408 459 411 462 
rect 408 462 411 465 
rect 408 465 411 468 
rect 408 468 411 471 
rect 408 471 411 474 
rect 408 474 411 477 
rect 408 477 411 480 
rect 408 480 411 483 
rect 408 483 411 486 
rect 408 486 411 489 
rect 408 489 411 492 
rect 408 492 411 495 
rect 408 495 411 498 
rect 408 498 411 501 
rect 408 501 411 504 
rect 408 504 411 507 
rect 408 507 411 510 
rect 411 0 414 3 
rect 411 3 414 6 
rect 411 6 414 9 
rect 411 9 414 12 
rect 411 12 414 15 
rect 411 15 414 18 
rect 411 18 414 21 
rect 411 21 414 24 
rect 411 24 414 27 
rect 411 27 414 30 
rect 411 30 414 33 
rect 411 33 414 36 
rect 411 36 414 39 
rect 411 39 414 42 
rect 411 42 414 45 
rect 411 45 414 48 
rect 411 48 414 51 
rect 411 51 414 54 
rect 411 54 414 57 
rect 411 57 414 60 
rect 411 60 414 63 
rect 411 63 414 66 
rect 411 66 414 69 
rect 411 69 414 72 
rect 411 72 414 75 
rect 411 75 414 78 
rect 411 78 414 81 
rect 411 81 414 84 
rect 411 84 414 87 
rect 411 87 414 90 
rect 411 90 414 93 
rect 411 93 414 96 
rect 411 96 414 99 
rect 411 99 414 102 
rect 411 102 414 105 
rect 411 105 414 108 
rect 411 108 414 111 
rect 411 111 414 114 
rect 411 114 414 117 
rect 411 117 414 120 
rect 411 120 414 123 
rect 411 123 414 126 
rect 411 126 414 129 
rect 411 129 414 132 
rect 411 132 414 135 
rect 411 135 414 138 
rect 411 138 414 141 
rect 411 141 414 144 
rect 411 144 414 147 
rect 411 147 414 150 
rect 411 150 414 153 
rect 411 153 414 156 
rect 411 156 414 159 
rect 411 159 414 162 
rect 411 162 414 165 
rect 411 165 414 168 
rect 411 168 414 171 
rect 411 171 414 174 
rect 411 174 414 177 
rect 411 177 414 180 
rect 411 180 414 183 
rect 411 183 414 186 
rect 411 186 414 189 
rect 411 189 414 192 
rect 411 192 414 195 
rect 411 195 414 198 
rect 411 198 414 201 
rect 411 201 414 204 
rect 411 204 414 207 
rect 411 207 414 210 
rect 411 210 414 213 
rect 411 213 414 216 
rect 411 216 414 219 
rect 411 219 414 222 
rect 411 222 414 225 
rect 411 225 414 228 
rect 411 228 414 231 
rect 411 231 414 234 
rect 411 234 414 237 
rect 411 237 414 240 
rect 411 240 414 243 
rect 411 243 414 246 
rect 411 246 414 249 
rect 411 249 414 252 
rect 411 252 414 255 
rect 411 255 414 258 
rect 411 258 414 261 
rect 411 261 414 264 
rect 411 264 414 267 
rect 411 267 414 270 
rect 411 270 414 273 
rect 411 273 414 276 
rect 411 276 414 279 
rect 411 279 414 282 
rect 411 282 414 285 
rect 411 285 414 288 
rect 411 288 414 291 
rect 411 291 414 294 
rect 411 294 414 297 
rect 411 297 414 300 
rect 411 300 414 303 
rect 411 303 414 306 
rect 411 306 414 309 
rect 411 309 414 312 
rect 411 312 414 315 
rect 411 315 414 318 
rect 411 318 414 321 
rect 411 321 414 324 
rect 411 324 414 327 
rect 411 327 414 330 
rect 411 330 414 333 
rect 411 333 414 336 
rect 411 336 414 339 
rect 411 339 414 342 
rect 411 342 414 345 
rect 411 345 414 348 
rect 411 348 414 351 
rect 411 351 414 354 
rect 411 354 414 357 
rect 411 357 414 360 
rect 411 360 414 363 
rect 411 363 414 366 
rect 411 366 414 369 
rect 411 369 414 372 
rect 411 372 414 375 
rect 411 375 414 378 
rect 411 378 414 381 
rect 411 381 414 384 
rect 411 384 414 387 
rect 411 387 414 390 
rect 411 390 414 393 
rect 411 393 414 396 
rect 411 396 414 399 
rect 411 399 414 402 
rect 411 402 414 405 
rect 411 405 414 408 
rect 411 408 414 411 
rect 411 411 414 414 
rect 411 414 414 417 
rect 411 417 414 420 
rect 411 420 414 423 
rect 411 423 414 426 
rect 411 426 414 429 
rect 411 429 414 432 
rect 411 432 414 435 
rect 411 435 414 438 
rect 411 438 414 441 
rect 411 441 414 444 
rect 411 444 414 447 
rect 411 447 414 450 
rect 411 450 414 453 
rect 411 453 414 456 
rect 411 456 414 459 
rect 411 459 414 462 
rect 411 462 414 465 
rect 411 465 414 468 
rect 411 468 414 471 
rect 411 471 414 474 
rect 411 474 414 477 
rect 411 477 414 480 
rect 411 480 414 483 
rect 411 483 414 486 
rect 411 486 414 489 
rect 411 489 414 492 
rect 411 492 414 495 
rect 411 495 414 498 
rect 411 498 414 501 
rect 411 501 414 504 
rect 411 504 414 507 
rect 411 507 414 510 
rect 414 0 417 3 
rect 414 3 417 6 
rect 414 6 417 9 
rect 414 9 417 12 
rect 414 12 417 15 
rect 414 15 417 18 
rect 414 18 417 21 
rect 414 21 417 24 
rect 414 24 417 27 
rect 414 27 417 30 
rect 414 30 417 33 
rect 414 33 417 36 
rect 414 36 417 39 
rect 414 39 417 42 
rect 414 42 417 45 
rect 414 45 417 48 
rect 414 48 417 51 
rect 414 51 417 54 
rect 414 54 417 57 
rect 414 57 417 60 
rect 414 60 417 63 
rect 414 63 417 66 
rect 414 66 417 69 
rect 414 69 417 72 
rect 414 72 417 75 
rect 414 75 417 78 
rect 414 78 417 81 
rect 414 81 417 84 
rect 414 84 417 87 
rect 414 87 417 90 
rect 414 90 417 93 
rect 414 93 417 96 
rect 414 96 417 99 
rect 414 99 417 102 
rect 414 102 417 105 
rect 414 105 417 108 
rect 414 108 417 111 
rect 414 111 417 114 
rect 414 114 417 117 
rect 414 117 417 120 
rect 414 120 417 123 
rect 414 123 417 126 
rect 414 126 417 129 
rect 414 129 417 132 
rect 414 132 417 135 
rect 414 135 417 138 
rect 414 138 417 141 
rect 414 141 417 144 
rect 414 144 417 147 
rect 414 147 417 150 
rect 414 150 417 153 
rect 414 153 417 156 
rect 414 156 417 159 
rect 414 159 417 162 
rect 414 162 417 165 
rect 414 165 417 168 
rect 414 168 417 171 
rect 414 171 417 174 
rect 414 174 417 177 
rect 414 177 417 180 
rect 414 180 417 183 
rect 414 183 417 186 
rect 414 186 417 189 
rect 414 189 417 192 
rect 414 192 417 195 
rect 414 195 417 198 
rect 414 198 417 201 
rect 414 201 417 204 
rect 414 204 417 207 
rect 414 207 417 210 
rect 414 210 417 213 
rect 414 213 417 216 
rect 414 216 417 219 
rect 414 219 417 222 
rect 414 222 417 225 
rect 414 225 417 228 
rect 414 228 417 231 
rect 414 231 417 234 
rect 414 234 417 237 
rect 414 237 417 240 
rect 414 240 417 243 
rect 414 243 417 246 
rect 414 246 417 249 
rect 414 249 417 252 
rect 414 252 417 255 
rect 414 255 417 258 
rect 414 258 417 261 
rect 414 261 417 264 
rect 414 264 417 267 
rect 414 267 417 270 
rect 414 270 417 273 
rect 414 273 417 276 
rect 414 276 417 279 
rect 414 279 417 282 
rect 414 282 417 285 
rect 414 285 417 288 
rect 414 288 417 291 
rect 414 291 417 294 
rect 414 294 417 297 
rect 414 297 417 300 
rect 414 300 417 303 
rect 414 303 417 306 
rect 414 306 417 309 
rect 414 309 417 312 
rect 414 312 417 315 
rect 414 315 417 318 
rect 414 318 417 321 
rect 414 321 417 324 
rect 414 324 417 327 
rect 414 327 417 330 
rect 414 330 417 333 
rect 414 333 417 336 
rect 414 336 417 339 
rect 414 339 417 342 
rect 414 342 417 345 
rect 414 345 417 348 
rect 414 348 417 351 
rect 414 351 417 354 
rect 414 354 417 357 
rect 414 357 417 360 
rect 414 360 417 363 
rect 414 363 417 366 
rect 414 366 417 369 
rect 414 369 417 372 
rect 414 372 417 375 
rect 414 375 417 378 
rect 414 378 417 381 
rect 414 381 417 384 
rect 414 384 417 387 
rect 414 387 417 390 
rect 414 390 417 393 
rect 414 393 417 396 
rect 414 396 417 399 
rect 414 399 417 402 
rect 414 402 417 405 
rect 414 405 417 408 
rect 414 408 417 411 
rect 414 411 417 414 
rect 414 414 417 417 
rect 414 417 417 420 
rect 414 420 417 423 
rect 414 423 417 426 
rect 414 426 417 429 
rect 414 429 417 432 
rect 414 432 417 435 
rect 414 435 417 438 
rect 414 438 417 441 
rect 414 441 417 444 
rect 414 444 417 447 
rect 414 447 417 450 
rect 414 450 417 453 
rect 414 453 417 456 
rect 414 456 417 459 
rect 414 459 417 462 
rect 414 462 417 465 
rect 414 465 417 468 
rect 414 468 417 471 
rect 414 471 417 474 
rect 414 474 417 477 
rect 414 477 417 480 
rect 414 480 417 483 
rect 414 483 417 486 
rect 414 486 417 489 
rect 414 489 417 492 
rect 414 492 417 495 
rect 414 495 417 498 
rect 414 498 417 501 
rect 414 501 417 504 
rect 414 504 417 507 
rect 414 507 417 510 
rect 417 0 420 3 
rect 417 3 420 6 
rect 417 6 420 9 
rect 417 9 420 12 
rect 417 12 420 15 
rect 417 15 420 18 
rect 417 18 420 21 
rect 417 21 420 24 
rect 417 24 420 27 
rect 417 27 420 30 
rect 417 30 420 33 
rect 417 33 420 36 
rect 417 36 420 39 
rect 417 39 420 42 
rect 417 42 420 45 
rect 417 45 420 48 
rect 417 48 420 51 
rect 417 51 420 54 
rect 417 54 420 57 
rect 417 57 420 60 
rect 417 60 420 63 
rect 417 63 420 66 
rect 417 66 420 69 
rect 417 69 420 72 
rect 417 72 420 75 
rect 417 75 420 78 
rect 417 78 420 81 
rect 417 81 420 84 
rect 417 84 420 87 
rect 417 87 420 90 
rect 417 90 420 93 
rect 417 93 420 96 
rect 417 96 420 99 
rect 417 99 420 102 
rect 417 102 420 105 
rect 417 105 420 108 
rect 417 108 420 111 
rect 417 111 420 114 
rect 417 114 420 117 
rect 417 117 420 120 
rect 417 120 420 123 
rect 417 123 420 126 
rect 417 126 420 129 
rect 417 129 420 132 
rect 417 132 420 135 
rect 417 135 420 138 
rect 417 138 420 141 
rect 417 141 420 144 
rect 417 144 420 147 
rect 417 147 420 150 
rect 417 150 420 153 
rect 417 153 420 156 
rect 417 156 420 159 
rect 417 159 420 162 
rect 417 162 420 165 
rect 417 165 420 168 
rect 417 168 420 171 
rect 417 171 420 174 
rect 417 174 420 177 
rect 417 177 420 180 
rect 417 180 420 183 
rect 417 183 420 186 
rect 417 186 420 189 
rect 417 189 420 192 
rect 417 192 420 195 
rect 417 195 420 198 
rect 417 198 420 201 
rect 417 201 420 204 
rect 417 204 420 207 
rect 417 207 420 210 
rect 417 210 420 213 
rect 417 213 420 216 
rect 417 216 420 219 
rect 417 219 420 222 
rect 417 222 420 225 
rect 417 225 420 228 
rect 417 228 420 231 
rect 417 231 420 234 
rect 417 234 420 237 
rect 417 237 420 240 
rect 417 240 420 243 
rect 417 243 420 246 
rect 417 246 420 249 
rect 417 249 420 252 
rect 417 252 420 255 
rect 417 255 420 258 
rect 417 258 420 261 
rect 417 261 420 264 
rect 417 264 420 267 
rect 417 267 420 270 
rect 417 270 420 273 
rect 417 273 420 276 
rect 417 276 420 279 
rect 417 279 420 282 
rect 417 282 420 285 
rect 417 285 420 288 
rect 417 288 420 291 
rect 417 291 420 294 
rect 417 294 420 297 
rect 417 297 420 300 
rect 417 300 420 303 
rect 417 303 420 306 
rect 417 306 420 309 
rect 417 309 420 312 
rect 417 312 420 315 
rect 417 315 420 318 
rect 417 318 420 321 
rect 417 321 420 324 
rect 417 324 420 327 
rect 417 327 420 330 
rect 417 330 420 333 
rect 417 333 420 336 
rect 417 336 420 339 
rect 417 339 420 342 
rect 417 342 420 345 
rect 417 345 420 348 
rect 417 348 420 351 
rect 417 351 420 354 
rect 417 354 420 357 
rect 417 357 420 360 
rect 417 360 420 363 
rect 417 363 420 366 
rect 417 366 420 369 
rect 417 369 420 372 
rect 417 372 420 375 
rect 417 375 420 378 
rect 417 378 420 381 
rect 417 381 420 384 
rect 417 384 420 387 
rect 417 387 420 390 
rect 417 390 420 393 
rect 417 393 420 396 
rect 417 396 420 399 
rect 417 399 420 402 
rect 417 402 420 405 
rect 417 405 420 408 
rect 417 408 420 411 
rect 417 411 420 414 
rect 417 414 420 417 
rect 417 417 420 420 
rect 417 420 420 423 
rect 417 423 420 426 
rect 417 426 420 429 
rect 417 429 420 432 
rect 417 432 420 435 
rect 417 435 420 438 
rect 417 438 420 441 
rect 417 441 420 444 
rect 417 444 420 447 
rect 417 447 420 450 
rect 417 450 420 453 
rect 417 453 420 456 
rect 417 456 420 459 
rect 417 459 420 462 
rect 417 462 420 465 
rect 417 465 420 468 
rect 417 468 420 471 
rect 417 471 420 474 
rect 417 474 420 477 
rect 417 477 420 480 
rect 417 480 420 483 
rect 417 483 420 486 
rect 417 486 420 489 
rect 417 489 420 492 
rect 417 492 420 495 
rect 417 495 420 498 
rect 417 498 420 501 
rect 417 501 420 504 
rect 417 504 420 507 
rect 417 507 420 510 
rect 420 0 423 3 
rect 420 3 423 6 
rect 420 6 423 9 
rect 420 9 423 12 
rect 420 12 423 15 
rect 420 15 423 18 
rect 420 18 423 21 
rect 420 21 423 24 
rect 420 24 423 27 
rect 420 27 423 30 
rect 420 30 423 33 
rect 420 33 423 36 
rect 420 36 423 39 
rect 420 39 423 42 
rect 420 42 423 45 
rect 420 45 423 48 
rect 420 48 423 51 
rect 420 51 423 54 
rect 420 54 423 57 
rect 420 57 423 60 
rect 420 60 423 63 
rect 420 63 423 66 
rect 420 66 423 69 
rect 420 69 423 72 
rect 420 72 423 75 
rect 420 75 423 78 
rect 420 78 423 81 
rect 420 81 423 84 
rect 420 84 423 87 
rect 420 87 423 90 
rect 420 90 423 93 
rect 420 93 423 96 
rect 420 96 423 99 
rect 420 99 423 102 
rect 420 102 423 105 
rect 420 105 423 108 
rect 420 108 423 111 
rect 420 111 423 114 
rect 420 114 423 117 
rect 420 117 423 120 
rect 420 120 423 123 
rect 420 123 423 126 
rect 420 126 423 129 
rect 420 129 423 132 
rect 420 132 423 135 
rect 420 135 423 138 
rect 420 138 423 141 
rect 420 141 423 144 
rect 420 144 423 147 
rect 420 147 423 150 
rect 420 150 423 153 
rect 420 153 423 156 
rect 420 156 423 159 
rect 420 159 423 162 
rect 420 162 423 165 
rect 420 165 423 168 
rect 420 168 423 171 
rect 420 171 423 174 
rect 420 174 423 177 
rect 420 177 423 180 
rect 420 180 423 183 
rect 420 183 423 186 
rect 420 186 423 189 
rect 420 189 423 192 
rect 420 192 423 195 
rect 420 195 423 198 
rect 420 198 423 201 
rect 420 201 423 204 
rect 420 204 423 207 
rect 420 207 423 210 
rect 420 210 423 213 
rect 420 213 423 216 
rect 420 216 423 219 
rect 420 219 423 222 
rect 420 222 423 225 
rect 420 225 423 228 
rect 420 228 423 231 
rect 420 231 423 234 
rect 420 234 423 237 
rect 420 237 423 240 
rect 420 240 423 243 
rect 420 243 423 246 
rect 420 246 423 249 
rect 420 249 423 252 
rect 420 252 423 255 
rect 420 255 423 258 
rect 420 258 423 261 
rect 420 261 423 264 
rect 420 264 423 267 
rect 420 267 423 270 
rect 420 270 423 273 
rect 420 273 423 276 
rect 420 276 423 279 
rect 420 279 423 282 
rect 420 282 423 285 
rect 420 285 423 288 
rect 420 288 423 291 
rect 420 291 423 294 
rect 420 294 423 297 
rect 420 297 423 300 
rect 420 300 423 303 
rect 420 303 423 306 
rect 420 306 423 309 
rect 420 309 423 312 
rect 420 312 423 315 
rect 420 315 423 318 
rect 420 318 423 321 
rect 420 321 423 324 
rect 420 324 423 327 
rect 420 327 423 330 
rect 420 330 423 333 
rect 420 333 423 336 
rect 420 336 423 339 
rect 420 339 423 342 
rect 420 342 423 345 
rect 420 345 423 348 
rect 420 348 423 351 
rect 420 351 423 354 
rect 420 354 423 357 
rect 420 357 423 360 
rect 420 360 423 363 
rect 420 363 423 366 
rect 420 366 423 369 
rect 420 369 423 372 
rect 420 372 423 375 
rect 420 375 423 378 
rect 420 378 423 381 
rect 420 381 423 384 
rect 420 384 423 387 
rect 420 387 423 390 
rect 420 390 423 393 
rect 420 393 423 396 
rect 420 396 423 399 
rect 420 399 423 402 
rect 420 402 423 405 
rect 420 405 423 408 
rect 420 408 423 411 
rect 420 411 423 414 
rect 420 414 423 417 
rect 420 417 423 420 
rect 420 420 423 423 
rect 420 423 423 426 
rect 420 426 423 429 
rect 420 429 423 432 
rect 420 432 423 435 
rect 420 435 423 438 
rect 420 438 423 441 
rect 420 441 423 444 
rect 420 444 423 447 
rect 420 447 423 450 
rect 420 450 423 453 
rect 420 453 423 456 
rect 420 456 423 459 
rect 420 459 423 462 
rect 420 462 423 465 
rect 420 465 423 468 
rect 420 468 423 471 
rect 420 471 423 474 
rect 420 474 423 477 
rect 420 477 423 480 
rect 420 480 423 483 
rect 420 483 423 486 
rect 420 486 423 489 
rect 420 489 423 492 
rect 420 492 423 495 
rect 420 495 423 498 
rect 420 498 423 501 
rect 420 501 423 504 
rect 420 504 423 507 
rect 420 507 423 510 
rect 423 0 426 3 
rect 423 3 426 6 
rect 423 6 426 9 
rect 423 9 426 12 
rect 423 12 426 15 
rect 423 15 426 18 
rect 423 18 426 21 
rect 423 21 426 24 
rect 423 24 426 27 
rect 423 27 426 30 
rect 423 30 426 33 
rect 423 33 426 36 
rect 423 36 426 39 
rect 423 39 426 42 
rect 423 42 426 45 
rect 423 45 426 48 
rect 423 48 426 51 
rect 423 51 426 54 
rect 423 54 426 57 
rect 423 57 426 60 
rect 423 60 426 63 
rect 423 63 426 66 
rect 423 66 426 69 
rect 423 69 426 72 
rect 423 72 426 75 
rect 423 75 426 78 
rect 423 78 426 81 
rect 423 81 426 84 
rect 423 84 426 87 
rect 423 87 426 90 
rect 423 90 426 93 
rect 423 93 426 96 
rect 423 96 426 99 
rect 423 99 426 102 
rect 423 102 426 105 
rect 423 105 426 108 
rect 423 108 426 111 
rect 423 111 426 114 
rect 423 114 426 117 
rect 423 117 426 120 
rect 423 120 426 123 
rect 423 123 426 126 
rect 423 126 426 129 
rect 423 129 426 132 
rect 423 132 426 135 
rect 423 135 426 138 
rect 423 138 426 141 
rect 423 141 426 144 
rect 423 144 426 147 
rect 423 147 426 150 
rect 423 150 426 153 
rect 423 153 426 156 
rect 423 156 426 159 
rect 423 159 426 162 
rect 423 162 426 165 
rect 423 165 426 168 
rect 423 168 426 171 
rect 423 171 426 174 
rect 423 174 426 177 
rect 423 177 426 180 
rect 423 180 426 183 
rect 423 183 426 186 
rect 423 186 426 189 
rect 423 189 426 192 
rect 423 192 426 195 
rect 423 195 426 198 
rect 423 198 426 201 
rect 423 201 426 204 
rect 423 204 426 207 
rect 423 207 426 210 
rect 423 210 426 213 
rect 423 213 426 216 
rect 423 216 426 219 
rect 423 219 426 222 
rect 423 222 426 225 
rect 423 225 426 228 
rect 423 228 426 231 
rect 423 231 426 234 
rect 423 234 426 237 
rect 423 237 426 240 
rect 423 240 426 243 
rect 423 243 426 246 
rect 423 246 426 249 
rect 423 249 426 252 
rect 423 252 426 255 
rect 423 255 426 258 
rect 423 258 426 261 
rect 423 261 426 264 
rect 423 264 426 267 
rect 423 267 426 270 
rect 423 270 426 273 
rect 423 273 426 276 
rect 423 276 426 279 
rect 423 279 426 282 
rect 423 282 426 285 
rect 423 285 426 288 
rect 423 288 426 291 
rect 423 291 426 294 
rect 423 294 426 297 
rect 423 297 426 300 
rect 423 300 426 303 
rect 423 303 426 306 
rect 423 306 426 309 
rect 423 309 426 312 
rect 423 312 426 315 
rect 423 315 426 318 
rect 423 318 426 321 
rect 423 321 426 324 
rect 423 324 426 327 
rect 423 327 426 330 
rect 423 330 426 333 
rect 423 333 426 336 
rect 423 336 426 339 
rect 423 339 426 342 
rect 423 342 426 345 
rect 423 345 426 348 
rect 423 348 426 351 
rect 423 351 426 354 
rect 423 354 426 357 
rect 423 357 426 360 
rect 423 360 426 363 
rect 423 363 426 366 
rect 423 366 426 369 
rect 423 369 426 372 
rect 423 372 426 375 
rect 423 375 426 378 
rect 423 378 426 381 
rect 423 381 426 384 
rect 423 384 426 387 
rect 423 387 426 390 
rect 423 390 426 393 
rect 423 393 426 396 
rect 423 396 426 399 
rect 423 399 426 402 
rect 423 402 426 405 
rect 423 405 426 408 
rect 423 408 426 411 
rect 423 411 426 414 
rect 423 414 426 417 
rect 423 417 426 420 
rect 423 420 426 423 
rect 423 423 426 426 
rect 423 426 426 429 
rect 423 429 426 432 
rect 423 432 426 435 
rect 423 435 426 438 
rect 423 438 426 441 
rect 423 441 426 444 
rect 423 444 426 447 
rect 423 447 426 450 
rect 423 450 426 453 
rect 423 453 426 456 
rect 423 456 426 459 
rect 423 459 426 462 
rect 423 462 426 465 
rect 423 465 426 468 
rect 423 468 426 471 
rect 423 471 426 474 
rect 423 474 426 477 
rect 423 477 426 480 
rect 423 480 426 483 
rect 423 483 426 486 
rect 423 486 426 489 
rect 423 489 426 492 
rect 423 492 426 495 
rect 423 495 426 498 
rect 423 498 426 501 
rect 423 501 426 504 
rect 423 504 426 507 
rect 423 507 426 510 
rect 426 0 429 3 
rect 426 3 429 6 
rect 426 6 429 9 
rect 426 9 429 12 
rect 426 12 429 15 
rect 426 15 429 18 
rect 426 18 429 21 
rect 426 21 429 24 
rect 426 24 429 27 
rect 426 27 429 30 
rect 426 30 429 33 
rect 426 33 429 36 
rect 426 36 429 39 
rect 426 39 429 42 
rect 426 42 429 45 
rect 426 45 429 48 
rect 426 48 429 51 
rect 426 51 429 54 
rect 426 54 429 57 
rect 426 57 429 60 
rect 426 60 429 63 
rect 426 63 429 66 
rect 426 66 429 69 
rect 426 69 429 72 
rect 426 72 429 75 
rect 426 75 429 78 
rect 426 78 429 81 
rect 426 81 429 84 
rect 426 84 429 87 
rect 426 87 429 90 
rect 426 90 429 93 
rect 426 93 429 96 
rect 426 96 429 99 
rect 426 99 429 102 
rect 426 102 429 105 
rect 426 105 429 108 
rect 426 108 429 111 
rect 426 111 429 114 
rect 426 114 429 117 
rect 426 117 429 120 
rect 426 120 429 123 
rect 426 123 429 126 
rect 426 126 429 129 
rect 426 129 429 132 
rect 426 132 429 135 
rect 426 135 429 138 
rect 426 138 429 141 
rect 426 141 429 144 
rect 426 144 429 147 
rect 426 147 429 150 
rect 426 150 429 153 
rect 426 153 429 156 
rect 426 156 429 159 
rect 426 159 429 162 
rect 426 162 429 165 
rect 426 165 429 168 
rect 426 168 429 171 
rect 426 171 429 174 
rect 426 174 429 177 
rect 426 177 429 180 
rect 426 180 429 183 
rect 426 183 429 186 
rect 426 186 429 189 
rect 426 189 429 192 
rect 426 192 429 195 
rect 426 195 429 198 
rect 426 198 429 201 
rect 426 201 429 204 
rect 426 204 429 207 
rect 426 207 429 210 
rect 426 210 429 213 
rect 426 213 429 216 
rect 426 216 429 219 
rect 426 219 429 222 
rect 426 222 429 225 
rect 426 225 429 228 
rect 426 228 429 231 
rect 426 231 429 234 
rect 426 234 429 237 
rect 426 237 429 240 
rect 426 240 429 243 
rect 426 243 429 246 
rect 426 246 429 249 
rect 426 249 429 252 
rect 426 252 429 255 
rect 426 255 429 258 
rect 426 258 429 261 
rect 426 261 429 264 
rect 426 264 429 267 
rect 426 267 429 270 
rect 426 270 429 273 
rect 426 273 429 276 
rect 426 276 429 279 
rect 426 279 429 282 
rect 426 282 429 285 
rect 426 285 429 288 
rect 426 288 429 291 
rect 426 291 429 294 
rect 426 294 429 297 
rect 426 297 429 300 
rect 426 300 429 303 
rect 426 303 429 306 
rect 426 306 429 309 
rect 426 309 429 312 
rect 426 312 429 315 
rect 426 315 429 318 
rect 426 318 429 321 
rect 426 321 429 324 
rect 426 324 429 327 
rect 426 327 429 330 
rect 426 330 429 333 
rect 426 333 429 336 
rect 426 336 429 339 
rect 426 339 429 342 
rect 426 342 429 345 
rect 426 345 429 348 
rect 426 348 429 351 
rect 426 351 429 354 
rect 426 354 429 357 
rect 426 357 429 360 
rect 426 360 429 363 
rect 426 363 429 366 
rect 426 366 429 369 
rect 426 369 429 372 
rect 426 372 429 375 
rect 426 375 429 378 
rect 426 378 429 381 
rect 426 381 429 384 
rect 426 384 429 387 
rect 426 387 429 390 
rect 426 390 429 393 
rect 426 393 429 396 
rect 426 396 429 399 
rect 426 399 429 402 
rect 426 402 429 405 
rect 426 405 429 408 
rect 426 408 429 411 
rect 426 411 429 414 
rect 426 414 429 417 
rect 426 417 429 420 
rect 426 420 429 423 
rect 426 423 429 426 
rect 426 426 429 429 
rect 426 429 429 432 
rect 426 432 429 435 
rect 426 435 429 438 
rect 426 438 429 441 
rect 426 441 429 444 
rect 426 444 429 447 
rect 426 447 429 450 
rect 426 450 429 453 
rect 426 453 429 456 
rect 426 456 429 459 
rect 426 459 429 462 
rect 426 462 429 465 
rect 426 465 429 468 
rect 426 468 429 471 
rect 426 471 429 474 
rect 426 474 429 477 
rect 426 477 429 480 
rect 426 480 429 483 
rect 426 483 429 486 
rect 426 486 429 489 
rect 426 489 429 492 
rect 426 492 429 495 
rect 426 495 429 498 
rect 426 498 429 501 
rect 426 501 429 504 
rect 426 504 429 507 
rect 426 507 429 510 
rect 429 0 432 3 
rect 429 3 432 6 
rect 429 6 432 9 
rect 429 9 432 12 
rect 429 12 432 15 
rect 429 15 432 18 
rect 429 18 432 21 
rect 429 21 432 24 
rect 429 24 432 27 
rect 429 27 432 30 
rect 429 30 432 33 
rect 429 33 432 36 
rect 429 36 432 39 
rect 429 39 432 42 
rect 429 42 432 45 
rect 429 45 432 48 
rect 429 48 432 51 
rect 429 51 432 54 
rect 429 54 432 57 
rect 429 57 432 60 
rect 429 60 432 63 
rect 429 63 432 66 
rect 429 66 432 69 
rect 429 69 432 72 
rect 429 72 432 75 
rect 429 75 432 78 
rect 429 78 432 81 
rect 429 81 432 84 
rect 429 84 432 87 
rect 429 87 432 90 
rect 429 90 432 93 
rect 429 93 432 96 
rect 429 96 432 99 
rect 429 99 432 102 
rect 429 102 432 105 
rect 429 105 432 108 
rect 429 108 432 111 
rect 429 111 432 114 
rect 429 114 432 117 
rect 429 117 432 120 
rect 429 120 432 123 
rect 429 123 432 126 
rect 429 126 432 129 
rect 429 129 432 132 
rect 429 132 432 135 
rect 429 135 432 138 
rect 429 138 432 141 
rect 429 141 432 144 
rect 429 144 432 147 
rect 429 147 432 150 
rect 429 150 432 153 
rect 429 153 432 156 
rect 429 156 432 159 
rect 429 159 432 162 
rect 429 162 432 165 
rect 429 165 432 168 
rect 429 168 432 171 
rect 429 171 432 174 
rect 429 174 432 177 
rect 429 177 432 180 
rect 429 180 432 183 
rect 429 183 432 186 
rect 429 186 432 189 
rect 429 189 432 192 
rect 429 192 432 195 
rect 429 195 432 198 
rect 429 198 432 201 
rect 429 201 432 204 
rect 429 204 432 207 
rect 429 207 432 210 
rect 429 210 432 213 
rect 429 213 432 216 
rect 429 216 432 219 
rect 429 219 432 222 
rect 429 222 432 225 
rect 429 225 432 228 
rect 429 228 432 231 
rect 429 231 432 234 
rect 429 234 432 237 
rect 429 237 432 240 
rect 429 240 432 243 
rect 429 243 432 246 
rect 429 246 432 249 
rect 429 249 432 252 
rect 429 252 432 255 
rect 429 255 432 258 
rect 429 258 432 261 
rect 429 261 432 264 
rect 429 264 432 267 
rect 429 267 432 270 
rect 429 270 432 273 
rect 429 273 432 276 
rect 429 276 432 279 
rect 429 279 432 282 
rect 429 282 432 285 
rect 429 285 432 288 
rect 429 288 432 291 
rect 429 291 432 294 
rect 429 294 432 297 
rect 429 297 432 300 
rect 429 300 432 303 
rect 429 303 432 306 
rect 429 306 432 309 
rect 429 309 432 312 
rect 429 312 432 315 
rect 429 315 432 318 
rect 429 318 432 321 
rect 429 321 432 324 
rect 429 324 432 327 
rect 429 327 432 330 
rect 429 330 432 333 
rect 429 333 432 336 
rect 429 336 432 339 
rect 429 339 432 342 
rect 429 342 432 345 
rect 429 345 432 348 
rect 429 348 432 351 
rect 429 351 432 354 
rect 429 354 432 357 
rect 429 357 432 360 
rect 429 360 432 363 
rect 429 363 432 366 
rect 429 366 432 369 
rect 429 369 432 372 
rect 429 372 432 375 
rect 429 375 432 378 
rect 429 378 432 381 
rect 429 381 432 384 
rect 429 384 432 387 
rect 429 387 432 390 
rect 429 390 432 393 
rect 429 393 432 396 
rect 429 396 432 399 
rect 429 399 432 402 
rect 429 402 432 405 
rect 429 405 432 408 
rect 429 408 432 411 
rect 429 411 432 414 
rect 429 414 432 417 
rect 429 417 432 420 
rect 429 420 432 423 
rect 429 423 432 426 
rect 429 426 432 429 
rect 429 429 432 432 
rect 429 432 432 435 
rect 429 435 432 438 
rect 429 438 432 441 
rect 429 441 432 444 
rect 429 444 432 447 
rect 429 447 432 450 
rect 429 450 432 453 
rect 429 453 432 456 
rect 429 456 432 459 
rect 429 459 432 462 
rect 429 462 432 465 
rect 429 465 432 468 
rect 429 468 432 471 
rect 429 471 432 474 
rect 429 474 432 477 
rect 429 477 432 480 
rect 429 480 432 483 
rect 429 483 432 486 
rect 429 486 432 489 
rect 429 489 432 492 
rect 429 492 432 495 
rect 429 495 432 498 
rect 429 498 432 501 
rect 429 501 432 504 
rect 429 504 432 507 
rect 429 507 432 510 
rect 432 0 435 3 
rect 432 3 435 6 
rect 432 6 435 9 
rect 432 9 435 12 
rect 432 12 435 15 
rect 432 15 435 18 
rect 432 18 435 21 
rect 432 21 435 24 
rect 432 24 435 27 
rect 432 27 435 30 
rect 432 30 435 33 
rect 432 33 435 36 
rect 432 36 435 39 
rect 432 39 435 42 
rect 432 42 435 45 
rect 432 45 435 48 
rect 432 48 435 51 
rect 432 51 435 54 
rect 432 54 435 57 
rect 432 57 435 60 
rect 432 60 435 63 
rect 432 63 435 66 
rect 432 66 435 69 
rect 432 69 435 72 
rect 432 72 435 75 
rect 432 75 435 78 
rect 432 78 435 81 
rect 432 81 435 84 
rect 432 84 435 87 
rect 432 87 435 90 
rect 432 90 435 93 
rect 432 93 435 96 
rect 432 96 435 99 
rect 432 99 435 102 
rect 432 102 435 105 
rect 432 105 435 108 
rect 432 108 435 111 
rect 432 111 435 114 
rect 432 114 435 117 
rect 432 117 435 120 
rect 432 120 435 123 
rect 432 123 435 126 
rect 432 126 435 129 
rect 432 129 435 132 
rect 432 132 435 135 
rect 432 135 435 138 
rect 432 138 435 141 
rect 432 141 435 144 
rect 432 144 435 147 
rect 432 147 435 150 
rect 432 150 435 153 
rect 432 153 435 156 
rect 432 156 435 159 
rect 432 159 435 162 
rect 432 162 435 165 
rect 432 165 435 168 
rect 432 168 435 171 
rect 432 171 435 174 
rect 432 174 435 177 
rect 432 177 435 180 
rect 432 180 435 183 
rect 432 183 435 186 
rect 432 186 435 189 
rect 432 189 435 192 
rect 432 192 435 195 
rect 432 195 435 198 
rect 432 198 435 201 
rect 432 201 435 204 
rect 432 204 435 207 
rect 432 207 435 210 
rect 432 210 435 213 
rect 432 213 435 216 
rect 432 216 435 219 
rect 432 219 435 222 
rect 432 222 435 225 
rect 432 225 435 228 
rect 432 228 435 231 
rect 432 231 435 234 
rect 432 234 435 237 
rect 432 237 435 240 
rect 432 240 435 243 
rect 432 243 435 246 
rect 432 246 435 249 
rect 432 249 435 252 
rect 432 252 435 255 
rect 432 255 435 258 
rect 432 258 435 261 
rect 432 261 435 264 
rect 432 264 435 267 
rect 432 267 435 270 
rect 432 270 435 273 
rect 432 273 435 276 
rect 432 276 435 279 
rect 432 279 435 282 
rect 432 282 435 285 
rect 432 285 435 288 
rect 432 288 435 291 
rect 432 291 435 294 
rect 432 294 435 297 
rect 432 297 435 300 
rect 432 300 435 303 
rect 432 303 435 306 
rect 432 306 435 309 
rect 432 309 435 312 
rect 432 312 435 315 
rect 432 315 435 318 
rect 432 318 435 321 
rect 432 321 435 324 
rect 432 324 435 327 
rect 432 327 435 330 
rect 432 330 435 333 
rect 432 333 435 336 
rect 432 336 435 339 
rect 432 339 435 342 
rect 432 342 435 345 
rect 432 345 435 348 
rect 432 348 435 351 
rect 432 351 435 354 
rect 432 354 435 357 
rect 432 357 435 360 
rect 432 360 435 363 
rect 432 363 435 366 
rect 432 366 435 369 
rect 432 369 435 372 
rect 432 372 435 375 
rect 432 375 435 378 
rect 432 378 435 381 
rect 432 381 435 384 
rect 432 384 435 387 
rect 432 387 435 390 
rect 432 390 435 393 
rect 432 393 435 396 
rect 432 396 435 399 
rect 432 399 435 402 
rect 432 402 435 405 
rect 432 405 435 408 
rect 432 408 435 411 
rect 432 411 435 414 
rect 432 414 435 417 
rect 432 417 435 420 
rect 432 420 435 423 
rect 432 423 435 426 
rect 432 426 435 429 
rect 432 429 435 432 
rect 432 432 435 435 
rect 432 435 435 438 
rect 432 438 435 441 
rect 432 441 435 444 
rect 432 444 435 447 
rect 432 447 435 450 
rect 432 450 435 453 
rect 432 453 435 456 
rect 432 456 435 459 
rect 432 459 435 462 
rect 432 462 435 465 
rect 432 465 435 468 
rect 432 468 435 471 
rect 432 471 435 474 
rect 432 474 435 477 
rect 432 477 435 480 
rect 432 480 435 483 
rect 432 483 435 486 
rect 432 486 435 489 
rect 432 489 435 492 
rect 432 492 435 495 
rect 432 495 435 498 
rect 432 498 435 501 
rect 432 501 435 504 
rect 432 504 435 507 
rect 432 507 435 510 
rect 435 0 438 3 
rect 435 3 438 6 
rect 435 6 438 9 
rect 435 9 438 12 
rect 435 12 438 15 
rect 435 15 438 18 
rect 435 18 438 21 
rect 435 21 438 24 
rect 435 24 438 27 
rect 435 27 438 30 
rect 435 30 438 33 
rect 435 33 438 36 
rect 435 36 438 39 
rect 435 39 438 42 
rect 435 42 438 45 
rect 435 45 438 48 
rect 435 48 438 51 
rect 435 51 438 54 
rect 435 54 438 57 
rect 435 57 438 60 
rect 435 60 438 63 
rect 435 63 438 66 
rect 435 66 438 69 
rect 435 69 438 72 
rect 435 72 438 75 
rect 435 75 438 78 
rect 435 78 438 81 
rect 435 81 438 84 
rect 435 84 438 87 
rect 435 87 438 90 
rect 435 90 438 93 
rect 435 93 438 96 
rect 435 96 438 99 
rect 435 99 438 102 
rect 435 102 438 105 
rect 435 105 438 108 
rect 435 108 438 111 
rect 435 111 438 114 
rect 435 114 438 117 
rect 435 117 438 120 
rect 435 120 438 123 
rect 435 123 438 126 
rect 435 126 438 129 
rect 435 129 438 132 
rect 435 132 438 135 
rect 435 135 438 138 
rect 435 138 438 141 
rect 435 141 438 144 
rect 435 144 438 147 
rect 435 147 438 150 
rect 435 150 438 153 
rect 435 153 438 156 
rect 435 156 438 159 
rect 435 159 438 162 
rect 435 162 438 165 
rect 435 165 438 168 
rect 435 168 438 171 
rect 435 171 438 174 
rect 435 174 438 177 
rect 435 177 438 180 
rect 435 180 438 183 
rect 435 183 438 186 
rect 435 186 438 189 
rect 435 189 438 192 
rect 435 192 438 195 
rect 435 195 438 198 
rect 435 198 438 201 
rect 435 201 438 204 
rect 435 204 438 207 
rect 435 207 438 210 
rect 435 210 438 213 
rect 435 213 438 216 
rect 435 216 438 219 
rect 435 219 438 222 
rect 435 222 438 225 
rect 435 225 438 228 
rect 435 228 438 231 
rect 435 231 438 234 
rect 435 234 438 237 
rect 435 237 438 240 
rect 435 240 438 243 
rect 435 243 438 246 
rect 435 246 438 249 
rect 435 249 438 252 
rect 435 252 438 255 
rect 435 255 438 258 
rect 435 258 438 261 
rect 435 261 438 264 
rect 435 264 438 267 
rect 435 267 438 270 
rect 435 270 438 273 
rect 435 273 438 276 
rect 435 276 438 279 
rect 435 279 438 282 
rect 435 282 438 285 
rect 435 285 438 288 
rect 435 288 438 291 
rect 435 291 438 294 
rect 435 294 438 297 
rect 435 297 438 300 
rect 435 300 438 303 
rect 435 303 438 306 
rect 435 306 438 309 
rect 435 309 438 312 
rect 435 312 438 315 
rect 435 315 438 318 
rect 435 318 438 321 
rect 435 321 438 324 
rect 435 324 438 327 
rect 435 327 438 330 
rect 435 330 438 333 
rect 435 333 438 336 
rect 435 336 438 339 
rect 435 339 438 342 
rect 435 342 438 345 
rect 435 345 438 348 
rect 435 348 438 351 
rect 435 351 438 354 
rect 435 354 438 357 
rect 435 357 438 360 
rect 435 360 438 363 
rect 435 363 438 366 
rect 435 366 438 369 
rect 435 369 438 372 
rect 435 372 438 375 
rect 435 375 438 378 
rect 435 378 438 381 
rect 435 381 438 384 
rect 435 384 438 387 
rect 435 387 438 390 
rect 435 390 438 393 
rect 435 393 438 396 
rect 435 396 438 399 
rect 435 399 438 402 
rect 435 402 438 405 
rect 435 405 438 408 
rect 435 408 438 411 
rect 435 411 438 414 
rect 435 414 438 417 
rect 435 417 438 420 
rect 435 420 438 423 
rect 435 423 438 426 
rect 435 426 438 429 
rect 435 429 438 432 
rect 435 432 438 435 
rect 435 435 438 438 
rect 435 438 438 441 
rect 435 441 438 444 
rect 435 444 438 447 
rect 435 447 438 450 
rect 435 450 438 453 
rect 435 453 438 456 
rect 435 456 438 459 
rect 435 459 438 462 
rect 435 462 438 465 
rect 435 465 438 468 
rect 435 468 438 471 
rect 435 471 438 474 
rect 435 474 438 477 
rect 435 477 438 480 
rect 435 480 438 483 
rect 435 483 438 486 
rect 435 486 438 489 
rect 435 489 438 492 
rect 435 492 438 495 
rect 435 495 438 498 
rect 435 498 438 501 
rect 435 501 438 504 
rect 435 504 438 507 
rect 435 507 438 510 
rect 438 0 441 3 
rect 438 3 441 6 
rect 438 6 441 9 
rect 438 9 441 12 
rect 438 12 441 15 
rect 438 15 441 18 
rect 438 18 441 21 
rect 438 21 441 24 
rect 438 24 441 27 
rect 438 27 441 30 
rect 438 30 441 33 
rect 438 33 441 36 
rect 438 36 441 39 
rect 438 39 441 42 
rect 438 42 441 45 
rect 438 45 441 48 
rect 438 48 441 51 
rect 438 51 441 54 
rect 438 54 441 57 
rect 438 57 441 60 
rect 438 60 441 63 
rect 438 63 441 66 
rect 438 66 441 69 
rect 438 69 441 72 
rect 438 72 441 75 
rect 438 75 441 78 
rect 438 78 441 81 
rect 438 81 441 84 
rect 438 84 441 87 
rect 438 87 441 90 
rect 438 90 441 93 
rect 438 93 441 96 
rect 438 96 441 99 
rect 438 99 441 102 
rect 438 102 441 105 
rect 438 105 441 108 
rect 438 108 441 111 
rect 438 111 441 114 
rect 438 114 441 117 
rect 438 117 441 120 
rect 438 120 441 123 
rect 438 123 441 126 
rect 438 126 441 129 
rect 438 129 441 132 
rect 438 132 441 135 
rect 438 135 441 138 
rect 438 138 441 141 
rect 438 141 441 144 
rect 438 144 441 147 
rect 438 147 441 150 
rect 438 150 441 153 
rect 438 153 441 156 
rect 438 156 441 159 
rect 438 159 441 162 
rect 438 162 441 165 
rect 438 165 441 168 
rect 438 168 441 171 
rect 438 171 441 174 
rect 438 174 441 177 
rect 438 177 441 180 
rect 438 180 441 183 
rect 438 183 441 186 
rect 438 186 441 189 
rect 438 189 441 192 
rect 438 192 441 195 
rect 438 195 441 198 
rect 438 198 441 201 
rect 438 201 441 204 
rect 438 204 441 207 
rect 438 207 441 210 
rect 438 210 441 213 
rect 438 213 441 216 
rect 438 216 441 219 
rect 438 219 441 222 
rect 438 222 441 225 
rect 438 225 441 228 
rect 438 228 441 231 
rect 438 231 441 234 
rect 438 234 441 237 
rect 438 237 441 240 
rect 438 240 441 243 
rect 438 243 441 246 
rect 438 246 441 249 
rect 438 249 441 252 
rect 438 252 441 255 
rect 438 255 441 258 
rect 438 258 441 261 
rect 438 261 441 264 
rect 438 264 441 267 
rect 438 267 441 270 
rect 438 270 441 273 
rect 438 273 441 276 
rect 438 276 441 279 
rect 438 279 441 282 
rect 438 282 441 285 
rect 438 285 441 288 
rect 438 288 441 291 
rect 438 291 441 294 
rect 438 294 441 297 
rect 438 297 441 300 
rect 438 300 441 303 
rect 438 303 441 306 
rect 438 306 441 309 
rect 438 309 441 312 
rect 438 312 441 315 
rect 438 315 441 318 
rect 438 318 441 321 
rect 438 321 441 324 
rect 438 324 441 327 
rect 438 327 441 330 
rect 438 330 441 333 
rect 438 333 441 336 
rect 438 336 441 339 
rect 438 339 441 342 
rect 438 342 441 345 
rect 438 345 441 348 
rect 438 348 441 351 
rect 438 351 441 354 
rect 438 354 441 357 
rect 438 357 441 360 
rect 438 360 441 363 
rect 438 363 441 366 
rect 438 366 441 369 
rect 438 369 441 372 
rect 438 372 441 375 
rect 438 375 441 378 
rect 438 378 441 381 
rect 438 381 441 384 
rect 438 384 441 387 
rect 438 387 441 390 
rect 438 390 441 393 
rect 438 393 441 396 
rect 438 396 441 399 
rect 438 399 441 402 
rect 438 402 441 405 
rect 438 405 441 408 
rect 438 408 441 411 
rect 438 411 441 414 
rect 438 414 441 417 
rect 438 417 441 420 
rect 438 420 441 423 
rect 438 423 441 426 
rect 438 426 441 429 
rect 438 429 441 432 
rect 438 432 441 435 
rect 438 435 441 438 
rect 438 438 441 441 
rect 438 441 441 444 
rect 438 444 441 447 
rect 438 447 441 450 
rect 438 450 441 453 
rect 438 453 441 456 
rect 438 456 441 459 
rect 438 459 441 462 
rect 438 462 441 465 
rect 438 465 441 468 
rect 438 468 441 471 
rect 438 471 441 474 
rect 438 474 441 477 
rect 438 477 441 480 
rect 438 480 441 483 
rect 438 483 441 486 
rect 438 486 441 489 
rect 438 489 441 492 
rect 438 492 441 495 
rect 438 495 441 498 
rect 438 498 441 501 
rect 438 501 441 504 
rect 438 504 441 507 
rect 438 507 441 510 
rect 441 0 444 3 
rect 441 3 444 6 
rect 441 6 444 9 
rect 441 9 444 12 
rect 441 12 444 15 
rect 441 15 444 18 
rect 441 18 444 21 
rect 441 21 444 24 
rect 441 24 444 27 
rect 441 27 444 30 
rect 441 30 444 33 
rect 441 33 444 36 
rect 441 36 444 39 
rect 441 39 444 42 
rect 441 42 444 45 
rect 441 45 444 48 
rect 441 48 444 51 
rect 441 51 444 54 
rect 441 54 444 57 
rect 441 57 444 60 
rect 441 60 444 63 
rect 441 63 444 66 
rect 441 66 444 69 
rect 441 69 444 72 
rect 441 72 444 75 
rect 441 75 444 78 
rect 441 78 444 81 
rect 441 81 444 84 
rect 441 84 444 87 
rect 441 87 444 90 
rect 441 90 444 93 
rect 441 93 444 96 
rect 441 96 444 99 
rect 441 99 444 102 
rect 441 102 444 105 
rect 441 105 444 108 
rect 441 108 444 111 
rect 441 111 444 114 
rect 441 114 444 117 
rect 441 117 444 120 
rect 441 120 444 123 
rect 441 123 444 126 
rect 441 126 444 129 
rect 441 129 444 132 
rect 441 132 444 135 
rect 441 135 444 138 
rect 441 138 444 141 
rect 441 141 444 144 
rect 441 144 444 147 
rect 441 147 444 150 
rect 441 150 444 153 
rect 441 153 444 156 
rect 441 156 444 159 
rect 441 159 444 162 
rect 441 162 444 165 
rect 441 165 444 168 
rect 441 168 444 171 
rect 441 171 444 174 
rect 441 174 444 177 
rect 441 177 444 180 
rect 441 180 444 183 
rect 441 183 444 186 
rect 441 186 444 189 
rect 441 189 444 192 
rect 441 192 444 195 
rect 441 195 444 198 
rect 441 198 444 201 
rect 441 201 444 204 
rect 441 204 444 207 
rect 441 207 444 210 
rect 441 210 444 213 
rect 441 213 444 216 
rect 441 216 444 219 
rect 441 219 444 222 
rect 441 222 444 225 
rect 441 225 444 228 
rect 441 228 444 231 
rect 441 231 444 234 
rect 441 234 444 237 
rect 441 237 444 240 
rect 441 240 444 243 
rect 441 243 444 246 
rect 441 246 444 249 
rect 441 249 444 252 
rect 441 252 444 255 
rect 441 255 444 258 
rect 441 258 444 261 
rect 441 261 444 264 
rect 441 264 444 267 
rect 441 267 444 270 
rect 441 270 444 273 
rect 441 273 444 276 
rect 441 276 444 279 
rect 441 279 444 282 
rect 441 282 444 285 
rect 441 285 444 288 
rect 441 288 444 291 
rect 441 291 444 294 
rect 441 294 444 297 
rect 441 297 444 300 
rect 441 300 444 303 
rect 441 303 444 306 
rect 441 306 444 309 
rect 441 309 444 312 
rect 441 312 444 315 
rect 441 315 444 318 
rect 441 318 444 321 
rect 441 321 444 324 
rect 441 324 444 327 
rect 441 327 444 330 
rect 441 330 444 333 
rect 441 333 444 336 
rect 441 336 444 339 
rect 441 339 444 342 
rect 441 342 444 345 
rect 441 345 444 348 
rect 441 348 444 351 
rect 441 351 444 354 
rect 441 354 444 357 
rect 441 357 444 360 
rect 441 360 444 363 
rect 441 363 444 366 
rect 441 366 444 369 
rect 441 369 444 372 
rect 441 372 444 375 
rect 441 375 444 378 
rect 441 378 444 381 
rect 441 381 444 384 
rect 441 384 444 387 
rect 441 387 444 390 
rect 441 390 444 393 
rect 441 393 444 396 
rect 441 396 444 399 
rect 441 399 444 402 
rect 441 402 444 405 
rect 441 405 444 408 
rect 441 408 444 411 
rect 441 411 444 414 
rect 441 414 444 417 
rect 441 417 444 420 
rect 441 420 444 423 
rect 441 423 444 426 
rect 441 426 444 429 
rect 441 429 444 432 
rect 441 432 444 435 
rect 441 435 444 438 
rect 441 438 444 441 
rect 441 441 444 444 
rect 441 444 444 447 
rect 441 447 444 450 
rect 441 450 444 453 
rect 441 453 444 456 
rect 441 456 444 459 
rect 441 459 444 462 
rect 441 462 444 465 
rect 441 465 444 468 
rect 441 468 444 471 
rect 441 471 444 474 
rect 441 474 444 477 
rect 441 477 444 480 
rect 441 480 444 483 
rect 441 483 444 486 
rect 441 486 444 489 
rect 441 489 444 492 
rect 441 492 444 495 
rect 441 495 444 498 
rect 441 498 444 501 
rect 441 501 444 504 
rect 441 504 444 507 
rect 441 507 444 510 
rect 444 0 447 3 
rect 444 3 447 6 
rect 444 6 447 9 
rect 444 9 447 12 
rect 444 12 447 15 
rect 444 15 447 18 
rect 444 18 447 21 
rect 444 21 447 24 
rect 444 24 447 27 
rect 444 27 447 30 
rect 444 30 447 33 
rect 444 33 447 36 
rect 444 36 447 39 
rect 444 39 447 42 
rect 444 42 447 45 
rect 444 45 447 48 
rect 444 48 447 51 
rect 444 51 447 54 
rect 444 54 447 57 
rect 444 57 447 60 
rect 444 60 447 63 
rect 444 63 447 66 
rect 444 66 447 69 
rect 444 69 447 72 
rect 444 72 447 75 
rect 444 75 447 78 
rect 444 78 447 81 
rect 444 81 447 84 
rect 444 84 447 87 
rect 444 87 447 90 
rect 444 90 447 93 
rect 444 93 447 96 
rect 444 96 447 99 
rect 444 99 447 102 
rect 444 102 447 105 
rect 444 105 447 108 
rect 444 108 447 111 
rect 444 111 447 114 
rect 444 114 447 117 
rect 444 117 447 120 
rect 444 120 447 123 
rect 444 123 447 126 
rect 444 126 447 129 
rect 444 129 447 132 
rect 444 132 447 135 
rect 444 135 447 138 
rect 444 138 447 141 
rect 444 141 447 144 
rect 444 144 447 147 
rect 444 147 447 150 
rect 444 150 447 153 
rect 444 153 447 156 
rect 444 156 447 159 
rect 444 159 447 162 
rect 444 162 447 165 
rect 444 165 447 168 
rect 444 168 447 171 
rect 444 171 447 174 
rect 444 174 447 177 
rect 444 177 447 180 
rect 444 180 447 183 
rect 444 183 447 186 
rect 444 186 447 189 
rect 444 189 447 192 
rect 444 192 447 195 
rect 444 195 447 198 
rect 444 198 447 201 
rect 444 201 447 204 
rect 444 204 447 207 
rect 444 207 447 210 
rect 444 210 447 213 
rect 444 213 447 216 
rect 444 216 447 219 
rect 444 219 447 222 
rect 444 222 447 225 
rect 444 225 447 228 
rect 444 228 447 231 
rect 444 231 447 234 
rect 444 234 447 237 
rect 444 237 447 240 
rect 444 240 447 243 
rect 444 243 447 246 
rect 444 246 447 249 
rect 444 249 447 252 
rect 444 252 447 255 
rect 444 255 447 258 
rect 444 258 447 261 
rect 444 261 447 264 
rect 444 264 447 267 
rect 444 267 447 270 
rect 444 270 447 273 
rect 444 273 447 276 
rect 444 276 447 279 
rect 444 279 447 282 
rect 444 282 447 285 
rect 444 285 447 288 
rect 444 288 447 291 
rect 444 291 447 294 
rect 444 294 447 297 
rect 444 297 447 300 
rect 444 300 447 303 
rect 444 303 447 306 
rect 444 306 447 309 
rect 444 309 447 312 
rect 444 312 447 315 
rect 444 315 447 318 
rect 444 318 447 321 
rect 444 321 447 324 
rect 444 324 447 327 
rect 444 327 447 330 
rect 444 330 447 333 
rect 444 333 447 336 
rect 444 336 447 339 
rect 444 339 447 342 
rect 444 342 447 345 
rect 444 345 447 348 
rect 444 348 447 351 
rect 444 351 447 354 
rect 444 354 447 357 
rect 444 357 447 360 
rect 444 360 447 363 
rect 444 363 447 366 
rect 444 366 447 369 
rect 444 369 447 372 
rect 444 372 447 375 
rect 444 375 447 378 
rect 444 378 447 381 
rect 444 381 447 384 
rect 444 384 447 387 
rect 444 387 447 390 
rect 444 390 447 393 
rect 444 393 447 396 
rect 444 396 447 399 
rect 444 399 447 402 
rect 444 402 447 405 
rect 444 405 447 408 
rect 444 408 447 411 
rect 444 411 447 414 
rect 444 414 447 417 
rect 444 417 447 420 
rect 444 420 447 423 
rect 444 423 447 426 
rect 444 426 447 429 
rect 444 429 447 432 
rect 444 432 447 435 
rect 444 435 447 438 
rect 444 438 447 441 
rect 444 441 447 444 
rect 444 444 447 447 
rect 444 447 447 450 
rect 444 450 447 453 
rect 444 453 447 456 
rect 444 456 447 459 
rect 444 459 447 462 
rect 444 462 447 465 
rect 444 465 447 468 
rect 444 468 447 471 
rect 444 471 447 474 
rect 444 474 447 477 
rect 444 477 447 480 
rect 444 480 447 483 
rect 444 483 447 486 
rect 444 486 447 489 
rect 444 489 447 492 
rect 444 492 447 495 
rect 444 495 447 498 
rect 444 498 447 501 
rect 444 501 447 504 
rect 444 504 447 507 
rect 444 507 447 510 
rect 447 0 450 3 
rect 447 3 450 6 
rect 447 6 450 9 
rect 447 9 450 12 
rect 447 12 450 15 
rect 447 15 450 18 
rect 447 18 450 21 
rect 447 21 450 24 
rect 447 24 450 27 
rect 447 27 450 30 
rect 447 30 450 33 
rect 447 33 450 36 
rect 447 36 450 39 
rect 447 39 450 42 
rect 447 42 450 45 
rect 447 45 450 48 
rect 447 48 450 51 
rect 447 51 450 54 
rect 447 54 450 57 
rect 447 57 450 60 
rect 447 60 450 63 
rect 447 63 450 66 
rect 447 66 450 69 
rect 447 69 450 72 
rect 447 72 450 75 
rect 447 75 450 78 
rect 447 78 450 81 
rect 447 81 450 84 
rect 447 84 450 87 
rect 447 87 450 90 
rect 447 90 450 93 
rect 447 93 450 96 
rect 447 96 450 99 
rect 447 99 450 102 
rect 447 102 450 105 
rect 447 105 450 108 
rect 447 108 450 111 
rect 447 111 450 114 
rect 447 114 450 117 
rect 447 117 450 120 
rect 447 120 450 123 
rect 447 123 450 126 
rect 447 126 450 129 
rect 447 129 450 132 
rect 447 132 450 135 
rect 447 135 450 138 
rect 447 138 450 141 
rect 447 141 450 144 
rect 447 144 450 147 
rect 447 147 450 150 
rect 447 150 450 153 
rect 447 153 450 156 
rect 447 156 450 159 
rect 447 159 450 162 
rect 447 162 450 165 
rect 447 165 450 168 
rect 447 168 450 171 
rect 447 171 450 174 
rect 447 174 450 177 
rect 447 177 450 180 
rect 447 180 450 183 
rect 447 183 450 186 
rect 447 186 450 189 
rect 447 189 450 192 
rect 447 192 450 195 
rect 447 195 450 198 
rect 447 198 450 201 
rect 447 201 450 204 
rect 447 204 450 207 
rect 447 207 450 210 
rect 447 210 450 213 
rect 447 213 450 216 
rect 447 216 450 219 
rect 447 219 450 222 
rect 447 222 450 225 
rect 447 225 450 228 
rect 447 228 450 231 
rect 447 231 450 234 
rect 447 234 450 237 
rect 447 237 450 240 
rect 447 240 450 243 
rect 447 243 450 246 
rect 447 246 450 249 
rect 447 249 450 252 
rect 447 252 450 255 
rect 447 255 450 258 
rect 447 258 450 261 
rect 447 261 450 264 
rect 447 264 450 267 
rect 447 267 450 270 
rect 447 270 450 273 
rect 447 273 450 276 
rect 447 276 450 279 
rect 447 279 450 282 
rect 447 282 450 285 
rect 447 285 450 288 
rect 447 288 450 291 
rect 447 291 450 294 
rect 447 294 450 297 
rect 447 297 450 300 
rect 447 300 450 303 
rect 447 303 450 306 
rect 447 306 450 309 
rect 447 309 450 312 
rect 447 312 450 315 
rect 447 315 450 318 
rect 447 318 450 321 
rect 447 321 450 324 
rect 447 324 450 327 
rect 447 327 450 330 
rect 447 330 450 333 
rect 447 333 450 336 
rect 447 336 450 339 
rect 447 339 450 342 
rect 447 342 450 345 
rect 447 345 450 348 
rect 447 348 450 351 
rect 447 351 450 354 
rect 447 354 450 357 
rect 447 357 450 360 
rect 447 360 450 363 
rect 447 363 450 366 
rect 447 366 450 369 
rect 447 369 450 372 
rect 447 372 450 375 
rect 447 375 450 378 
rect 447 378 450 381 
rect 447 381 450 384 
rect 447 384 450 387 
rect 447 387 450 390 
rect 447 390 450 393 
rect 447 393 450 396 
rect 447 396 450 399 
rect 447 399 450 402 
rect 447 402 450 405 
rect 447 405 450 408 
rect 447 408 450 411 
rect 447 411 450 414 
rect 447 414 450 417 
rect 447 417 450 420 
rect 447 420 450 423 
rect 447 423 450 426 
rect 447 426 450 429 
rect 447 429 450 432 
rect 447 432 450 435 
rect 447 435 450 438 
rect 447 438 450 441 
rect 447 441 450 444 
rect 447 444 450 447 
rect 447 447 450 450 
rect 447 450 450 453 
rect 447 453 450 456 
rect 447 456 450 459 
rect 447 459 450 462 
rect 447 462 450 465 
rect 447 465 450 468 
rect 447 468 450 471 
rect 447 471 450 474 
rect 447 474 450 477 
rect 447 477 450 480 
rect 447 480 450 483 
rect 447 483 450 486 
rect 447 486 450 489 
rect 447 489 450 492 
rect 447 492 450 495 
rect 447 495 450 498 
rect 447 498 450 501 
rect 447 501 450 504 
rect 447 504 450 507 
rect 447 507 450 510 
rect 450 0 453 3 
rect 450 3 453 6 
rect 450 6 453 9 
rect 450 9 453 12 
rect 450 12 453 15 
rect 450 15 453 18 
rect 450 18 453 21 
rect 450 21 453 24 
rect 450 24 453 27 
rect 450 27 453 30 
rect 450 30 453 33 
rect 450 33 453 36 
rect 450 36 453 39 
rect 450 39 453 42 
rect 450 42 453 45 
rect 450 45 453 48 
rect 450 48 453 51 
rect 450 51 453 54 
rect 450 54 453 57 
rect 450 57 453 60 
rect 450 60 453 63 
rect 450 63 453 66 
rect 450 66 453 69 
rect 450 69 453 72 
rect 450 72 453 75 
rect 450 75 453 78 
rect 450 78 453 81 
rect 450 81 453 84 
rect 450 84 453 87 
rect 450 87 453 90 
rect 450 90 453 93 
rect 450 93 453 96 
rect 450 96 453 99 
rect 450 99 453 102 
rect 450 102 453 105 
rect 450 105 453 108 
rect 450 108 453 111 
rect 450 111 453 114 
rect 450 114 453 117 
rect 450 117 453 120 
rect 450 120 453 123 
rect 450 123 453 126 
rect 450 126 453 129 
rect 450 129 453 132 
rect 450 132 453 135 
rect 450 135 453 138 
rect 450 138 453 141 
rect 450 141 453 144 
rect 450 144 453 147 
rect 450 147 453 150 
rect 450 150 453 153 
rect 450 153 453 156 
rect 450 156 453 159 
rect 450 159 453 162 
rect 450 162 453 165 
rect 450 165 453 168 
rect 450 168 453 171 
rect 450 171 453 174 
rect 450 174 453 177 
rect 450 177 453 180 
rect 450 180 453 183 
rect 450 183 453 186 
rect 450 186 453 189 
rect 450 189 453 192 
rect 450 192 453 195 
rect 450 195 453 198 
rect 450 198 453 201 
rect 450 201 453 204 
rect 450 204 453 207 
rect 450 207 453 210 
rect 450 210 453 213 
rect 450 213 453 216 
rect 450 216 453 219 
rect 450 219 453 222 
rect 450 222 453 225 
rect 450 225 453 228 
rect 450 228 453 231 
rect 450 231 453 234 
rect 450 234 453 237 
rect 450 237 453 240 
rect 450 240 453 243 
rect 450 243 453 246 
rect 450 246 453 249 
rect 450 249 453 252 
rect 450 252 453 255 
rect 450 255 453 258 
rect 450 258 453 261 
rect 450 261 453 264 
rect 450 264 453 267 
rect 450 267 453 270 
rect 450 270 453 273 
rect 450 273 453 276 
rect 450 276 453 279 
rect 450 279 453 282 
rect 450 282 453 285 
rect 450 285 453 288 
rect 450 288 453 291 
rect 450 291 453 294 
rect 450 294 453 297 
rect 450 297 453 300 
rect 450 300 453 303 
rect 450 303 453 306 
rect 450 306 453 309 
rect 450 309 453 312 
rect 450 312 453 315 
rect 450 315 453 318 
rect 450 318 453 321 
rect 450 321 453 324 
rect 450 324 453 327 
rect 450 327 453 330 
rect 450 330 453 333 
rect 450 333 453 336 
rect 450 336 453 339 
rect 450 339 453 342 
rect 450 342 453 345 
rect 450 345 453 348 
rect 450 348 453 351 
rect 450 351 453 354 
rect 450 354 453 357 
rect 450 357 453 360 
rect 450 360 453 363 
rect 450 363 453 366 
rect 450 366 453 369 
rect 450 369 453 372 
rect 450 372 453 375 
rect 450 375 453 378 
rect 450 378 453 381 
rect 450 381 453 384 
rect 450 384 453 387 
rect 450 387 453 390 
rect 450 390 453 393 
rect 450 393 453 396 
rect 450 396 453 399 
rect 450 399 453 402 
rect 450 402 453 405 
rect 450 405 453 408 
rect 450 408 453 411 
rect 450 411 453 414 
rect 450 414 453 417 
rect 450 417 453 420 
rect 450 420 453 423 
rect 450 423 453 426 
rect 450 426 453 429 
rect 450 429 453 432 
rect 450 432 453 435 
rect 450 435 453 438 
rect 450 438 453 441 
rect 450 441 453 444 
rect 450 444 453 447 
rect 450 447 453 450 
rect 450 450 453 453 
rect 450 453 453 456 
rect 450 456 453 459 
rect 450 459 453 462 
rect 450 462 453 465 
rect 450 465 453 468 
rect 450 468 453 471 
rect 450 471 453 474 
rect 450 474 453 477 
rect 450 477 453 480 
rect 450 480 453 483 
rect 450 483 453 486 
rect 450 486 453 489 
rect 450 489 453 492 
rect 450 492 453 495 
rect 450 495 453 498 
rect 450 498 453 501 
rect 450 501 453 504 
rect 450 504 453 507 
rect 450 507 453 510 
rect 453 0 456 3 
rect 453 3 456 6 
rect 453 6 456 9 
rect 453 9 456 12 
rect 453 12 456 15 
rect 453 15 456 18 
rect 453 18 456 21 
rect 453 21 456 24 
rect 453 24 456 27 
rect 453 27 456 30 
rect 453 30 456 33 
rect 453 33 456 36 
rect 453 36 456 39 
rect 453 39 456 42 
rect 453 42 456 45 
rect 453 45 456 48 
rect 453 48 456 51 
rect 453 51 456 54 
rect 453 54 456 57 
rect 453 57 456 60 
rect 453 60 456 63 
rect 453 63 456 66 
rect 453 66 456 69 
rect 453 69 456 72 
rect 453 72 456 75 
rect 453 75 456 78 
rect 453 78 456 81 
rect 453 81 456 84 
rect 453 84 456 87 
rect 453 87 456 90 
rect 453 90 456 93 
rect 453 93 456 96 
rect 453 96 456 99 
rect 453 99 456 102 
rect 453 102 456 105 
rect 453 105 456 108 
rect 453 108 456 111 
rect 453 111 456 114 
rect 453 114 456 117 
rect 453 117 456 120 
rect 453 120 456 123 
rect 453 123 456 126 
rect 453 126 456 129 
rect 453 129 456 132 
rect 453 132 456 135 
rect 453 135 456 138 
rect 453 138 456 141 
rect 453 141 456 144 
rect 453 144 456 147 
rect 453 147 456 150 
rect 453 150 456 153 
rect 453 153 456 156 
rect 453 156 456 159 
rect 453 159 456 162 
rect 453 162 456 165 
rect 453 165 456 168 
rect 453 168 456 171 
rect 453 171 456 174 
rect 453 174 456 177 
rect 453 177 456 180 
rect 453 180 456 183 
rect 453 183 456 186 
rect 453 186 456 189 
rect 453 189 456 192 
rect 453 192 456 195 
rect 453 195 456 198 
rect 453 198 456 201 
rect 453 201 456 204 
rect 453 204 456 207 
rect 453 207 456 210 
rect 453 210 456 213 
rect 453 213 456 216 
rect 453 216 456 219 
rect 453 219 456 222 
rect 453 222 456 225 
rect 453 225 456 228 
rect 453 228 456 231 
rect 453 231 456 234 
rect 453 234 456 237 
rect 453 237 456 240 
rect 453 240 456 243 
rect 453 243 456 246 
rect 453 246 456 249 
rect 453 249 456 252 
rect 453 252 456 255 
rect 453 255 456 258 
rect 453 258 456 261 
rect 453 261 456 264 
rect 453 264 456 267 
rect 453 267 456 270 
rect 453 270 456 273 
rect 453 273 456 276 
rect 453 276 456 279 
rect 453 279 456 282 
rect 453 282 456 285 
rect 453 285 456 288 
rect 453 288 456 291 
rect 453 291 456 294 
rect 453 294 456 297 
rect 453 297 456 300 
rect 453 300 456 303 
rect 453 303 456 306 
rect 453 306 456 309 
rect 453 309 456 312 
rect 453 312 456 315 
rect 453 315 456 318 
rect 453 318 456 321 
rect 453 321 456 324 
rect 453 324 456 327 
rect 453 327 456 330 
rect 453 330 456 333 
rect 453 333 456 336 
rect 453 336 456 339 
rect 453 339 456 342 
rect 453 342 456 345 
rect 453 345 456 348 
rect 453 348 456 351 
rect 453 351 456 354 
rect 453 354 456 357 
rect 453 357 456 360 
rect 453 360 456 363 
rect 453 363 456 366 
rect 453 366 456 369 
rect 453 369 456 372 
rect 453 372 456 375 
rect 453 375 456 378 
rect 453 378 456 381 
rect 453 381 456 384 
rect 453 384 456 387 
rect 453 387 456 390 
rect 453 390 456 393 
rect 453 393 456 396 
rect 453 396 456 399 
rect 453 399 456 402 
rect 453 402 456 405 
rect 453 405 456 408 
rect 453 408 456 411 
rect 453 411 456 414 
rect 453 414 456 417 
rect 453 417 456 420 
rect 453 420 456 423 
rect 453 423 456 426 
rect 453 426 456 429 
rect 453 429 456 432 
rect 453 432 456 435 
rect 453 435 456 438 
rect 453 438 456 441 
rect 453 441 456 444 
rect 453 444 456 447 
rect 453 447 456 450 
rect 453 450 456 453 
rect 453 453 456 456 
rect 453 456 456 459 
rect 453 459 456 462 
rect 453 462 456 465 
rect 453 465 456 468 
rect 453 468 456 471 
rect 453 471 456 474 
rect 453 474 456 477 
rect 453 477 456 480 
rect 453 480 456 483 
rect 453 483 456 486 
rect 453 486 456 489 
rect 453 489 456 492 
rect 453 492 456 495 
rect 453 495 456 498 
rect 453 498 456 501 
rect 453 501 456 504 
rect 453 504 456 507 
rect 453 507 456 510 
rect 456 0 459 3 
rect 456 3 459 6 
rect 456 6 459 9 
rect 456 9 459 12 
rect 456 12 459 15 
rect 456 15 459 18 
rect 456 18 459 21 
rect 456 21 459 24 
rect 456 24 459 27 
rect 456 27 459 30 
rect 456 30 459 33 
rect 456 33 459 36 
rect 456 36 459 39 
rect 456 39 459 42 
rect 456 42 459 45 
rect 456 45 459 48 
rect 456 48 459 51 
rect 456 51 459 54 
rect 456 54 459 57 
rect 456 57 459 60 
rect 456 60 459 63 
rect 456 63 459 66 
rect 456 66 459 69 
rect 456 69 459 72 
rect 456 72 459 75 
rect 456 75 459 78 
rect 456 78 459 81 
rect 456 81 459 84 
rect 456 84 459 87 
rect 456 87 459 90 
rect 456 90 459 93 
rect 456 93 459 96 
rect 456 96 459 99 
rect 456 99 459 102 
rect 456 102 459 105 
rect 456 105 459 108 
rect 456 108 459 111 
rect 456 111 459 114 
rect 456 114 459 117 
rect 456 117 459 120 
rect 456 120 459 123 
rect 456 123 459 126 
rect 456 126 459 129 
rect 456 129 459 132 
rect 456 132 459 135 
rect 456 135 459 138 
rect 456 138 459 141 
rect 456 141 459 144 
rect 456 144 459 147 
rect 456 147 459 150 
rect 456 150 459 153 
rect 456 153 459 156 
rect 456 156 459 159 
rect 456 159 459 162 
rect 456 162 459 165 
rect 456 165 459 168 
rect 456 168 459 171 
rect 456 171 459 174 
rect 456 174 459 177 
rect 456 177 459 180 
rect 456 180 459 183 
rect 456 183 459 186 
rect 456 186 459 189 
rect 456 189 459 192 
rect 456 192 459 195 
rect 456 195 459 198 
rect 456 198 459 201 
rect 456 201 459 204 
rect 456 204 459 207 
rect 456 207 459 210 
rect 456 210 459 213 
rect 456 213 459 216 
rect 456 216 459 219 
rect 456 219 459 222 
rect 456 222 459 225 
rect 456 225 459 228 
rect 456 228 459 231 
rect 456 231 459 234 
rect 456 234 459 237 
rect 456 237 459 240 
rect 456 240 459 243 
rect 456 243 459 246 
rect 456 246 459 249 
rect 456 249 459 252 
rect 456 252 459 255 
rect 456 255 459 258 
rect 456 258 459 261 
rect 456 261 459 264 
rect 456 264 459 267 
rect 456 267 459 270 
rect 456 270 459 273 
rect 456 273 459 276 
rect 456 276 459 279 
rect 456 279 459 282 
rect 456 282 459 285 
rect 456 285 459 288 
rect 456 288 459 291 
rect 456 291 459 294 
rect 456 294 459 297 
rect 456 297 459 300 
rect 456 300 459 303 
rect 456 303 459 306 
rect 456 306 459 309 
rect 456 309 459 312 
rect 456 312 459 315 
rect 456 315 459 318 
rect 456 318 459 321 
rect 456 321 459 324 
rect 456 324 459 327 
rect 456 327 459 330 
rect 456 330 459 333 
rect 456 333 459 336 
rect 456 336 459 339 
rect 456 339 459 342 
rect 456 342 459 345 
rect 456 345 459 348 
rect 456 348 459 351 
rect 456 351 459 354 
rect 456 354 459 357 
rect 456 357 459 360 
rect 456 360 459 363 
rect 456 363 459 366 
rect 456 366 459 369 
rect 456 369 459 372 
rect 456 372 459 375 
rect 456 375 459 378 
rect 456 378 459 381 
rect 456 381 459 384 
rect 456 384 459 387 
rect 456 387 459 390 
rect 456 390 459 393 
rect 456 393 459 396 
rect 456 396 459 399 
rect 456 399 459 402 
rect 456 402 459 405 
rect 456 405 459 408 
rect 456 408 459 411 
rect 456 411 459 414 
rect 456 414 459 417 
rect 456 417 459 420 
rect 456 420 459 423 
rect 456 423 459 426 
rect 456 426 459 429 
rect 456 429 459 432 
rect 456 432 459 435 
rect 456 435 459 438 
rect 456 438 459 441 
rect 456 441 459 444 
rect 456 444 459 447 
rect 456 447 459 450 
rect 456 450 459 453 
rect 456 453 459 456 
rect 456 456 459 459 
rect 456 459 459 462 
rect 456 462 459 465 
rect 456 465 459 468 
rect 456 468 459 471 
rect 456 471 459 474 
rect 456 474 459 477 
rect 456 477 459 480 
rect 456 480 459 483 
rect 456 483 459 486 
rect 456 486 459 489 
rect 456 489 459 492 
rect 456 492 459 495 
rect 456 495 459 498 
rect 456 498 459 501 
rect 456 501 459 504 
rect 456 504 459 507 
rect 456 507 459 510 
rect 459 0 462 3 
rect 459 3 462 6 
rect 459 6 462 9 
rect 459 9 462 12 
rect 459 12 462 15 
rect 459 15 462 18 
rect 459 18 462 21 
rect 459 21 462 24 
rect 459 24 462 27 
rect 459 27 462 30 
rect 459 30 462 33 
rect 459 33 462 36 
rect 459 36 462 39 
rect 459 39 462 42 
rect 459 42 462 45 
rect 459 45 462 48 
rect 459 48 462 51 
rect 459 51 462 54 
rect 459 54 462 57 
rect 459 57 462 60 
rect 459 60 462 63 
rect 459 63 462 66 
rect 459 66 462 69 
rect 459 69 462 72 
rect 459 72 462 75 
rect 459 75 462 78 
rect 459 78 462 81 
rect 459 81 462 84 
rect 459 84 462 87 
rect 459 87 462 90 
rect 459 90 462 93 
rect 459 93 462 96 
rect 459 96 462 99 
rect 459 99 462 102 
rect 459 102 462 105 
rect 459 105 462 108 
rect 459 108 462 111 
rect 459 111 462 114 
rect 459 114 462 117 
rect 459 117 462 120 
rect 459 120 462 123 
rect 459 123 462 126 
rect 459 126 462 129 
rect 459 129 462 132 
rect 459 132 462 135 
rect 459 135 462 138 
rect 459 138 462 141 
rect 459 141 462 144 
rect 459 144 462 147 
rect 459 147 462 150 
rect 459 150 462 153 
rect 459 153 462 156 
rect 459 156 462 159 
rect 459 159 462 162 
rect 459 162 462 165 
rect 459 165 462 168 
rect 459 168 462 171 
rect 459 171 462 174 
rect 459 174 462 177 
rect 459 177 462 180 
rect 459 180 462 183 
rect 459 183 462 186 
rect 459 186 462 189 
rect 459 189 462 192 
rect 459 192 462 195 
rect 459 195 462 198 
rect 459 198 462 201 
rect 459 201 462 204 
rect 459 204 462 207 
rect 459 207 462 210 
rect 459 210 462 213 
rect 459 213 462 216 
rect 459 216 462 219 
rect 459 219 462 222 
rect 459 222 462 225 
rect 459 225 462 228 
rect 459 228 462 231 
rect 459 231 462 234 
rect 459 234 462 237 
rect 459 237 462 240 
rect 459 240 462 243 
rect 459 243 462 246 
rect 459 246 462 249 
rect 459 249 462 252 
rect 459 252 462 255 
rect 459 255 462 258 
rect 459 258 462 261 
rect 459 261 462 264 
rect 459 264 462 267 
rect 459 267 462 270 
rect 459 270 462 273 
rect 459 273 462 276 
rect 459 276 462 279 
rect 459 279 462 282 
rect 459 282 462 285 
rect 459 285 462 288 
rect 459 288 462 291 
rect 459 291 462 294 
rect 459 294 462 297 
rect 459 297 462 300 
rect 459 300 462 303 
rect 459 303 462 306 
rect 459 306 462 309 
rect 459 309 462 312 
rect 459 312 462 315 
rect 459 315 462 318 
rect 459 318 462 321 
rect 459 321 462 324 
rect 459 324 462 327 
rect 459 327 462 330 
rect 459 330 462 333 
rect 459 333 462 336 
rect 459 336 462 339 
rect 459 339 462 342 
rect 459 342 462 345 
rect 459 345 462 348 
rect 459 348 462 351 
rect 459 351 462 354 
rect 459 354 462 357 
rect 459 357 462 360 
rect 459 360 462 363 
rect 459 363 462 366 
rect 459 366 462 369 
rect 459 369 462 372 
rect 459 372 462 375 
rect 459 375 462 378 
rect 459 378 462 381 
rect 459 381 462 384 
rect 459 384 462 387 
rect 459 387 462 390 
rect 459 390 462 393 
rect 459 393 462 396 
rect 459 396 462 399 
rect 459 399 462 402 
rect 459 402 462 405 
rect 459 405 462 408 
rect 459 408 462 411 
rect 459 411 462 414 
rect 459 414 462 417 
rect 459 417 462 420 
rect 459 420 462 423 
rect 459 423 462 426 
rect 459 426 462 429 
rect 459 429 462 432 
rect 459 432 462 435 
rect 459 435 462 438 
rect 459 438 462 441 
rect 459 441 462 444 
rect 459 444 462 447 
rect 459 447 462 450 
rect 459 450 462 453 
rect 459 453 462 456 
rect 459 456 462 459 
rect 459 459 462 462 
rect 459 462 462 465 
rect 459 465 462 468 
rect 459 468 462 471 
rect 459 471 462 474 
rect 459 474 462 477 
rect 459 477 462 480 
rect 459 480 462 483 
rect 459 483 462 486 
rect 459 486 462 489 
rect 459 489 462 492 
rect 459 492 462 495 
rect 459 495 462 498 
rect 459 498 462 501 
rect 459 501 462 504 
rect 459 504 462 507 
rect 459 507 462 510 
rect 462 0 465 3 
rect 462 3 465 6 
rect 462 6 465 9 
rect 462 9 465 12 
rect 462 12 465 15 
rect 462 15 465 18 
rect 462 18 465 21 
rect 462 21 465 24 
rect 462 24 465 27 
rect 462 27 465 30 
rect 462 30 465 33 
rect 462 33 465 36 
rect 462 36 465 39 
rect 462 39 465 42 
rect 462 42 465 45 
rect 462 45 465 48 
rect 462 48 465 51 
rect 462 51 465 54 
rect 462 54 465 57 
rect 462 57 465 60 
rect 462 60 465 63 
rect 462 63 465 66 
rect 462 66 465 69 
rect 462 69 465 72 
rect 462 72 465 75 
rect 462 75 465 78 
rect 462 78 465 81 
rect 462 81 465 84 
rect 462 84 465 87 
rect 462 87 465 90 
rect 462 90 465 93 
rect 462 93 465 96 
rect 462 96 465 99 
rect 462 99 465 102 
rect 462 102 465 105 
rect 462 105 465 108 
rect 462 108 465 111 
rect 462 111 465 114 
rect 462 114 465 117 
rect 462 117 465 120 
rect 462 120 465 123 
rect 462 123 465 126 
rect 462 126 465 129 
rect 462 129 465 132 
rect 462 132 465 135 
rect 462 135 465 138 
rect 462 138 465 141 
rect 462 141 465 144 
rect 462 144 465 147 
rect 462 147 465 150 
rect 462 150 465 153 
rect 462 153 465 156 
rect 462 156 465 159 
rect 462 159 465 162 
rect 462 162 465 165 
rect 462 165 465 168 
rect 462 168 465 171 
rect 462 171 465 174 
rect 462 174 465 177 
rect 462 177 465 180 
rect 462 180 465 183 
rect 462 183 465 186 
rect 462 186 465 189 
rect 462 189 465 192 
rect 462 192 465 195 
rect 462 195 465 198 
rect 462 198 465 201 
rect 462 201 465 204 
rect 462 204 465 207 
rect 462 207 465 210 
rect 462 210 465 213 
rect 462 213 465 216 
rect 462 216 465 219 
rect 462 219 465 222 
rect 462 222 465 225 
rect 462 225 465 228 
rect 462 228 465 231 
rect 462 231 465 234 
rect 462 234 465 237 
rect 462 237 465 240 
rect 462 240 465 243 
rect 462 243 465 246 
rect 462 246 465 249 
rect 462 249 465 252 
rect 462 252 465 255 
rect 462 255 465 258 
rect 462 258 465 261 
rect 462 261 465 264 
rect 462 264 465 267 
rect 462 267 465 270 
rect 462 270 465 273 
rect 462 273 465 276 
rect 462 276 465 279 
rect 462 279 465 282 
rect 462 282 465 285 
rect 462 285 465 288 
rect 462 288 465 291 
rect 462 291 465 294 
rect 462 294 465 297 
rect 462 297 465 300 
rect 462 300 465 303 
rect 462 303 465 306 
rect 462 306 465 309 
rect 462 309 465 312 
rect 462 312 465 315 
rect 462 315 465 318 
rect 462 318 465 321 
rect 462 321 465 324 
rect 462 324 465 327 
rect 462 327 465 330 
rect 462 330 465 333 
rect 462 333 465 336 
rect 462 336 465 339 
rect 462 339 465 342 
rect 462 342 465 345 
rect 462 345 465 348 
rect 462 348 465 351 
rect 462 351 465 354 
rect 462 354 465 357 
rect 462 357 465 360 
rect 462 360 465 363 
rect 462 363 465 366 
rect 462 366 465 369 
rect 462 369 465 372 
rect 462 372 465 375 
rect 462 375 465 378 
rect 462 378 465 381 
rect 462 381 465 384 
rect 462 384 465 387 
rect 462 387 465 390 
rect 462 390 465 393 
rect 462 393 465 396 
rect 462 396 465 399 
rect 462 399 465 402 
rect 462 402 465 405 
rect 462 405 465 408 
rect 462 408 465 411 
rect 462 411 465 414 
rect 462 414 465 417 
rect 462 417 465 420 
rect 462 420 465 423 
rect 462 423 465 426 
rect 462 426 465 429 
rect 462 429 465 432 
rect 462 432 465 435 
rect 462 435 465 438 
rect 462 438 465 441 
rect 462 441 465 444 
rect 462 444 465 447 
rect 462 447 465 450 
rect 462 450 465 453 
rect 462 453 465 456 
rect 462 456 465 459 
rect 462 459 465 462 
rect 462 462 465 465 
rect 462 465 465 468 
rect 462 468 465 471 
rect 462 471 465 474 
rect 462 474 465 477 
rect 462 477 465 480 
rect 462 480 465 483 
rect 462 483 465 486 
rect 462 486 465 489 
rect 462 489 465 492 
rect 462 492 465 495 
rect 462 495 465 498 
rect 462 498 465 501 
rect 462 501 465 504 
rect 462 504 465 507 
rect 462 507 465 510 
rect 465 0 468 3 
rect 465 3 468 6 
rect 465 6 468 9 
rect 465 9 468 12 
rect 465 12 468 15 
rect 465 15 468 18 
rect 465 18 468 21 
rect 465 21 468 24 
rect 465 24 468 27 
rect 465 27 468 30 
rect 465 30 468 33 
rect 465 33 468 36 
rect 465 36 468 39 
rect 465 39 468 42 
rect 465 42 468 45 
rect 465 45 468 48 
rect 465 48 468 51 
rect 465 51 468 54 
rect 465 54 468 57 
rect 465 57 468 60 
rect 465 60 468 63 
rect 465 63 468 66 
rect 465 66 468 69 
rect 465 69 468 72 
rect 465 72 468 75 
rect 465 75 468 78 
rect 465 78 468 81 
rect 465 81 468 84 
rect 465 84 468 87 
rect 465 87 468 90 
rect 465 90 468 93 
rect 465 93 468 96 
rect 465 96 468 99 
rect 465 99 468 102 
rect 465 102 468 105 
rect 465 105 468 108 
rect 465 108 468 111 
rect 465 111 468 114 
rect 465 114 468 117 
rect 465 117 468 120 
rect 465 120 468 123 
rect 465 123 468 126 
rect 465 126 468 129 
rect 465 129 468 132 
rect 465 132 468 135 
rect 465 135 468 138 
rect 465 138 468 141 
rect 465 141 468 144 
rect 465 144 468 147 
rect 465 147 468 150 
rect 465 150 468 153 
rect 465 153 468 156 
rect 465 156 468 159 
rect 465 159 468 162 
rect 465 162 468 165 
rect 465 165 468 168 
rect 465 168 468 171 
rect 465 171 468 174 
rect 465 174 468 177 
rect 465 177 468 180 
rect 465 180 468 183 
rect 465 183 468 186 
rect 465 186 468 189 
rect 465 189 468 192 
rect 465 192 468 195 
rect 465 195 468 198 
rect 465 198 468 201 
rect 465 201 468 204 
rect 465 204 468 207 
rect 465 207 468 210 
rect 465 210 468 213 
rect 465 213 468 216 
rect 465 216 468 219 
rect 465 219 468 222 
rect 465 222 468 225 
rect 465 225 468 228 
rect 465 228 468 231 
rect 465 231 468 234 
rect 465 234 468 237 
rect 465 237 468 240 
rect 465 240 468 243 
rect 465 243 468 246 
rect 465 246 468 249 
rect 465 249 468 252 
rect 465 252 468 255 
rect 465 255 468 258 
rect 465 258 468 261 
rect 465 261 468 264 
rect 465 264 468 267 
rect 465 267 468 270 
rect 465 270 468 273 
rect 465 273 468 276 
rect 465 276 468 279 
rect 465 279 468 282 
rect 465 282 468 285 
rect 465 285 468 288 
rect 465 288 468 291 
rect 465 291 468 294 
rect 465 294 468 297 
rect 465 297 468 300 
rect 465 300 468 303 
rect 465 303 468 306 
rect 465 306 468 309 
rect 465 309 468 312 
rect 465 312 468 315 
rect 465 315 468 318 
rect 465 318 468 321 
rect 465 321 468 324 
rect 465 324 468 327 
rect 465 327 468 330 
rect 465 330 468 333 
rect 465 333 468 336 
rect 465 336 468 339 
rect 465 339 468 342 
rect 465 342 468 345 
rect 465 345 468 348 
rect 465 348 468 351 
rect 465 351 468 354 
rect 465 354 468 357 
rect 465 357 468 360 
rect 465 360 468 363 
rect 465 363 468 366 
rect 465 366 468 369 
rect 465 369 468 372 
rect 465 372 468 375 
rect 465 375 468 378 
rect 465 378 468 381 
rect 465 381 468 384 
rect 465 384 468 387 
rect 465 387 468 390 
rect 465 390 468 393 
rect 465 393 468 396 
rect 465 396 468 399 
rect 465 399 468 402 
rect 465 402 468 405 
rect 465 405 468 408 
rect 465 408 468 411 
rect 465 411 468 414 
rect 465 414 468 417 
rect 465 417 468 420 
rect 465 420 468 423 
rect 465 423 468 426 
rect 465 426 468 429 
rect 465 429 468 432 
rect 465 432 468 435 
rect 465 435 468 438 
rect 465 438 468 441 
rect 465 441 468 444 
rect 465 444 468 447 
rect 465 447 468 450 
rect 465 450 468 453 
rect 465 453 468 456 
rect 465 456 468 459 
rect 465 459 468 462 
rect 465 462 468 465 
rect 465 465 468 468 
rect 465 468 468 471 
rect 465 471 468 474 
rect 465 474 468 477 
rect 465 477 468 480 
rect 465 480 468 483 
rect 465 483 468 486 
rect 465 486 468 489 
rect 465 489 468 492 
rect 465 492 468 495 
rect 465 495 468 498 
rect 465 498 468 501 
rect 465 501 468 504 
rect 465 504 468 507 
rect 465 507 468 510 
rect 468 0 471 3 
rect 468 3 471 6 
rect 468 6 471 9 
rect 468 9 471 12 
rect 468 12 471 15 
rect 468 15 471 18 
rect 468 18 471 21 
rect 468 21 471 24 
rect 468 24 471 27 
rect 468 27 471 30 
rect 468 30 471 33 
rect 468 33 471 36 
rect 468 36 471 39 
rect 468 39 471 42 
rect 468 42 471 45 
rect 468 45 471 48 
rect 468 48 471 51 
rect 468 51 471 54 
rect 468 54 471 57 
rect 468 57 471 60 
rect 468 60 471 63 
rect 468 63 471 66 
rect 468 66 471 69 
rect 468 69 471 72 
rect 468 72 471 75 
rect 468 75 471 78 
rect 468 78 471 81 
rect 468 81 471 84 
rect 468 84 471 87 
rect 468 87 471 90 
rect 468 90 471 93 
rect 468 93 471 96 
rect 468 96 471 99 
rect 468 99 471 102 
rect 468 102 471 105 
rect 468 105 471 108 
rect 468 108 471 111 
rect 468 111 471 114 
rect 468 114 471 117 
rect 468 117 471 120 
rect 468 120 471 123 
rect 468 123 471 126 
rect 468 126 471 129 
rect 468 129 471 132 
rect 468 132 471 135 
rect 468 135 471 138 
rect 468 138 471 141 
rect 468 141 471 144 
rect 468 144 471 147 
rect 468 147 471 150 
rect 468 150 471 153 
rect 468 153 471 156 
rect 468 156 471 159 
rect 468 159 471 162 
rect 468 162 471 165 
rect 468 165 471 168 
rect 468 168 471 171 
rect 468 171 471 174 
rect 468 174 471 177 
rect 468 177 471 180 
rect 468 180 471 183 
rect 468 183 471 186 
rect 468 186 471 189 
rect 468 189 471 192 
rect 468 192 471 195 
rect 468 195 471 198 
rect 468 198 471 201 
rect 468 201 471 204 
rect 468 204 471 207 
rect 468 207 471 210 
rect 468 210 471 213 
rect 468 213 471 216 
rect 468 216 471 219 
rect 468 219 471 222 
rect 468 222 471 225 
rect 468 225 471 228 
rect 468 228 471 231 
rect 468 231 471 234 
rect 468 234 471 237 
rect 468 237 471 240 
rect 468 240 471 243 
rect 468 243 471 246 
rect 468 246 471 249 
rect 468 249 471 252 
rect 468 252 471 255 
rect 468 255 471 258 
rect 468 258 471 261 
rect 468 261 471 264 
rect 468 264 471 267 
rect 468 267 471 270 
rect 468 270 471 273 
rect 468 273 471 276 
rect 468 276 471 279 
rect 468 279 471 282 
rect 468 282 471 285 
rect 468 285 471 288 
rect 468 288 471 291 
rect 468 291 471 294 
rect 468 294 471 297 
rect 468 297 471 300 
rect 468 300 471 303 
rect 468 303 471 306 
rect 468 306 471 309 
rect 468 309 471 312 
rect 468 312 471 315 
rect 468 315 471 318 
rect 468 318 471 321 
rect 468 321 471 324 
rect 468 324 471 327 
rect 468 327 471 330 
rect 468 330 471 333 
rect 468 333 471 336 
rect 468 336 471 339 
rect 468 339 471 342 
rect 468 342 471 345 
rect 468 345 471 348 
rect 468 348 471 351 
rect 468 351 471 354 
rect 468 354 471 357 
rect 468 357 471 360 
rect 468 360 471 363 
rect 468 363 471 366 
rect 468 366 471 369 
rect 468 369 471 372 
rect 468 372 471 375 
rect 468 375 471 378 
rect 468 378 471 381 
rect 468 381 471 384 
rect 468 384 471 387 
rect 468 387 471 390 
rect 468 390 471 393 
rect 468 393 471 396 
rect 468 396 471 399 
rect 468 399 471 402 
rect 468 402 471 405 
rect 468 405 471 408 
rect 468 408 471 411 
rect 468 411 471 414 
rect 468 414 471 417 
rect 468 417 471 420 
rect 468 420 471 423 
rect 468 423 471 426 
rect 468 426 471 429 
rect 468 429 471 432 
rect 468 432 471 435 
rect 468 435 471 438 
rect 468 438 471 441 
rect 468 441 471 444 
rect 468 444 471 447 
rect 468 447 471 450 
rect 468 450 471 453 
rect 468 453 471 456 
rect 468 456 471 459 
rect 468 459 471 462 
rect 468 462 471 465 
rect 468 465 471 468 
rect 468 468 471 471 
rect 468 471 471 474 
rect 468 474 471 477 
rect 468 477 471 480 
rect 468 480 471 483 
rect 468 483 471 486 
rect 468 486 471 489 
rect 468 489 471 492 
rect 468 492 471 495 
rect 468 495 471 498 
rect 468 498 471 501 
rect 468 501 471 504 
rect 468 504 471 507 
rect 468 507 471 510 
rect 471 0 474 3 
rect 471 3 474 6 
rect 471 6 474 9 
rect 471 9 474 12 
rect 471 12 474 15 
rect 471 15 474 18 
rect 471 18 474 21 
rect 471 21 474 24 
rect 471 24 474 27 
rect 471 27 474 30 
rect 471 30 474 33 
rect 471 33 474 36 
rect 471 36 474 39 
rect 471 39 474 42 
rect 471 42 474 45 
rect 471 45 474 48 
rect 471 48 474 51 
rect 471 51 474 54 
rect 471 54 474 57 
rect 471 57 474 60 
rect 471 60 474 63 
rect 471 63 474 66 
rect 471 66 474 69 
rect 471 69 474 72 
rect 471 72 474 75 
rect 471 75 474 78 
rect 471 78 474 81 
rect 471 81 474 84 
rect 471 84 474 87 
rect 471 87 474 90 
rect 471 90 474 93 
rect 471 93 474 96 
rect 471 96 474 99 
rect 471 99 474 102 
rect 471 102 474 105 
rect 471 105 474 108 
rect 471 108 474 111 
rect 471 111 474 114 
rect 471 114 474 117 
rect 471 117 474 120 
rect 471 120 474 123 
rect 471 123 474 126 
rect 471 126 474 129 
rect 471 129 474 132 
rect 471 132 474 135 
rect 471 135 474 138 
rect 471 138 474 141 
rect 471 141 474 144 
rect 471 144 474 147 
rect 471 147 474 150 
rect 471 150 474 153 
rect 471 153 474 156 
rect 471 156 474 159 
rect 471 159 474 162 
rect 471 162 474 165 
rect 471 165 474 168 
rect 471 168 474 171 
rect 471 171 474 174 
rect 471 174 474 177 
rect 471 177 474 180 
rect 471 180 474 183 
rect 471 183 474 186 
rect 471 186 474 189 
rect 471 189 474 192 
rect 471 192 474 195 
rect 471 195 474 198 
rect 471 198 474 201 
rect 471 201 474 204 
rect 471 204 474 207 
rect 471 207 474 210 
rect 471 210 474 213 
rect 471 213 474 216 
rect 471 216 474 219 
rect 471 219 474 222 
rect 471 222 474 225 
rect 471 225 474 228 
rect 471 228 474 231 
rect 471 231 474 234 
rect 471 234 474 237 
rect 471 237 474 240 
rect 471 240 474 243 
rect 471 243 474 246 
rect 471 246 474 249 
rect 471 249 474 252 
rect 471 252 474 255 
rect 471 255 474 258 
rect 471 258 474 261 
rect 471 261 474 264 
rect 471 264 474 267 
rect 471 267 474 270 
rect 471 270 474 273 
rect 471 273 474 276 
rect 471 276 474 279 
rect 471 279 474 282 
rect 471 282 474 285 
rect 471 285 474 288 
rect 471 288 474 291 
rect 471 291 474 294 
rect 471 294 474 297 
rect 471 297 474 300 
rect 471 300 474 303 
rect 471 303 474 306 
rect 471 306 474 309 
rect 471 309 474 312 
rect 471 312 474 315 
rect 471 315 474 318 
rect 471 318 474 321 
rect 471 321 474 324 
rect 471 324 474 327 
rect 471 327 474 330 
rect 471 330 474 333 
rect 471 333 474 336 
rect 471 336 474 339 
rect 471 339 474 342 
rect 471 342 474 345 
rect 471 345 474 348 
rect 471 348 474 351 
rect 471 351 474 354 
rect 471 354 474 357 
rect 471 357 474 360 
rect 471 360 474 363 
rect 471 363 474 366 
rect 471 366 474 369 
rect 471 369 474 372 
rect 471 372 474 375 
rect 471 375 474 378 
rect 471 378 474 381 
rect 471 381 474 384 
rect 471 384 474 387 
rect 471 387 474 390 
rect 471 390 474 393 
rect 471 393 474 396 
rect 471 396 474 399 
rect 471 399 474 402 
rect 471 402 474 405 
rect 471 405 474 408 
rect 471 408 474 411 
rect 471 411 474 414 
rect 471 414 474 417 
rect 471 417 474 420 
rect 471 420 474 423 
rect 471 423 474 426 
rect 471 426 474 429 
rect 471 429 474 432 
rect 471 432 474 435 
rect 471 435 474 438 
rect 471 438 474 441 
rect 471 441 474 444 
rect 471 444 474 447 
rect 471 447 474 450 
rect 471 450 474 453 
rect 471 453 474 456 
rect 471 456 474 459 
rect 471 459 474 462 
rect 471 462 474 465 
rect 471 465 474 468 
rect 471 468 474 471 
rect 471 471 474 474 
rect 471 474 474 477 
rect 471 477 474 480 
rect 471 480 474 483 
rect 471 483 474 486 
rect 471 486 474 489 
rect 471 489 474 492 
rect 471 492 474 495 
rect 471 495 474 498 
rect 471 498 474 501 
rect 471 501 474 504 
rect 471 504 474 507 
rect 471 507 474 510 
rect 474 0 477 3 
rect 474 3 477 6 
rect 474 6 477 9 
rect 474 9 477 12 
rect 474 12 477 15 
rect 474 15 477 18 
rect 474 18 477 21 
rect 474 21 477 24 
rect 474 24 477 27 
rect 474 27 477 30 
rect 474 30 477 33 
rect 474 33 477 36 
rect 474 36 477 39 
rect 474 39 477 42 
rect 474 42 477 45 
rect 474 45 477 48 
rect 474 48 477 51 
rect 474 51 477 54 
rect 474 54 477 57 
rect 474 57 477 60 
rect 474 60 477 63 
rect 474 63 477 66 
rect 474 66 477 69 
rect 474 69 477 72 
rect 474 72 477 75 
rect 474 75 477 78 
rect 474 78 477 81 
rect 474 81 477 84 
rect 474 84 477 87 
rect 474 87 477 90 
rect 474 90 477 93 
rect 474 93 477 96 
rect 474 96 477 99 
rect 474 99 477 102 
rect 474 102 477 105 
rect 474 105 477 108 
rect 474 108 477 111 
rect 474 111 477 114 
rect 474 114 477 117 
rect 474 117 477 120 
rect 474 120 477 123 
rect 474 123 477 126 
rect 474 126 477 129 
rect 474 129 477 132 
rect 474 132 477 135 
rect 474 135 477 138 
rect 474 138 477 141 
rect 474 141 477 144 
rect 474 144 477 147 
rect 474 147 477 150 
rect 474 150 477 153 
rect 474 153 477 156 
rect 474 156 477 159 
rect 474 159 477 162 
rect 474 162 477 165 
rect 474 165 477 168 
rect 474 168 477 171 
rect 474 171 477 174 
rect 474 174 477 177 
rect 474 177 477 180 
rect 474 180 477 183 
rect 474 183 477 186 
rect 474 186 477 189 
rect 474 189 477 192 
rect 474 192 477 195 
rect 474 195 477 198 
rect 474 198 477 201 
rect 474 201 477 204 
rect 474 204 477 207 
rect 474 207 477 210 
rect 474 210 477 213 
rect 474 213 477 216 
rect 474 216 477 219 
rect 474 219 477 222 
rect 474 222 477 225 
rect 474 225 477 228 
rect 474 228 477 231 
rect 474 231 477 234 
rect 474 234 477 237 
rect 474 237 477 240 
rect 474 240 477 243 
rect 474 243 477 246 
rect 474 246 477 249 
rect 474 249 477 252 
rect 474 252 477 255 
rect 474 255 477 258 
rect 474 258 477 261 
rect 474 261 477 264 
rect 474 264 477 267 
rect 474 267 477 270 
rect 474 270 477 273 
rect 474 273 477 276 
rect 474 276 477 279 
rect 474 279 477 282 
rect 474 282 477 285 
rect 474 285 477 288 
rect 474 288 477 291 
rect 474 291 477 294 
rect 474 294 477 297 
rect 474 297 477 300 
rect 474 300 477 303 
rect 474 303 477 306 
rect 474 306 477 309 
rect 474 309 477 312 
rect 474 312 477 315 
rect 474 315 477 318 
rect 474 318 477 321 
rect 474 321 477 324 
rect 474 324 477 327 
rect 474 327 477 330 
rect 474 330 477 333 
rect 474 333 477 336 
rect 474 336 477 339 
rect 474 339 477 342 
rect 474 342 477 345 
rect 474 345 477 348 
rect 474 348 477 351 
rect 474 351 477 354 
rect 474 354 477 357 
rect 474 357 477 360 
rect 474 360 477 363 
rect 474 363 477 366 
rect 474 366 477 369 
rect 474 369 477 372 
rect 474 372 477 375 
rect 474 375 477 378 
rect 474 378 477 381 
rect 474 381 477 384 
rect 474 384 477 387 
rect 474 387 477 390 
rect 474 390 477 393 
rect 474 393 477 396 
rect 474 396 477 399 
rect 474 399 477 402 
rect 474 402 477 405 
rect 474 405 477 408 
rect 474 408 477 411 
rect 474 411 477 414 
rect 474 414 477 417 
rect 474 417 477 420 
rect 474 420 477 423 
rect 474 423 477 426 
rect 474 426 477 429 
rect 474 429 477 432 
rect 474 432 477 435 
rect 474 435 477 438 
rect 474 438 477 441 
rect 474 441 477 444 
rect 474 444 477 447 
rect 474 447 477 450 
rect 474 450 477 453 
rect 474 453 477 456 
rect 474 456 477 459 
rect 474 459 477 462 
rect 474 462 477 465 
rect 474 465 477 468 
rect 474 468 477 471 
rect 474 471 477 474 
rect 474 474 477 477 
rect 474 477 477 480 
rect 474 480 477 483 
rect 474 483 477 486 
rect 474 486 477 489 
rect 474 489 477 492 
rect 474 492 477 495 
rect 474 495 477 498 
rect 474 498 477 501 
rect 474 501 477 504 
rect 474 504 477 507 
rect 474 507 477 510 
rect 477 0 480 3 
rect 477 3 480 6 
rect 477 6 480 9 
rect 477 9 480 12 
rect 477 12 480 15 
rect 477 15 480 18 
rect 477 18 480 21 
rect 477 21 480 24 
rect 477 24 480 27 
rect 477 27 480 30 
rect 477 30 480 33 
rect 477 33 480 36 
rect 477 36 480 39 
rect 477 39 480 42 
rect 477 42 480 45 
rect 477 45 480 48 
rect 477 48 480 51 
rect 477 51 480 54 
rect 477 54 480 57 
rect 477 57 480 60 
rect 477 60 480 63 
rect 477 63 480 66 
rect 477 66 480 69 
rect 477 69 480 72 
rect 477 72 480 75 
rect 477 75 480 78 
rect 477 78 480 81 
rect 477 81 480 84 
rect 477 84 480 87 
rect 477 87 480 90 
rect 477 90 480 93 
rect 477 93 480 96 
rect 477 96 480 99 
rect 477 99 480 102 
rect 477 102 480 105 
rect 477 105 480 108 
rect 477 108 480 111 
rect 477 111 480 114 
rect 477 114 480 117 
rect 477 117 480 120 
rect 477 120 480 123 
rect 477 123 480 126 
rect 477 126 480 129 
rect 477 129 480 132 
rect 477 132 480 135 
rect 477 135 480 138 
rect 477 138 480 141 
rect 477 141 480 144 
rect 477 144 480 147 
rect 477 147 480 150 
rect 477 150 480 153 
rect 477 153 480 156 
rect 477 156 480 159 
rect 477 159 480 162 
rect 477 162 480 165 
rect 477 165 480 168 
rect 477 168 480 171 
rect 477 171 480 174 
rect 477 174 480 177 
rect 477 177 480 180 
rect 477 180 480 183 
rect 477 183 480 186 
rect 477 186 480 189 
rect 477 189 480 192 
rect 477 192 480 195 
rect 477 195 480 198 
rect 477 198 480 201 
rect 477 201 480 204 
rect 477 204 480 207 
rect 477 207 480 210 
rect 477 210 480 213 
rect 477 213 480 216 
rect 477 216 480 219 
rect 477 219 480 222 
rect 477 222 480 225 
rect 477 225 480 228 
rect 477 228 480 231 
rect 477 231 480 234 
rect 477 234 480 237 
rect 477 237 480 240 
rect 477 240 480 243 
rect 477 243 480 246 
rect 477 246 480 249 
rect 477 249 480 252 
rect 477 252 480 255 
rect 477 255 480 258 
rect 477 258 480 261 
rect 477 261 480 264 
rect 477 264 480 267 
rect 477 267 480 270 
rect 477 270 480 273 
rect 477 273 480 276 
rect 477 276 480 279 
rect 477 279 480 282 
rect 477 282 480 285 
rect 477 285 480 288 
rect 477 288 480 291 
rect 477 291 480 294 
rect 477 294 480 297 
rect 477 297 480 300 
rect 477 300 480 303 
rect 477 303 480 306 
rect 477 306 480 309 
rect 477 309 480 312 
rect 477 312 480 315 
rect 477 315 480 318 
rect 477 318 480 321 
rect 477 321 480 324 
rect 477 324 480 327 
rect 477 327 480 330 
rect 477 330 480 333 
rect 477 333 480 336 
rect 477 336 480 339 
rect 477 339 480 342 
rect 477 342 480 345 
rect 477 345 480 348 
rect 477 348 480 351 
rect 477 351 480 354 
rect 477 354 480 357 
rect 477 357 480 360 
rect 477 360 480 363 
rect 477 363 480 366 
rect 477 366 480 369 
rect 477 369 480 372 
rect 477 372 480 375 
rect 477 375 480 378 
rect 477 378 480 381 
rect 477 381 480 384 
rect 477 384 480 387 
rect 477 387 480 390 
rect 477 390 480 393 
rect 477 393 480 396 
rect 477 396 480 399 
rect 477 399 480 402 
rect 477 402 480 405 
rect 477 405 480 408 
rect 477 408 480 411 
rect 477 411 480 414 
rect 477 414 480 417 
rect 477 417 480 420 
rect 477 420 480 423 
rect 477 423 480 426 
rect 477 426 480 429 
rect 477 429 480 432 
rect 477 432 480 435 
rect 477 435 480 438 
rect 477 438 480 441 
rect 477 441 480 444 
rect 477 444 480 447 
rect 477 447 480 450 
rect 477 450 480 453 
rect 477 453 480 456 
rect 477 456 480 459 
rect 477 459 480 462 
rect 477 462 480 465 
rect 477 465 480 468 
rect 477 468 480 471 
rect 477 471 480 474 
rect 477 474 480 477 
rect 477 477 480 480 
rect 477 480 480 483 
rect 477 483 480 486 
rect 477 486 480 489 
rect 477 489 480 492 
rect 477 492 480 495 
rect 477 495 480 498 
rect 477 498 480 501 
rect 477 501 480 504 
rect 477 504 480 507 
rect 477 507 480 510 
rect 480 0 483 3 
rect 480 3 483 6 
rect 480 6 483 9 
rect 480 9 483 12 
rect 480 12 483 15 
rect 480 15 483 18 
rect 480 18 483 21 
rect 480 21 483 24 
rect 480 24 483 27 
rect 480 27 483 30 
rect 480 30 483 33 
rect 480 33 483 36 
rect 480 36 483 39 
rect 480 39 483 42 
rect 480 42 483 45 
rect 480 45 483 48 
rect 480 48 483 51 
rect 480 51 483 54 
rect 480 54 483 57 
rect 480 57 483 60 
rect 480 60 483 63 
rect 480 63 483 66 
rect 480 66 483 69 
rect 480 69 483 72 
rect 480 72 483 75 
rect 480 75 483 78 
rect 480 78 483 81 
rect 480 81 483 84 
rect 480 84 483 87 
rect 480 87 483 90 
rect 480 90 483 93 
rect 480 93 483 96 
rect 480 96 483 99 
rect 480 99 483 102 
rect 480 102 483 105 
rect 480 105 483 108 
rect 480 108 483 111 
rect 480 111 483 114 
rect 480 114 483 117 
rect 480 117 483 120 
rect 480 120 483 123 
rect 480 123 483 126 
rect 480 126 483 129 
rect 480 129 483 132 
rect 480 132 483 135 
rect 480 135 483 138 
rect 480 138 483 141 
rect 480 141 483 144 
rect 480 144 483 147 
rect 480 147 483 150 
rect 480 150 483 153 
rect 480 153 483 156 
rect 480 156 483 159 
rect 480 159 483 162 
rect 480 162 483 165 
rect 480 165 483 168 
rect 480 168 483 171 
rect 480 171 483 174 
rect 480 174 483 177 
rect 480 177 483 180 
rect 480 180 483 183 
rect 480 183 483 186 
rect 480 186 483 189 
rect 480 189 483 192 
rect 480 192 483 195 
rect 480 195 483 198 
rect 480 198 483 201 
rect 480 201 483 204 
rect 480 204 483 207 
rect 480 207 483 210 
rect 480 210 483 213 
rect 480 213 483 216 
rect 480 216 483 219 
rect 480 219 483 222 
rect 480 222 483 225 
rect 480 225 483 228 
rect 480 228 483 231 
rect 480 231 483 234 
rect 480 234 483 237 
rect 480 237 483 240 
rect 480 240 483 243 
rect 480 243 483 246 
rect 480 246 483 249 
rect 480 249 483 252 
rect 480 252 483 255 
rect 480 255 483 258 
rect 480 258 483 261 
rect 480 261 483 264 
rect 480 264 483 267 
rect 480 267 483 270 
rect 480 270 483 273 
rect 480 273 483 276 
rect 480 276 483 279 
rect 480 279 483 282 
rect 480 282 483 285 
rect 480 285 483 288 
rect 480 288 483 291 
rect 480 291 483 294 
rect 480 294 483 297 
rect 480 297 483 300 
rect 480 300 483 303 
rect 480 303 483 306 
rect 480 306 483 309 
rect 480 309 483 312 
rect 480 312 483 315 
rect 480 315 483 318 
rect 480 318 483 321 
rect 480 321 483 324 
rect 480 324 483 327 
rect 480 327 483 330 
rect 480 330 483 333 
rect 480 333 483 336 
rect 480 336 483 339 
rect 480 339 483 342 
rect 480 342 483 345 
rect 480 345 483 348 
rect 480 348 483 351 
rect 480 351 483 354 
rect 480 354 483 357 
rect 480 357 483 360 
rect 480 360 483 363 
rect 480 363 483 366 
rect 480 366 483 369 
rect 480 369 483 372 
rect 480 372 483 375 
rect 480 375 483 378 
rect 480 378 483 381 
rect 480 381 483 384 
rect 480 384 483 387 
rect 480 387 483 390 
rect 480 390 483 393 
rect 480 393 483 396 
rect 480 396 483 399 
rect 480 399 483 402 
rect 480 402 483 405 
rect 480 405 483 408 
rect 480 408 483 411 
rect 480 411 483 414 
rect 480 414 483 417 
rect 480 417 483 420 
rect 480 420 483 423 
rect 480 423 483 426 
rect 480 426 483 429 
rect 480 429 483 432 
rect 480 432 483 435 
rect 480 435 483 438 
rect 480 438 483 441 
rect 480 441 483 444 
rect 480 444 483 447 
rect 480 447 483 450 
rect 480 450 483 453 
rect 480 453 483 456 
rect 480 456 483 459 
rect 480 459 483 462 
rect 480 462 483 465 
rect 480 465 483 468 
rect 480 468 483 471 
rect 480 471 483 474 
rect 480 474 483 477 
rect 480 477 483 480 
rect 480 480 483 483 
rect 480 483 483 486 
rect 480 486 483 489 
rect 480 489 483 492 
rect 480 492 483 495 
rect 480 495 483 498 
rect 480 498 483 501 
rect 480 501 483 504 
rect 480 504 483 507 
rect 480 507 483 510 
rect 483 0 486 3 
rect 483 3 486 6 
rect 483 6 486 9 
rect 483 9 486 12 
rect 483 12 486 15 
rect 483 15 486 18 
rect 483 18 486 21 
rect 483 21 486 24 
rect 483 24 486 27 
rect 483 27 486 30 
rect 483 30 486 33 
rect 483 33 486 36 
rect 483 36 486 39 
rect 483 39 486 42 
rect 483 42 486 45 
rect 483 45 486 48 
rect 483 48 486 51 
rect 483 51 486 54 
rect 483 54 486 57 
rect 483 57 486 60 
rect 483 60 486 63 
rect 483 63 486 66 
rect 483 66 486 69 
rect 483 69 486 72 
rect 483 72 486 75 
rect 483 75 486 78 
rect 483 78 486 81 
rect 483 81 486 84 
rect 483 84 486 87 
rect 483 87 486 90 
rect 483 90 486 93 
rect 483 93 486 96 
rect 483 96 486 99 
rect 483 99 486 102 
rect 483 102 486 105 
rect 483 105 486 108 
rect 483 108 486 111 
rect 483 111 486 114 
rect 483 114 486 117 
rect 483 117 486 120 
rect 483 120 486 123 
rect 483 123 486 126 
rect 483 126 486 129 
rect 483 129 486 132 
rect 483 132 486 135 
rect 483 135 486 138 
rect 483 138 486 141 
rect 483 141 486 144 
rect 483 144 486 147 
rect 483 147 486 150 
rect 483 150 486 153 
rect 483 153 486 156 
rect 483 156 486 159 
rect 483 159 486 162 
rect 483 162 486 165 
rect 483 165 486 168 
rect 483 168 486 171 
rect 483 171 486 174 
rect 483 174 486 177 
rect 483 177 486 180 
rect 483 180 486 183 
rect 483 183 486 186 
rect 483 186 486 189 
rect 483 189 486 192 
rect 483 192 486 195 
rect 483 195 486 198 
rect 483 198 486 201 
rect 483 201 486 204 
rect 483 204 486 207 
rect 483 207 486 210 
rect 483 210 486 213 
rect 483 213 486 216 
rect 483 216 486 219 
rect 483 219 486 222 
rect 483 222 486 225 
rect 483 225 486 228 
rect 483 228 486 231 
rect 483 231 486 234 
rect 483 234 486 237 
rect 483 237 486 240 
rect 483 240 486 243 
rect 483 243 486 246 
rect 483 246 486 249 
rect 483 249 486 252 
rect 483 252 486 255 
rect 483 255 486 258 
rect 483 258 486 261 
rect 483 261 486 264 
rect 483 264 486 267 
rect 483 267 486 270 
rect 483 270 486 273 
rect 483 273 486 276 
rect 483 276 486 279 
rect 483 279 486 282 
rect 483 282 486 285 
rect 483 285 486 288 
rect 483 288 486 291 
rect 483 291 486 294 
rect 483 294 486 297 
rect 483 297 486 300 
rect 483 300 486 303 
rect 483 303 486 306 
rect 483 306 486 309 
rect 483 309 486 312 
rect 483 312 486 315 
rect 483 315 486 318 
rect 483 318 486 321 
rect 483 321 486 324 
rect 483 324 486 327 
rect 483 327 486 330 
rect 483 330 486 333 
rect 483 333 486 336 
rect 483 336 486 339 
rect 483 339 486 342 
rect 483 342 486 345 
rect 483 345 486 348 
rect 483 348 486 351 
rect 483 351 486 354 
rect 483 354 486 357 
rect 483 357 486 360 
rect 483 360 486 363 
rect 483 363 486 366 
rect 483 366 486 369 
rect 483 369 486 372 
rect 483 372 486 375 
rect 483 375 486 378 
rect 483 378 486 381 
rect 483 381 486 384 
rect 483 384 486 387 
rect 483 387 486 390 
rect 483 390 486 393 
rect 483 393 486 396 
rect 483 396 486 399 
rect 483 399 486 402 
rect 483 402 486 405 
rect 483 405 486 408 
rect 483 408 486 411 
rect 483 411 486 414 
rect 483 414 486 417 
rect 483 417 486 420 
rect 483 420 486 423 
rect 483 423 486 426 
rect 483 426 486 429 
rect 483 429 486 432 
rect 483 432 486 435 
rect 483 435 486 438 
rect 483 438 486 441 
rect 483 441 486 444 
rect 483 444 486 447 
rect 483 447 486 450 
rect 483 450 486 453 
rect 483 453 486 456 
rect 483 456 486 459 
rect 483 459 486 462 
rect 483 462 486 465 
rect 483 465 486 468 
rect 483 468 486 471 
rect 483 471 486 474 
rect 483 474 486 477 
rect 483 477 486 480 
rect 483 480 486 483 
rect 483 483 486 486 
rect 483 486 486 489 
rect 483 489 486 492 
rect 483 492 486 495 
rect 483 495 486 498 
rect 483 498 486 501 
rect 483 501 486 504 
rect 483 504 486 507 
rect 483 507 486 510 
rect 486 0 489 3 
rect 486 3 489 6 
rect 486 6 489 9 
rect 486 9 489 12 
rect 486 12 489 15 
rect 486 15 489 18 
rect 486 18 489 21 
rect 486 21 489 24 
rect 486 24 489 27 
rect 486 27 489 30 
rect 486 30 489 33 
rect 486 33 489 36 
rect 486 36 489 39 
rect 486 39 489 42 
rect 486 42 489 45 
rect 486 45 489 48 
rect 486 48 489 51 
rect 486 51 489 54 
rect 486 54 489 57 
rect 486 57 489 60 
rect 486 60 489 63 
rect 486 63 489 66 
rect 486 66 489 69 
rect 486 69 489 72 
rect 486 72 489 75 
rect 486 75 489 78 
rect 486 78 489 81 
rect 486 81 489 84 
rect 486 84 489 87 
rect 486 87 489 90 
rect 486 90 489 93 
rect 486 93 489 96 
rect 486 96 489 99 
rect 486 99 489 102 
rect 486 102 489 105 
rect 486 105 489 108 
rect 486 108 489 111 
rect 486 111 489 114 
rect 486 114 489 117 
rect 486 117 489 120 
rect 486 120 489 123 
rect 486 123 489 126 
rect 486 126 489 129 
rect 486 129 489 132 
rect 486 132 489 135 
rect 486 135 489 138 
rect 486 138 489 141 
rect 486 141 489 144 
rect 486 144 489 147 
rect 486 147 489 150 
rect 486 150 489 153 
rect 486 153 489 156 
rect 486 156 489 159 
rect 486 159 489 162 
rect 486 162 489 165 
rect 486 165 489 168 
rect 486 168 489 171 
rect 486 171 489 174 
rect 486 174 489 177 
rect 486 177 489 180 
rect 486 180 489 183 
rect 486 183 489 186 
rect 486 186 489 189 
rect 486 189 489 192 
rect 486 192 489 195 
rect 486 195 489 198 
rect 486 198 489 201 
rect 486 201 489 204 
rect 486 204 489 207 
rect 486 207 489 210 
rect 486 210 489 213 
rect 486 213 489 216 
rect 486 216 489 219 
rect 486 219 489 222 
rect 486 222 489 225 
rect 486 225 489 228 
rect 486 228 489 231 
rect 486 231 489 234 
rect 486 234 489 237 
rect 486 237 489 240 
rect 486 240 489 243 
rect 486 243 489 246 
rect 486 246 489 249 
rect 486 249 489 252 
rect 486 252 489 255 
rect 486 255 489 258 
rect 486 258 489 261 
rect 486 261 489 264 
rect 486 264 489 267 
rect 486 267 489 270 
rect 486 270 489 273 
rect 486 273 489 276 
rect 486 276 489 279 
rect 486 279 489 282 
rect 486 282 489 285 
rect 486 285 489 288 
rect 486 288 489 291 
rect 486 291 489 294 
rect 486 294 489 297 
rect 486 297 489 300 
rect 486 300 489 303 
rect 486 303 489 306 
rect 486 306 489 309 
rect 486 309 489 312 
rect 486 312 489 315 
rect 486 315 489 318 
rect 486 318 489 321 
rect 486 321 489 324 
rect 486 324 489 327 
rect 486 327 489 330 
rect 486 330 489 333 
rect 486 333 489 336 
rect 486 336 489 339 
rect 486 339 489 342 
rect 486 342 489 345 
rect 486 345 489 348 
rect 486 348 489 351 
rect 486 351 489 354 
rect 486 354 489 357 
rect 486 357 489 360 
rect 486 360 489 363 
rect 486 363 489 366 
rect 486 366 489 369 
rect 486 369 489 372 
rect 486 372 489 375 
rect 486 375 489 378 
rect 486 378 489 381 
rect 486 381 489 384 
rect 486 384 489 387 
rect 486 387 489 390 
rect 486 390 489 393 
rect 486 393 489 396 
rect 486 396 489 399 
rect 486 399 489 402 
rect 486 402 489 405 
rect 486 405 489 408 
rect 486 408 489 411 
rect 486 411 489 414 
rect 486 414 489 417 
rect 486 417 489 420 
rect 486 420 489 423 
rect 486 423 489 426 
rect 486 426 489 429 
rect 486 429 489 432 
rect 486 432 489 435 
rect 486 435 489 438 
rect 486 438 489 441 
rect 486 441 489 444 
rect 486 444 489 447 
rect 486 447 489 450 
rect 486 450 489 453 
rect 486 453 489 456 
rect 486 456 489 459 
rect 486 459 489 462 
rect 486 462 489 465 
rect 486 465 489 468 
rect 486 468 489 471 
rect 486 471 489 474 
rect 486 474 489 477 
rect 486 477 489 480 
rect 486 480 489 483 
rect 486 483 489 486 
rect 486 486 489 489 
rect 486 489 489 492 
rect 486 492 489 495 
rect 486 495 489 498 
rect 486 498 489 501 
rect 486 501 489 504 
rect 486 504 489 507 
rect 486 507 489 510 
rect 489 0 492 3 
rect 489 3 492 6 
rect 489 6 492 9 
rect 489 9 492 12 
rect 489 12 492 15 
rect 489 15 492 18 
rect 489 18 492 21 
rect 489 21 492 24 
rect 489 24 492 27 
rect 489 27 492 30 
rect 489 30 492 33 
rect 489 33 492 36 
rect 489 36 492 39 
rect 489 39 492 42 
rect 489 42 492 45 
rect 489 45 492 48 
rect 489 48 492 51 
rect 489 51 492 54 
rect 489 54 492 57 
rect 489 57 492 60 
rect 489 60 492 63 
rect 489 63 492 66 
rect 489 66 492 69 
rect 489 69 492 72 
rect 489 72 492 75 
rect 489 75 492 78 
rect 489 78 492 81 
rect 489 81 492 84 
rect 489 84 492 87 
rect 489 87 492 90 
rect 489 90 492 93 
rect 489 93 492 96 
rect 489 96 492 99 
rect 489 99 492 102 
rect 489 102 492 105 
rect 489 105 492 108 
rect 489 108 492 111 
rect 489 111 492 114 
rect 489 114 492 117 
rect 489 117 492 120 
rect 489 120 492 123 
rect 489 123 492 126 
rect 489 126 492 129 
rect 489 129 492 132 
rect 489 132 492 135 
rect 489 135 492 138 
rect 489 138 492 141 
rect 489 141 492 144 
rect 489 144 492 147 
rect 489 147 492 150 
rect 489 150 492 153 
rect 489 153 492 156 
rect 489 156 492 159 
rect 489 159 492 162 
rect 489 162 492 165 
rect 489 165 492 168 
rect 489 168 492 171 
rect 489 171 492 174 
rect 489 174 492 177 
rect 489 177 492 180 
rect 489 180 492 183 
rect 489 183 492 186 
rect 489 186 492 189 
rect 489 189 492 192 
rect 489 192 492 195 
rect 489 195 492 198 
rect 489 198 492 201 
rect 489 201 492 204 
rect 489 204 492 207 
rect 489 207 492 210 
rect 489 210 492 213 
rect 489 213 492 216 
rect 489 216 492 219 
rect 489 219 492 222 
rect 489 222 492 225 
rect 489 225 492 228 
rect 489 228 492 231 
rect 489 231 492 234 
rect 489 234 492 237 
rect 489 237 492 240 
rect 489 240 492 243 
rect 489 243 492 246 
rect 489 246 492 249 
rect 489 249 492 252 
rect 489 252 492 255 
rect 489 255 492 258 
rect 489 258 492 261 
rect 489 261 492 264 
rect 489 264 492 267 
rect 489 267 492 270 
rect 489 270 492 273 
rect 489 273 492 276 
rect 489 276 492 279 
rect 489 279 492 282 
rect 489 282 492 285 
rect 489 285 492 288 
rect 489 288 492 291 
rect 489 291 492 294 
rect 489 294 492 297 
rect 489 297 492 300 
rect 489 300 492 303 
rect 489 303 492 306 
rect 489 306 492 309 
rect 489 309 492 312 
rect 489 312 492 315 
rect 489 315 492 318 
rect 489 318 492 321 
rect 489 321 492 324 
rect 489 324 492 327 
rect 489 327 492 330 
rect 489 330 492 333 
rect 489 333 492 336 
rect 489 336 492 339 
rect 489 339 492 342 
rect 489 342 492 345 
rect 489 345 492 348 
rect 489 348 492 351 
rect 489 351 492 354 
rect 489 354 492 357 
rect 489 357 492 360 
rect 489 360 492 363 
rect 489 363 492 366 
rect 489 366 492 369 
rect 489 369 492 372 
rect 489 372 492 375 
rect 489 375 492 378 
rect 489 378 492 381 
rect 489 381 492 384 
rect 489 384 492 387 
rect 489 387 492 390 
rect 489 390 492 393 
rect 489 393 492 396 
rect 489 396 492 399 
rect 489 399 492 402 
rect 489 402 492 405 
rect 489 405 492 408 
rect 489 408 492 411 
rect 489 411 492 414 
rect 489 414 492 417 
rect 489 417 492 420 
rect 489 420 492 423 
rect 489 423 492 426 
rect 489 426 492 429 
rect 489 429 492 432 
rect 489 432 492 435 
rect 489 435 492 438 
rect 489 438 492 441 
rect 489 441 492 444 
rect 489 444 492 447 
rect 489 447 492 450 
rect 489 450 492 453 
rect 489 453 492 456 
rect 489 456 492 459 
rect 489 459 492 462 
rect 489 462 492 465 
rect 489 465 492 468 
rect 489 468 492 471 
rect 489 471 492 474 
rect 489 474 492 477 
rect 489 477 492 480 
rect 489 480 492 483 
rect 489 483 492 486 
rect 489 486 492 489 
rect 489 489 492 492 
rect 489 492 492 495 
rect 489 495 492 498 
rect 489 498 492 501 
rect 489 501 492 504 
rect 489 504 492 507 
rect 489 507 492 510 
rect 492 0 495 3 
rect 492 3 495 6 
rect 492 6 495 9 
rect 492 9 495 12 
rect 492 12 495 15 
rect 492 15 495 18 
rect 492 18 495 21 
rect 492 21 495 24 
rect 492 24 495 27 
rect 492 27 495 30 
rect 492 30 495 33 
rect 492 33 495 36 
rect 492 36 495 39 
rect 492 39 495 42 
rect 492 42 495 45 
rect 492 45 495 48 
rect 492 48 495 51 
rect 492 51 495 54 
rect 492 54 495 57 
rect 492 57 495 60 
rect 492 60 495 63 
rect 492 63 495 66 
rect 492 66 495 69 
rect 492 69 495 72 
rect 492 72 495 75 
rect 492 75 495 78 
rect 492 78 495 81 
rect 492 81 495 84 
rect 492 84 495 87 
rect 492 87 495 90 
rect 492 90 495 93 
rect 492 93 495 96 
rect 492 96 495 99 
rect 492 99 495 102 
rect 492 102 495 105 
rect 492 105 495 108 
rect 492 108 495 111 
rect 492 111 495 114 
rect 492 114 495 117 
rect 492 117 495 120 
rect 492 120 495 123 
rect 492 123 495 126 
rect 492 126 495 129 
rect 492 129 495 132 
rect 492 132 495 135 
rect 492 135 495 138 
rect 492 138 495 141 
rect 492 141 495 144 
rect 492 144 495 147 
rect 492 147 495 150 
rect 492 150 495 153 
rect 492 153 495 156 
rect 492 156 495 159 
rect 492 159 495 162 
rect 492 162 495 165 
rect 492 165 495 168 
rect 492 168 495 171 
rect 492 171 495 174 
rect 492 174 495 177 
rect 492 177 495 180 
rect 492 180 495 183 
rect 492 183 495 186 
rect 492 186 495 189 
rect 492 189 495 192 
rect 492 192 495 195 
rect 492 195 495 198 
rect 492 198 495 201 
rect 492 201 495 204 
rect 492 204 495 207 
rect 492 207 495 210 
rect 492 210 495 213 
rect 492 213 495 216 
rect 492 216 495 219 
rect 492 219 495 222 
rect 492 222 495 225 
rect 492 225 495 228 
rect 492 228 495 231 
rect 492 231 495 234 
rect 492 234 495 237 
rect 492 237 495 240 
rect 492 240 495 243 
rect 492 243 495 246 
rect 492 246 495 249 
rect 492 249 495 252 
rect 492 252 495 255 
rect 492 255 495 258 
rect 492 258 495 261 
rect 492 261 495 264 
rect 492 264 495 267 
rect 492 267 495 270 
rect 492 270 495 273 
rect 492 273 495 276 
rect 492 276 495 279 
rect 492 279 495 282 
rect 492 282 495 285 
rect 492 285 495 288 
rect 492 288 495 291 
rect 492 291 495 294 
rect 492 294 495 297 
rect 492 297 495 300 
rect 492 300 495 303 
rect 492 303 495 306 
rect 492 306 495 309 
rect 492 309 495 312 
rect 492 312 495 315 
rect 492 315 495 318 
rect 492 318 495 321 
rect 492 321 495 324 
rect 492 324 495 327 
rect 492 327 495 330 
rect 492 330 495 333 
rect 492 333 495 336 
rect 492 336 495 339 
rect 492 339 495 342 
rect 492 342 495 345 
rect 492 345 495 348 
rect 492 348 495 351 
rect 492 351 495 354 
rect 492 354 495 357 
rect 492 357 495 360 
rect 492 360 495 363 
rect 492 363 495 366 
rect 492 366 495 369 
rect 492 369 495 372 
rect 492 372 495 375 
rect 492 375 495 378 
rect 492 378 495 381 
rect 492 381 495 384 
rect 492 384 495 387 
rect 492 387 495 390 
rect 492 390 495 393 
rect 492 393 495 396 
rect 492 396 495 399 
rect 492 399 495 402 
rect 492 402 495 405 
rect 492 405 495 408 
rect 492 408 495 411 
rect 492 411 495 414 
rect 492 414 495 417 
rect 492 417 495 420 
rect 492 420 495 423 
rect 492 423 495 426 
rect 492 426 495 429 
rect 492 429 495 432 
rect 492 432 495 435 
rect 492 435 495 438 
rect 492 438 495 441 
rect 492 441 495 444 
rect 492 444 495 447 
rect 492 447 495 450 
rect 492 450 495 453 
rect 492 453 495 456 
rect 492 456 495 459 
rect 492 459 495 462 
rect 492 462 495 465 
rect 492 465 495 468 
rect 492 468 495 471 
rect 492 471 495 474 
rect 492 474 495 477 
rect 492 477 495 480 
rect 492 480 495 483 
rect 492 483 495 486 
rect 492 486 495 489 
rect 492 489 495 492 
rect 492 492 495 495 
rect 492 495 495 498 
rect 492 498 495 501 
rect 492 501 495 504 
rect 492 504 495 507 
rect 492 507 495 510 
rect 495 0 498 3 
rect 495 3 498 6 
rect 495 6 498 9 
rect 495 9 498 12 
rect 495 12 498 15 
rect 495 15 498 18 
rect 495 18 498 21 
rect 495 21 498 24 
rect 495 24 498 27 
rect 495 27 498 30 
rect 495 30 498 33 
rect 495 33 498 36 
rect 495 36 498 39 
rect 495 39 498 42 
rect 495 42 498 45 
rect 495 45 498 48 
rect 495 48 498 51 
rect 495 51 498 54 
rect 495 54 498 57 
rect 495 57 498 60 
rect 495 60 498 63 
rect 495 63 498 66 
rect 495 66 498 69 
rect 495 69 498 72 
rect 495 72 498 75 
rect 495 75 498 78 
rect 495 78 498 81 
rect 495 81 498 84 
rect 495 84 498 87 
rect 495 87 498 90 
rect 495 90 498 93 
rect 495 93 498 96 
rect 495 96 498 99 
rect 495 99 498 102 
rect 495 102 498 105 
rect 495 105 498 108 
rect 495 108 498 111 
rect 495 111 498 114 
rect 495 114 498 117 
rect 495 117 498 120 
rect 495 120 498 123 
rect 495 123 498 126 
rect 495 126 498 129 
rect 495 129 498 132 
rect 495 132 498 135 
rect 495 135 498 138 
rect 495 138 498 141 
rect 495 141 498 144 
rect 495 144 498 147 
rect 495 147 498 150 
rect 495 150 498 153 
rect 495 153 498 156 
rect 495 156 498 159 
rect 495 159 498 162 
rect 495 162 498 165 
rect 495 165 498 168 
rect 495 168 498 171 
rect 495 171 498 174 
rect 495 174 498 177 
rect 495 177 498 180 
rect 495 180 498 183 
rect 495 183 498 186 
rect 495 186 498 189 
rect 495 189 498 192 
rect 495 192 498 195 
rect 495 195 498 198 
rect 495 198 498 201 
rect 495 201 498 204 
rect 495 204 498 207 
rect 495 207 498 210 
rect 495 210 498 213 
rect 495 213 498 216 
rect 495 216 498 219 
rect 495 219 498 222 
rect 495 222 498 225 
rect 495 225 498 228 
rect 495 228 498 231 
rect 495 231 498 234 
rect 495 234 498 237 
rect 495 237 498 240 
rect 495 240 498 243 
rect 495 243 498 246 
rect 495 246 498 249 
rect 495 249 498 252 
rect 495 252 498 255 
rect 495 255 498 258 
rect 495 258 498 261 
rect 495 261 498 264 
rect 495 264 498 267 
rect 495 267 498 270 
rect 495 270 498 273 
rect 495 273 498 276 
rect 495 276 498 279 
rect 495 279 498 282 
rect 495 282 498 285 
rect 495 285 498 288 
rect 495 288 498 291 
rect 495 291 498 294 
rect 495 294 498 297 
rect 495 297 498 300 
rect 495 300 498 303 
rect 495 303 498 306 
rect 495 306 498 309 
rect 495 309 498 312 
rect 495 312 498 315 
rect 495 315 498 318 
rect 495 318 498 321 
rect 495 321 498 324 
rect 495 324 498 327 
rect 495 327 498 330 
rect 495 330 498 333 
rect 495 333 498 336 
rect 495 336 498 339 
rect 495 339 498 342 
rect 495 342 498 345 
rect 495 345 498 348 
rect 495 348 498 351 
rect 495 351 498 354 
rect 495 354 498 357 
rect 495 357 498 360 
rect 495 360 498 363 
rect 495 363 498 366 
rect 495 366 498 369 
rect 495 369 498 372 
rect 495 372 498 375 
rect 495 375 498 378 
rect 495 378 498 381 
rect 495 381 498 384 
rect 495 384 498 387 
rect 495 387 498 390 
rect 495 390 498 393 
rect 495 393 498 396 
rect 495 396 498 399 
rect 495 399 498 402 
rect 495 402 498 405 
rect 495 405 498 408 
rect 495 408 498 411 
rect 495 411 498 414 
rect 495 414 498 417 
rect 495 417 498 420 
rect 495 420 498 423 
rect 495 423 498 426 
rect 495 426 498 429 
rect 495 429 498 432 
rect 495 432 498 435 
rect 495 435 498 438 
rect 495 438 498 441 
rect 495 441 498 444 
rect 495 444 498 447 
rect 495 447 498 450 
rect 495 450 498 453 
rect 495 453 498 456 
rect 495 456 498 459 
rect 495 459 498 462 
rect 495 462 498 465 
rect 495 465 498 468 
rect 495 468 498 471 
rect 495 471 498 474 
rect 495 474 498 477 
rect 495 477 498 480 
rect 495 480 498 483 
rect 495 483 498 486 
rect 495 486 498 489 
rect 495 489 498 492 
rect 495 492 498 495 
rect 495 495 498 498 
rect 495 498 498 501 
rect 495 501 498 504 
rect 495 504 498 507 
rect 495 507 498 510 
rect 498 0 501 3 
rect 498 3 501 6 
rect 498 6 501 9 
rect 498 9 501 12 
rect 498 12 501 15 
rect 498 15 501 18 
rect 498 18 501 21 
rect 498 21 501 24 
rect 498 24 501 27 
rect 498 27 501 30 
rect 498 30 501 33 
rect 498 33 501 36 
rect 498 36 501 39 
rect 498 39 501 42 
rect 498 42 501 45 
rect 498 45 501 48 
rect 498 48 501 51 
rect 498 51 501 54 
rect 498 54 501 57 
rect 498 57 501 60 
rect 498 60 501 63 
rect 498 63 501 66 
rect 498 66 501 69 
rect 498 69 501 72 
rect 498 72 501 75 
rect 498 75 501 78 
rect 498 78 501 81 
rect 498 81 501 84 
rect 498 84 501 87 
rect 498 87 501 90 
rect 498 90 501 93 
rect 498 93 501 96 
rect 498 96 501 99 
rect 498 99 501 102 
rect 498 102 501 105 
rect 498 105 501 108 
rect 498 108 501 111 
rect 498 111 501 114 
rect 498 114 501 117 
rect 498 117 501 120 
rect 498 120 501 123 
rect 498 123 501 126 
rect 498 126 501 129 
rect 498 129 501 132 
rect 498 132 501 135 
rect 498 135 501 138 
rect 498 138 501 141 
rect 498 141 501 144 
rect 498 144 501 147 
rect 498 147 501 150 
rect 498 150 501 153 
rect 498 153 501 156 
rect 498 156 501 159 
rect 498 159 501 162 
rect 498 162 501 165 
rect 498 165 501 168 
rect 498 168 501 171 
rect 498 171 501 174 
rect 498 174 501 177 
rect 498 177 501 180 
rect 498 180 501 183 
rect 498 183 501 186 
rect 498 186 501 189 
rect 498 189 501 192 
rect 498 192 501 195 
rect 498 195 501 198 
rect 498 198 501 201 
rect 498 201 501 204 
rect 498 204 501 207 
rect 498 207 501 210 
rect 498 210 501 213 
rect 498 213 501 216 
rect 498 216 501 219 
rect 498 219 501 222 
rect 498 222 501 225 
rect 498 225 501 228 
rect 498 228 501 231 
rect 498 231 501 234 
rect 498 234 501 237 
rect 498 237 501 240 
rect 498 240 501 243 
rect 498 243 501 246 
rect 498 246 501 249 
rect 498 249 501 252 
rect 498 252 501 255 
rect 498 255 501 258 
rect 498 258 501 261 
rect 498 261 501 264 
rect 498 264 501 267 
rect 498 267 501 270 
rect 498 270 501 273 
rect 498 273 501 276 
rect 498 276 501 279 
rect 498 279 501 282 
rect 498 282 501 285 
rect 498 285 501 288 
rect 498 288 501 291 
rect 498 291 501 294 
rect 498 294 501 297 
rect 498 297 501 300 
rect 498 300 501 303 
rect 498 303 501 306 
rect 498 306 501 309 
rect 498 309 501 312 
rect 498 312 501 315 
rect 498 315 501 318 
rect 498 318 501 321 
rect 498 321 501 324 
rect 498 324 501 327 
rect 498 327 501 330 
rect 498 330 501 333 
rect 498 333 501 336 
rect 498 336 501 339 
rect 498 339 501 342 
rect 498 342 501 345 
rect 498 345 501 348 
rect 498 348 501 351 
rect 498 351 501 354 
rect 498 354 501 357 
rect 498 357 501 360 
rect 498 360 501 363 
rect 498 363 501 366 
rect 498 366 501 369 
rect 498 369 501 372 
rect 498 372 501 375 
rect 498 375 501 378 
rect 498 378 501 381 
rect 498 381 501 384 
rect 498 384 501 387 
rect 498 387 501 390 
rect 498 390 501 393 
rect 498 393 501 396 
rect 498 396 501 399 
rect 498 399 501 402 
rect 498 402 501 405 
rect 498 405 501 408 
rect 498 408 501 411 
rect 498 411 501 414 
rect 498 414 501 417 
rect 498 417 501 420 
rect 498 420 501 423 
rect 498 423 501 426 
rect 498 426 501 429 
rect 498 429 501 432 
rect 498 432 501 435 
rect 498 435 501 438 
rect 498 438 501 441 
rect 498 441 501 444 
rect 498 444 501 447 
rect 498 447 501 450 
rect 498 450 501 453 
rect 498 453 501 456 
rect 498 456 501 459 
rect 498 459 501 462 
rect 498 462 501 465 
rect 498 465 501 468 
rect 498 468 501 471 
rect 498 471 501 474 
rect 498 474 501 477 
rect 498 477 501 480 
rect 498 480 501 483 
rect 498 483 501 486 
rect 498 486 501 489 
rect 498 489 501 492 
rect 498 492 501 495 
rect 498 495 501 498 
rect 498 498 501 501 
rect 498 501 501 504 
rect 498 504 501 507 
rect 498 507 501 510 
rect 501 0 504 3 
rect 501 3 504 6 
rect 501 6 504 9 
rect 501 9 504 12 
rect 501 12 504 15 
rect 501 15 504 18 
rect 501 18 504 21 
rect 501 21 504 24 
rect 501 24 504 27 
rect 501 27 504 30 
rect 501 30 504 33 
rect 501 33 504 36 
rect 501 36 504 39 
rect 501 39 504 42 
rect 501 42 504 45 
rect 501 45 504 48 
rect 501 48 504 51 
rect 501 51 504 54 
rect 501 54 504 57 
rect 501 57 504 60 
rect 501 60 504 63 
rect 501 63 504 66 
rect 501 66 504 69 
rect 501 69 504 72 
rect 501 72 504 75 
rect 501 75 504 78 
rect 501 78 504 81 
rect 501 81 504 84 
rect 501 84 504 87 
rect 501 87 504 90 
rect 501 90 504 93 
rect 501 93 504 96 
rect 501 96 504 99 
rect 501 99 504 102 
rect 501 102 504 105 
rect 501 105 504 108 
rect 501 108 504 111 
rect 501 111 504 114 
rect 501 114 504 117 
rect 501 117 504 120 
rect 501 120 504 123 
rect 501 123 504 126 
rect 501 126 504 129 
rect 501 129 504 132 
rect 501 132 504 135 
rect 501 135 504 138 
rect 501 138 504 141 
rect 501 141 504 144 
rect 501 144 504 147 
rect 501 147 504 150 
rect 501 150 504 153 
rect 501 153 504 156 
rect 501 156 504 159 
rect 501 159 504 162 
rect 501 162 504 165 
rect 501 165 504 168 
rect 501 168 504 171 
rect 501 171 504 174 
rect 501 174 504 177 
rect 501 177 504 180 
rect 501 180 504 183 
rect 501 183 504 186 
rect 501 186 504 189 
rect 501 189 504 192 
rect 501 192 504 195 
rect 501 195 504 198 
rect 501 198 504 201 
rect 501 201 504 204 
rect 501 204 504 207 
rect 501 207 504 210 
rect 501 210 504 213 
rect 501 213 504 216 
rect 501 216 504 219 
rect 501 219 504 222 
rect 501 222 504 225 
rect 501 225 504 228 
rect 501 228 504 231 
rect 501 231 504 234 
rect 501 234 504 237 
rect 501 237 504 240 
rect 501 240 504 243 
rect 501 243 504 246 
rect 501 246 504 249 
rect 501 249 504 252 
rect 501 252 504 255 
rect 501 255 504 258 
rect 501 258 504 261 
rect 501 261 504 264 
rect 501 264 504 267 
rect 501 267 504 270 
rect 501 270 504 273 
rect 501 273 504 276 
rect 501 276 504 279 
rect 501 279 504 282 
rect 501 282 504 285 
rect 501 285 504 288 
rect 501 288 504 291 
rect 501 291 504 294 
rect 501 294 504 297 
rect 501 297 504 300 
rect 501 300 504 303 
rect 501 303 504 306 
rect 501 306 504 309 
rect 501 309 504 312 
rect 501 312 504 315 
rect 501 315 504 318 
rect 501 318 504 321 
rect 501 321 504 324 
rect 501 324 504 327 
rect 501 327 504 330 
rect 501 330 504 333 
rect 501 333 504 336 
rect 501 336 504 339 
rect 501 339 504 342 
rect 501 342 504 345 
rect 501 345 504 348 
rect 501 348 504 351 
rect 501 351 504 354 
rect 501 354 504 357 
rect 501 357 504 360 
rect 501 360 504 363 
rect 501 363 504 366 
rect 501 366 504 369 
rect 501 369 504 372 
rect 501 372 504 375 
rect 501 375 504 378 
rect 501 378 504 381 
rect 501 381 504 384 
rect 501 384 504 387 
rect 501 387 504 390 
rect 501 390 504 393 
rect 501 393 504 396 
rect 501 396 504 399 
rect 501 399 504 402 
rect 501 402 504 405 
rect 501 405 504 408 
rect 501 408 504 411 
rect 501 411 504 414 
rect 501 414 504 417 
rect 501 417 504 420 
rect 501 420 504 423 
rect 501 423 504 426 
rect 501 426 504 429 
rect 501 429 504 432 
rect 501 432 504 435 
rect 501 435 504 438 
rect 501 438 504 441 
rect 501 441 504 444 
rect 501 444 504 447 
rect 501 447 504 450 
rect 501 450 504 453 
rect 501 453 504 456 
rect 501 456 504 459 
rect 501 459 504 462 
rect 501 462 504 465 
rect 501 465 504 468 
rect 501 468 504 471 
rect 501 471 504 474 
rect 501 474 504 477 
rect 501 477 504 480 
rect 501 480 504 483 
rect 501 483 504 486 
rect 501 486 504 489 
rect 501 489 504 492 
rect 501 492 504 495 
rect 501 495 504 498 
rect 501 498 504 501 
rect 501 501 504 504 
rect 501 504 504 507 
rect 501 507 504 510 
rect 504 0 507 3 
rect 504 3 507 6 
rect 504 6 507 9 
rect 504 9 507 12 
rect 504 12 507 15 
rect 504 15 507 18 
rect 504 18 507 21 
rect 504 21 507 24 
rect 504 24 507 27 
rect 504 27 507 30 
rect 504 30 507 33 
rect 504 33 507 36 
rect 504 36 507 39 
rect 504 39 507 42 
rect 504 42 507 45 
rect 504 45 507 48 
rect 504 48 507 51 
rect 504 51 507 54 
rect 504 54 507 57 
rect 504 57 507 60 
rect 504 60 507 63 
rect 504 63 507 66 
rect 504 66 507 69 
rect 504 69 507 72 
rect 504 72 507 75 
rect 504 75 507 78 
rect 504 78 507 81 
rect 504 81 507 84 
rect 504 84 507 87 
rect 504 87 507 90 
rect 504 90 507 93 
rect 504 93 507 96 
rect 504 96 507 99 
rect 504 99 507 102 
rect 504 102 507 105 
rect 504 105 507 108 
rect 504 108 507 111 
rect 504 111 507 114 
rect 504 114 507 117 
rect 504 117 507 120 
rect 504 120 507 123 
rect 504 123 507 126 
rect 504 126 507 129 
rect 504 129 507 132 
rect 504 132 507 135 
rect 504 135 507 138 
rect 504 138 507 141 
rect 504 141 507 144 
rect 504 144 507 147 
rect 504 147 507 150 
rect 504 150 507 153 
rect 504 153 507 156 
rect 504 156 507 159 
rect 504 159 507 162 
rect 504 162 507 165 
rect 504 165 507 168 
rect 504 168 507 171 
rect 504 171 507 174 
rect 504 174 507 177 
rect 504 177 507 180 
rect 504 180 507 183 
rect 504 183 507 186 
rect 504 186 507 189 
rect 504 189 507 192 
rect 504 192 507 195 
rect 504 195 507 198 
rect 504 198 507 201 
rect 504 201 507 204 
rect 504 204 507 207 
rect 504 207 507 210 
rect 504 210 507 213 
rect 504 213 507 216 
rect 504 216 507 219 
rect 504 219 507 222 
rect 504 222 507 225 
rect 504 225 507 228 
rect 504 228 507 231 
rect 504 231 507 234 
rect 504 234 507 237 
rect 504 237 507 240 
rect 504 240 507 243 
rect 504 243 507 246 
rect 504 246 507 249 
rect 504 249 507 252 
rect 504 252 507 255 
rect 504 255 507 258 
rect 504 258 507 261 
rect 504 261 507 264 
rect 504 264 507 267 
rect 504 267 507 270 
rect 504 270 507 273 
rect 504 273 507 276 
rect 504 276 507 279 
rect 504 279 507 282 
rect 504 282 507 285 
rect 504 285 507 288 
rect 504 288 507 291 
rect 504 291 507 294 
rect 504 294 507 297 
rect 504 297 507 300 
rect 504 300 507 303 
rect 504 303 507 306 
rect 504 306 507 309 
rect 504 309 507 312 
rect 504 312 507 315 
rect 504 315 507 318 
rect 504 318 507 321 
rect 504 321 507 324 
rect 504 324 507 327 
rect 504 327 507 330 
rect 504 330 507 333 
rect 504 333 507 336 
rect 504 336 507 339 
rect 504 339 507 342 
rect 504 342 507 345 
rect 504 345 507 348 
rect 504 348 507 351 
rect 504 351 507 354 
rect 504 354 507 357 
rect 504 357 507 360 
rect 504 360 507 363 
rect 504 363 507 366 
rect 504 366 507 369 
rect 504 369 507 372 
rect 504 372 507 375 
rect 504 375 507 378 
rect 504 378 507 381 
rect 504 381 507 384 
rect 504 384 507 387 
rect 504 387 507 390 
rect 504 390 507 393 
rect 504 393 507 396 
rect 504 396 507 399 
rect 504 399 507 402 
rect 504 402 507 405 
rect 504 405 507 408 
rect 504 408 507 411 
rect 504 411 507 414 
rect 504 414 507 417 
rect 504 417 507 420 
rect 504 420 507 423 
rect 504 423 507 426 
rect 504 426 507 429 
rect 504 429 507 432 
rect 504 432 507 435 
rect 504 435 507 438 
rect 504 438 507 441 
rect 504 441 507 444 
rect 504 444 507 447 
rect 504 447 507 450 
rect 504 450 507 453 
rect 504 453 507 456 
rect 504 456 507 459 
rect 504 459 507 462 
rect 504 462 507 465 
rect 504 465 507 468 
rect 504 468 507 471 
rect 504 471 507 474 
rect 504 474 507 477 
rect 504 477 507 480 
rect 504 480 507 483 
rect 504 483 507 486 
rect 504 486 507 489 
rect 504 489 507 492 
rect 504 492 507 495 
rect 504 495 507 498 
rect 504 498 507 501 
rect 504 501 507 504 
rect 504 504 507 507 
rect 504 507 507 510 
rect 507 0 510 3 
rect 507 3 510 6 
rect 507 6 510 9 
rect 507 9 510 12 
rect 507 12 510 15 
rect 507 15 510 18 
rect 507 18 510 21 
rect 507 21 510 24 
rect 507 24 510 27 
rect 507 27 510 30 
rect 507 30 510 33 
rect 507 33 510 36 
rect 507 36 510 39 
rect 507 39 510 42 
rect 507 42 510 45 
rect 507 45 510 48 
rect 507 48 510 51 
rect 507 51 510 54 
rect 507 54 510 57 
rect 507 57 510 60 
rect 507 60 510 63 
rect 507 63 510 66 
rect 507 66 510 69 
rect 507 69 510 72 
rect 507 72 510 75 
rect 507 75 510 78 
rect 507 78 510 81 
rect 507 81 510 84 
rect 507 84 510 87 
rect 507 87 510 90 
rect 507 90 510 93 
rect 507 93 510 96 
rect 507 96 510 99 
rect 507 99 510 102 
rect 507 102 510 105 
rect 507 105 510 108 
rect 507 108 510 111 
rect 507 111 510 114 
rect 507 114 510 117 
rect 507 117 510 120 
rect 507 120 510 123 
rect 507 123 510 126 
rect 507 126 510 129 
rect 507 129 510 132 
rect 507 132 510 135 
rect 507 135 510 138 
rect 507 138 510 141 
rect 507 141 510 144 
rect 507 144 510 147 
rect 507 147 510 150 
rect 507 150 510 153 
rect 507 153 510 156 
rect 507 156 510 159 
rect 507 159 510 162 
rect 507 162 510 165 
rect 507 165 510 168 
rect 507 168 510 171 
rect 507 171 510 174 
rect 507 174 510 177 
rect 507 177 510 180 
rect 507 180 510 183 
rect 507 183 510 186 
rect 507 186 510 189 
rect 507 189 510 192 
rect 507 192 510 195 
rect 507 195 510 198 
rect 507 198 510 201 
rect 507 201 510 204 
rect 507 204 510 207 
rect 507 207 510 210 
rect 507 210 510 213 
rect 507 213 510 216 
rect 507 216 510 219 
rect 507 219 510 222 
rect 507 222 510 225 
rect 507 225 510 228 
rect 507 228 510 231 
rect 507 231 510 234 
rect 507 234 510 237 
rect 507 237 510 240 
rect 507 240 510 243 
rect 507 243 510 246 
rect 507 246 510 249 
rect 507 249 510 252 
rect 507 252 510 255 
rect 507 255 510 258 
rect 507 258 510 261 
rect 507 261 510 264 
rect 507 264 510 267 
rect 507 267 510 270 
rect 507 270 510 273 
rect 507 273 510 276 
rect 507 276 510 279 
rect 507 279 510 282 
rect 507 282 510 285 
rect 507 285 510 288 
rect 507 288 510 291 
rect 507 291 510 294 
rect 507 294 510 297 
rect 507 297 510 300 
rect 507 300 510 303 
rect 507 303 510 306 
rect 507 306 510 309 
rect 507 309 510 312 
rect 507 312 510 315 
rect 507 315 510 318 
rect 507 318 510 321 
rect 507 321 510 324 
rect 507 324 510 327 
rect 507 327 510 330 
rect 507 330 510 333 
rect 507 333 510 336 
rect 507 336 510 339 
rect 507 339 510 342 
rect 507 342 510 345 
rect 507 345 510 348 
rect 507 348 510 351 
rect 507 351 510 354 
rect 507 354 510 357 
rect 507 357 510 360 
rect 507 360 510 363 
rect 507 363 510 366 
rect 507 366 510 369 
rect 507 369 510 372 
rect 507 372 510 375 
rect 507 375 510 378 
rect 507 378 510 381 
rect 507 381 510 384 
rect 507 384 510 387 
rect 507 387 510 390 
rect 507 390 510 393 
rect 507 393 510 396 
rect 507 396 510 399 
rect 507 399 510 402 
rect 507 402 510 405 
rect 507 405 510 408 
rect 507 408 510 411 
rect 507 411 510 414 
rect 507 414 510 417 
rect 507 417 510 420 
rect 507 420 510 423 
rect 507 423 510 426 
rect 507 426 510 429 
rect 507 429 510 432 
rect 507 432 510 435 
rect 507 435 510 438 
rect 507 438 510 441 
rect 507 441 510 444 
rect 507 444 510 447 
rect 507 447 510 450 
rect 507 450 510 453 
rect 507 453 510 456 
rect 507 456 510 459 
rect 507 459 510 462 
rect 507 462 510 465 
rect 507 465 510 468 
rect 507 468 510 471 
rect 507 471 510 474 
rect 507 474 510 477 
rect 507 477 510 480 
rect 507 480 510 483 
rect 507 483 510 486 
rect 507 486 510 489 
rect 507 489 510 492 
rect 507 492 510 495 
rect 507 495 510 498 
rect 507 498 510 501 
rect 507 501 510 504 
rect 507 504 510 507 
rect 507 507 510 510 
<< metal2 >>
rect 0 0 3 3 
rect 0 3 3 6 
rect 0 6 3 9 
rect 0 9 3 12 
rect 0 12 3 15 
rect 0 15 3 18 
rect 0 18 3 21 
rect 0 21 3 24 
rect 0 24 3 27 
rect 0 27 3 30 
rect 0 30 3 33 
rect 0 33 3 36 
rect 0 36 3 39 
rect 0 39 3 42 
rect 0 42 3 45 
rect 0 45 3 48 
rect 0 48 3 51 
rect 0 51 3 54 
rect 0 54 3 57 
rect 0 57 3 60 
rect 0 60 3 63 
rect 0 63 3 66 
rect 0 66 3 69 
rect 0 69 3 72 
rect 0 72 3 75 
rect 0 75 3 78 
rect 0 78 3 81 
rect 0 81 3 84 
rect 0 84 3 87 
rect 0 87 3 90 
rect 0 90 3 93 
rect 0 93 3 96 
rect 0 96 3 99 
rect 0 99 3 102 
rect 0 102 3 105 
rect 0 105 3 108 
rect 0 108 3 111 
rect 0 111 3 114 
rect 0 114 3 117 
rect 0 117 3 120 
rect 0 120 3 123 
rect 0 123 3 126 
rect 0 126 3 129 
rect 0 129 3 132 
rect 0 132 3 135 
rect 0 135 3 138 
rect 0 138 3 141 
rect 0 141 3 144 
rect 0 144 3 147 
rect 0 147 3 150 
rect 0 150 3 153 
rect 0 153 3 156 
rect 0 156 3 159 
rect 0 159 3 162 
rect 0 162 3 165 
rect 0 165 3 168 
rect 0 168 3 171 
rect 0 171 3 174 
rect 0 174 3 177 
rect 0 177 3 180 
rect 0 180 3 183 
rect 0 183 3 186 
rect 0 186 3 189 
rect 0 189 3 192 
rect 0 192 3 195 
rect 0 195 3 198 
rect 0 198 3 201 
rect 0 201 3 204 
rect 0 204 3 207 
rect 0 207 3 210 
rect 0 210 3 213 
rect 0 213 3 216 
rect 0 216 3 219 
rect 0 219 3 222 
rect 0 222 3 225 
rect 0 225 3 228 
rect 0 228 3 231 
rect 0 231 3 234 
rect 0 234 3 237 
rect 0 237 3 240 
rect 0 240 3 243 
rect 0 243 3 246 
rect 0 246 3 249 
rect 0 249 3 252 
rect 0 252 3 255 
rect 0 255 3 258 
rect 0 258 3 261 
rect 0 261 3 264 
rect 0 264 3 267 
rect 0 267 3 270 
rect 0 270 3 273 
rect 0 273 3 276 
rect 0 276 3 279 
rect 0 279 3 282 
rect 0 282 3 285 
rect 0 285 3 288 
rect 0 288 3 291 
rect 0 291 3 294 
rect 0 294 3 297 
rect 0 297 3 300 
rect 0 300 3 303 
rect 0 303 3 306 
rect 0 306 3 309 
rect 0 309 3 312 
rect 0 312 3 315 
rect 0 315 3 318 
rect 0 318 3 321 
rect 0 321 3 324 
rect 0 324 3 327 
rect 0 327 3 330 
rect 0 330 3 333 
rect 0 333 3 336 
rect 0 336 3 339 
rect 0 339 3 342 
rect 0 342 3 345 
rect 0 345 3 348 
rect 0 348 3 351 
rect 0 351 3 354 
rect 0 354 3 357 
rect 0 357 3 360 
rect 0 360 3 363 
rect 0 363 3 366 
rect 0 366 3 369 
rect 0 369 3 372 
rect 0 372 3 375 
rect 0 375 3 378 
rect 0 378 3 381 
rect 0 381 3 384 
rect 0 384 3 387 
rect 0 387 3 390 
rect 0 390 3 393 
rect 0 393 3 396 
rect 0 396 3 399 
rect 0 399 3 402 
rect 0 402 3 405 
rect 0 405 3 408 
rect 0 408 3 411 
rect 0 411 3 414 
rect 0 414 3 417 
rect 0 417 3 420 
rect 0 420 3 423 
rect 0 423 3 426 
rect 0 426 3 429 
rect 0 429 3 432 
rect 0 432 3 435 
rect 0 435 3 438 
rect 0 438 3 441 
rect 0 441 3 444 
rect 0 444 3 447 
rect 0 447 3 450 
rect 0 450 3 453 
rect 0 453 3 456 
rect 0 456 3 459 
rect 0 459 3 462 
rect 0 462 3 465 
rect 0 465 3 468 
rect 0 468 3 471 
rect 0 471 3 474 
rect 0 474 3 477 
rect 0 477 3 480 
rect 0 480 3 483 
rect 0 483 3 486 
rect 0 486 3 489 
rect 0 489 3 492 
rect 0 492 3 495 
rect 0 495 3 498 
rect 0 498 3 501 
rect 0 501 3 504 
rect 0 504 3 507 
rect 0 507 3 510 
rect 3 0 6 3 
rect 3 3 6 6 
rect 3 6 6 9 
rect 3 9 6 12 
rect 3 12 6 15 
rect 3 15 6 18 
rect 3 18 6 21 
rect 3 21 6 24 
rect 3 24 6 27 
rect 3 27 6 30 
rect 3 30 6 33 
rect 3 33 6 36 
rect 3 36 6 39 
rect 3 39 6 42 
rect 3 42 6 45 
rect 3 45 6 48 
rect 3 48 6 51 
rect 3 51 6 54 
rect 3 54 6 57 
rect 3 57 6 60 
rect 3 60 6 63 
rect 3 63 6 66 
rect 3 66 6 69 
rect 3 69 6 72 
rect 3 72 6 75 
rect 3 75 6 78 
rect 3 78 6 81 
rect 3 81 6 84 
rect 3 84 6 87 
rect 3 87 6 90 
rect 3 90 6 93 
rect 3 93 6 96 
rect 3 96 6 99 
rect 3 99 6 102 
rect 3 102 6 105 
rect 3 105 6 108 
rect 3 108 6 111 
rect 3 111 6 114 
rect 3 114 6 117 
rect 3 117 6 120 
rect 3 120 6 123 
rect 3 123 6 126 
rect 3 126 6 129 
rect 3 129 6 132 
rect 3 132 6 135 
rect 3 135 6 138 
rect 3 138 6 141 
rect 3 141 6 144 
rect 3 144 6 147 
rect 3 147 6 150 
rect 3 150 6 153 
rect 3 153 6 156 
rect 3 156 6 159 
rect 3 159 6 162 
rect 3 162 6 165 
rect 3 165 6 168 
rect 3 168 6 171 
rect 3 171 6 174 
rect 3 174 6 177 
rect 3 177 6 180 
rect 3 180 6 183 
rect 3 183 6 186 
rect 3 186 6 189 
rect 3 189 6 192 
rect 3 192 6 195 
rect 3 195 6 198 
rect 3 198 6 201 
rect 3 201 6 204 
rect 3 204 6 207 
rect 3 207 6 210 
rect 3 210 6 213 
rect 3 213 6 216 
rect 3 216 6 219 
rect 3 219 6 222 
rect 3 222 6 225 
rect 3 225 6 228 
rect 3 228 6 231 
rect 3 231 6 234 
rect 3 234 6 237 
rect 3 237 6 240 
rect 3 240 6 243 
rect 3 243 6 246 
rect 3 246 6 249 
rect 3 249 6 252 
rect 3 252 6 255 
rect 3 255 6 258 
rect 3 258 6 261 
rect 3 261 6 264 
rect 3 264 6 267 
rect 3 267 6 270 
rect 3 270 6 273 
rect 3 273 6 276 
rect 3 276 6 279 
rect 3 279 6 282 
rect 3 282 6 285 
rect 3 285 6 288 
rect 3 288 6 291 
rect 3 291 6 294 
rect 3 294 6 297 
rect 3 297 6 300 
rect 3 300 6 303 
rect 3 303 6 306 
rect 3 306 6 309 
rect 3 309 6 312 
rect 3 312 6 315 
rect 3 315 6 318 
rect 3 318 6 321 
rect 3 321 6 324 
rect 3 324 6 327 
rect 3 327 6 330 
rect 3 330 6 333 
rect 3 333 6 336 
rect 3 336 6 339 
rect 3 339 6 342 
rect 3 342 6 345 
rect 3 345 6 348 
rect 3 348 6 351 
rect 3 351 6 354 
rect 3 354 6 357 
rect 3 357 6 360 
rect 3 360 6 363 
rect 3 363 6 366 
rect 3 366 6 369 
rect 3 369 6 372 
rect 3 372 6 375 
rect 3 375 6 378 
rect 3 378 6 381 
rect 3 381 6 384 
rect 3 384 6 387 
rect 3 387 6 390 
rect 3 390 6 393 
rect 3 393 6 396 
rect 3 396 6 399 
rect 3 399 6 402 
rect 3 402 6 405 
rect 3 405 6 408 
rect 3 408 6 411 
rect 3 411 6 414 
rect 3 414 6 417 
rect 3 417 6 420 
rect 3 420 6 423 
rect 3 423 6 426 
rect 3 426 6 429 
rect 3 429 6 432 
rect 3 432 6 435 
rect 3 435 6 438 
rect 3 438 6 441 
rect 3 441 6 444 
rect 3 444 6 447 
rect 3 447 6 450 
rect 3 450 6 453 
rect 3 453 6 456 
rect 3 456 6 459 
rect 3 459 6 462 
rect 3 462 6 465 
rect 3 465 6 468 
rect 3 468 6 471 
rect 3 471 6 474 
rect 3 474 6 477 
rect 3 477 6 480 
rect 3 480 6 483 
rect 3 483 6 486 
rect 3 486 6 489 
rect 3 489 6 492 
rect 3 492 6 495 
rect 3 495 6 498 
rect 3 498 6 501 
rect 3 501 6 504 
rect 3 504 6 507 
rect 3 507 6 510 
rect 6 0 9 3 
rect 6 3 9 6 
rect 6 6 9 9 
rect 6 9 9 12 
rect 6 12 9 15 
rect 6 15 9 18 
rect 6 18 9 21 
rect 6 21 9 24 
rect 6 24 9 27 
rect 6 27 9 30 
rect 6 30 9 33 
rect 6 33 9 36 
rect 6 36 9 39 
rect 6 39 9 42 
rect 6 42 9 45 
rect 6 45 9 48 
rect 6 48 9 51 
rect 6 51 9 54 
rect 6 54 9 57 
rect 6 57 9 60 
rect 6 60 9 63 
rect 6 63 9 66 
rect 6 66 9 69 
rect 6 69 9 72 
rect 6 72 9 75 
rect 6 75 9 78 
rect 6 78 9 81 
rect 6 81 9 84 
rect 6 84 9 87 
rect 6 87 9 90 
rect 6 90 9 93 
rect 6 93 9 96 
rect 6 96 9 99 
rect 6 99 9 102 
rect 6 102 9 105 
rect 6 105 9 108 
rect 6 108 9 111 
rect 6 111 9 114 
rect 6 114 9 117 
rect 6 117 9 120 
rect 6 120 9 123 
rect 6 123 9 126 
rect 6 126 9 129 
rect 6 129 9 132 
rect 6 132 9 135 
rect 6 135 9 138 
rect 6 138 9 141 
rect 6 141 9 144 
rect 6 144 9 147 
rect 6 147 9 150 
rect 6 150 9 153 
rect 6 153 9 156 
rect 6 156 9 159 
rect 6 159 9 162 
rect 6 162 9 165 
rect 6 165 9 168 
rect 6 168 9 171 
rect 6 171 9 174 
rect 6 174 9 177 
rect 6 177 9 180 
rect 6 180 9 183 
rect 6 183 9 186 
rect 6 186 9 189 
rect 6 189 9 192 
rect 6 192 9 195 
rect 6 195 9 198 
rect 6 198 9 201 
rect 6 201 9 204 
rect 6 204 9 207 
rect 6 207 9 210 
rect 6 210 9 213 
rect 6 213 9 216 
rect 6 216 9 219 
rect 6 219 9 222 
rect 6 222 9 225 
rect 6 225 9 228 
rect 6 228 9 231 
rect 6 231 9 234 
rect 6 234 9 237 
rect 6 237 9 240 
rect 6 240 9 243 
rect 6 243 9 246 
rect 6 246 9 249 
rect 6 249 9 252 
rect 6 252 9 255 
rect 6 255 9 258 
rect 6 258 9 261 
rect 6 261 9 264 
rect 6 264 9 267 
rect 6 267 9 270 
rect 6 270 9 273 
rect 6 273 9 276 
rect 6 276 9 279 
rect 6 279 9 282 
rect 6 282 9 285 
rect 6 285 9 288 
rect 6 288 9 291 
rect 6 291 9 294 
rect 6 294 9 297 
rect 6 297 9 300 
rect 6 300 9 303 
rect 6 303 9 306 
rect 6 306 9 309 
rect 6 309 9 312 
rect 6 312 9 315 
rect 6 315 9 318 
rect 6 318 9 321 
rect 6 321 9 324 
rect 6 324 9 327 
rect 6 327 9 330 
rect 6 330 9 333 
rect 6 333 9 336 
rect 6 336 9 339 
rect 6 339 9 342 
rect 6 342 9 345 
rect 6 345 9 348 
rect 6 348 9 351 
rect 6 351 9 354 
rect 6 354 9 357 
rect 6 357 9 360 
rect 6 360 9 363 
rect 6 363 9 366 
rect 6 366 9 369 
rect 6 369 9 372 
rect 6 372 9 375 
rect 6 375 9 378 
rect 6 378 9 381 
rect 6 381 9 384 
rect 6 384 9 387 
rect 6 387 9 390 
rect 6 390 9 393 
rect 6 393 9 396 
rect 6 396 9 399 
rect 6 399 9 402 
rect 6 402 9 405 
rect 6 405 9 408 
rect 6 408 9 411 
rect 6 411 9 414 
rect 6 414 9 417 
rect 6 417 9 420 
rect 6 420 9 423 
rect 6 423 9 426 
rect 6 426 9 429 
rect 6 429 9 432 
rect 6 432 9 435 
rect 6 435 9 438 
rect 6 438 9 441 
rect 6 441 9 444 
rect 6 444 9 447 
rect 6 447 9 450 
rect 6 450 9 453 
rect 6 453 9 456 
rect 6 456 9 459 
rect 6 459 9 462 
rect 6 462 9 465 
rect 6 465 9 468 
rect 6 468 9 471 
rect 6 471 9 474 
rect 6 474 9 477 
rect 6 477 9 480 
rect 6 480 9 483 
rect 6 483 9 486 
rect 6 486 9 489 
rect 6 489 9 492 
rect 6 492 9 495 
rect 6 495 9 498 
rect 6 498 9 501 
rect 6 501 9 504 
rect 6 504 9 507 
rect 6 507 9 510 
rect 9 0 12 3 
rect 9 3 12 6 
rect 9 6 12 9 
rect 9 9 12 12 
rect 9 12 12 15 
rect 9 15 12 18 
rect 9 18 12 21 
rect 9 21 12 24 
rect 9 24 12 27 
rect 9 27 12 30 
rect 9 30 12 33 
rect 9 33 12 36 
rect 9 36 12 39 
rect 9 39 12 42 
rect 9 42 12 45 
rect 9 45 12 48 
rect 9 48 12 51 
rect 9 51 12 54 
rect 9 54 12 57 
rect 9 57 12 60 
rect 9 60 12 63 
rect 9 63 12 66 
rect 9 66 12 69 
rect 9 69 12 72 
rect 9 72 12 75 
rect 9 75 12 78 
rect 9 78 12 81 
rect 9 81 12 84 
rect 9 84 12 87 
rect 9 87 12 90 
rect 9 90 12 93 
rect 9 93 12 96 
rect 9 96 12 99 
rect 9 99 12 102 
rect 9 102 12 105 
rect 9 105 12 108 
rect 9 108 12 111 
rect 9 111 12 114 
rect 9 114 12 117 
rect 9 117 12 120 
rect 9 120 12 123 
rect 9 123 12 126 
rect 9 126 12 129 
rect 9 129 12 132 
rect 9 132 12 135 
rect 9 135 12 138 
rect 9 138 12 141 
rect 9 141 12 144 
rect 9 144 12 147 
rect 9 147 12 150 
rect 9 150 12 153 
rect 9 153 12 156 
rect 9 156 12 159 
rect 9 159 12 162 
rect 9 162 12 165 
rect 9 165 12 168 
rect 9 168 12 171 
rect 9 171 12 174 
rect 9 174 12 177 
rect 9 177 12 180 
rect 9 180 12 183 
rect 9 183 12 186 
rect 9 186 12 189 
rect 9 189 12 192 
rect 9 192 12 195 
rect 9 195 12 198 
rect 9 198 12 201 
rect 9 201 12 204 
rect 9 204 12 207 
rect 9 207 12 210 
rect 9 210 12 213 
rect 9 213 12 216 
rect 9 216 12 219 
rect 9 219 12 222 
rect 9 222 12 225 
rect 9 225 12 228 
rect 9 228 12 231 
rect 9 231 12 234 
rect 9 234 12 237 
rect 9 237 12 240 
rect 9 240 12 243 
rect 9 243 12 246 
rect 9 246 12 249 
rect 9 249 12 252 
rect 9 252 12 255 
rect 9 255 12 258 
rect 9 258 12 261 
rect 9 261 12 264 
rect 9 264 12 267 
rect 9 267 12 270 
rect 9 270 12 273 
rect 9 273 12 276 
rect 9 276 12 279 
rect 9 279 12 282 
rect 9 282 12 285 
rect 9 285 12 288 
rect 9 288 12 291 
rect 9 291 12 294 
rect 9 294 12 297 
rect 9 297 12 300 
rect 9 300 12 303 
rect 9 303 12 306 
rect 9 306 12 309 
rect 9 309 12 312 
rect 9 312 12 315 
rect 9 315 12 318 
rect 9 318 12 321 
rect 9 321 12 324 
rect 9 324 12 327 
rect 9 327 12 330 
rect 9 330 12 333 
rect 9 333 12 336 
rect 9 336 12 339 
rect 9 339 12 342 
rect 9 342 12 345 
rect 9 345 12 348 
rect 9 348 12 351 
rect 9 351 12 354 
rect 9 354 12 357 
rect 9 357 12 360 
rect 9 360 12 363 
rect 9 363 12 366 
rect 9 366 12 369 
rect 9 369 12 372 
rect 9 372 12 375 
rect 9 375 12 378 
rect 9 378 12 381 
rect 9 381 12 384 
rect 9 384 12 387 
rect 9 387 12 390 
rect 9 390 12 393 
rect 9 393 12 396 
rect 9 396 12 399 
rect 9 399 12 402 
rect 9 402 12 405 
rect 9 405 12 408 
rect 9 408 12 411 
rect 9 411 12 414 
rect 9 414 12 417 
rect 9 417 12 420 
rect 9 420 12 423 
rect 9 423 12 426 
rect 9 426 12 429 
rect 9 429 12 432 
rect 9 432 12 435 
rect 9 435 12 438 
rect 9 438 12 441 
rect 9 441 12 444 
rect 9 444 12 447 
rect 9 447 12 450 
rect 9 450 12 453 
rect 9 453 12 456 
rect 9 456 12 459 
rect 9 459 12 462 
rect 9 462 12 465 
rect 9 465 12 468 
rect 9 468 12 471 
rect 9 471 12 474 
rect 9 474 12 477 
rect 9 477 12 480 
rect 9 480 12 483 
rect 9 483 12 486 
rect 9 486 12 489 
rect 9 489 12 492 
rect 9 492 12 495 
rect 9 495 12 498 
rect 9 498 12 501 
rect 9 501 12 504 
rect 9 504 12 507 
rect 9 507 12 510 
rect 12 0 15 3 
rect 12 3 15 6 
rect 12 6 15 9 
rect 12 9 15 12 
rect 12 12 15 15 
rect 12 15 15 18 
rect 12 18 15 21 
rect 12 21 15 24 
rect 12 24 15 27 
rect 12 27 15 30 
rect 12 30 15 33 
rect 12 33 15 36 
rect 12 36 15 39 
rect 12 39 15 42 
rect 12 42 15 45 
rect 12 45 15 48 
rect 12 48 15 51 
rect 12 51 15 54 
rect 12 54 15 57 
rect 12 57 15 60 
rect 12 60 15 63 
rect 12 63 15 66 
rect 12 66 15 69 
rect 12 69 15 72 
rect 12 72 15 75 
rect 12 75 15 78 
rect 12 78 15 81 
rect 12 81 15 84 
rect 12 84 15 87 
rect 12 87 15 90 
rect 12 90 15 93 
rect 12 93 15 96 
rect 12 96 15 99 
rect 12 99 15 102 
rect 12 102 15 105 
rect 12 105 15 108 
rect 12 108 15 111 
rect 12 111 15 114 
rect 12 114 15 117 
rect 12 117 15 120 
rect 12 120 15 123 
rect 12 123 15 126 
rect 12 126 15 129 
rect 12 129 15 132 
rect 12 132 15 135 
rect 12 135 15 138 
rect 12 138 15 141 
rect 12 141 15 144 
rect 12 144 15 147 
rect 12 147 15 150 
rect 12 150 15 153 
rect 12 153 15 156 
rect 12 156 15 159 
rect 12 159 15 162 
rect 12 162 15 165 
rect 12 165 15 168 
rect 12 168 15 171 
rect 12 171 15 174 
rect 12 174 15 177 
rect 12 177 15 180 
rect 12 180 15 183 
rect 12 183 15 186 
rect 12 186 15 189 
rect 12 189 15 192 
rect 12 192 15 195 
rect 12 195 15 198 
rect 12 198 15 201 
rect 12 201 15 204 
rect 12 204 15 207 
rect 12 207 15 210 
rect 12 210 15 213 
rect 12 213 15 216 
rect 12 216 15 219 
rect 12 219 15 222 
rect 12 222 15 225 
rect 12 225 15 228 
rect 12 228 15 231 
rect 12 231 15 234 
rect 12 234 15 237 
rect 12 237 15 240 
rect 12 240 15 243 
rect 12 243 15 246 
rect 12 246 15 249 
rect 12 249 15 252 
rect 12 252 15 255 
rect 12 255 15 258 
rect 12 258 15 261 
rect 12 261 15 264 
rect 12 264 15 267 
rect 12 267 15 270 
rect 12 270 15 273 
rect 12 273 15 276 
rect 12 276 15 279 
rect 12 279 15 282 
rect 12 282 15 285 
rect 12 285 15 288 
rect 12 288 15 291 
rect 12 291 15 294 
rect 12 294 15 297 
rect 12 297 15 300 
rect 12 300 15 303 
rect 12 303 15 306 
rect 12 306 15 309 
rect 12 309 15 312 
rect 12 312 15 315 
rect 12 315 15 318 
rect 12 318 15 321 
rect 12 321 15 324 
rect 12 324 15 327 
rect 12 327 15 330 
rect 12 330 15 333 
rect 12 333 15 336 
rect 12 336 15 339 
rect 12 339 15 342 
rect 12 342 15 345 
rect 12 345 15 348 
rect 12 348 15 351 
rect 12 351 15 354 
rect 12 354 15 357 
rect 12 357 15 360 
rect 12 360 15 363 
rect 12 363 15 366 
rect 12 366 15 369 
rect 12 369 15 372 
rect 12 372 15 375 
rect 12 375 15 378 
rect 12 378 15 381 
rect 12 381 15 384 
rect 12 384 15 387 
rect 12 387 15 390 
rect 12 390 15 393 
rect 12 393 15 396 
rect 12 396 15 399 
rect 12 399 15 402 
rect 12 402 15 405 
rect 12 405 15 408 
rect 12 408 15 411 
rect 12 411 15 414 
rect 12 414 15 417 
rect 12 417 15 420 
rect 12 420 15 423 
rect 12 423 15 426 
rect 12 426 15 429 
rect 12 429 15 432 
rect 12 432 15 435 
rect 12 435 15 438 
rect 12 438 15 441 
rect 12 441 15 444 
rect 12 444 15 447 
rect 12 447 15 450 
rect 12 450 15 453 
rect 12 453 15 456 
rect 12 456 15 459 
rect 12 459 15 462 
rect 12 462 15 465 
rect 12 465 15 468 
rect 12 468 15 471 
rect 12 471 15 474 
rect 12 474 15 477 
rect 12 477 15 480 
rect 12 480 15 483 
rect 12 483 15 486 
rect 12 486 15 489 
rect 12 489 15 492 
rect 12 492 15 495 
rect 12 495 15 498 
rect 12 498 15 501 
rect 12 501 15 504 
rect 12 504 15 507 
rect 12 507 15 510 
rect 15 0 18 3 
rect 15 3 18 6 
rect 15 6 18 9 
rect 15 9 18 12 
rect 15 12 18 15 
rect 15 15 18 18 
rect 15 18 18 21 
rect 15 21 18 24 
rect 15 24 18 27 
rect 15 27 18 30 
rect 15 30 18 33 
rect 15 33 18 36 
rect 15 36 18 39 
rect 15 39 18 42 
rect 15 42 18 45 
rect 15 45 18 48 
rect 15 48 18 51 
rect 15 51 18 54 
rect 15 54 18 57 
rect 15 57 18 60 
rect 15 60 18 63 
rect 15 63 18 66 
rect 15 66 18 69 
rect 15 69 18 72 
rect 15 72 18 75 
rect 15 75 18 78 
rect 15 78 18 81 
rect 15 81 18 84 
rect 15 84 18 87 
rect 15 87 18 90 
rect 15 90 18 93 
rect 15 93 18 96 
rect 15 96 18 99 
rect 15 99 18 102 
rect 15 102 18 105 
rect 15 105 18 108 
rect 15 108 18 111 
rect 15 111 18 114 
rect 15 114 18 117 
rect 15 117 18 120 
rect 15 120 18 123 
rect 15 123 18 126 
rect 15 126 18 129 
rect 15 129 18 132 
rect 15 132 18 135 
rect 15 135 18 138 
rect 15 138 18 141 
rect 15 141 18 144 
rect 15 144 18 147 
rect 15 147 18 150 
rect 15 150 18 153 
rect 15 153 18 156 
rect 15 156 18 159 
rect 15 159 18 162 
rect 15 162 18 165 
rect 15 165 18 168 
rect 15 168 18 171 
rect 15 171 18 174 
rect 15 174 18 177 
rect 15 177 18 180 
rect 15 180 18 183 
rect 15 183 18 186 
rect 15 186 18 189 
rect 15 189 18 192 
rect 15 192 18 195 
rect 15 195 18 198 
rect 15 198 18 201 
rect 15 201 18 204 
rect 15 204 18 207 
rect 15 207 18 210 
rect 15 210 18 213 
rect 15 213 18 216 
rect 15 216 18 219 
rect 15 219 18 222 
rect 15 222 18 225 
rect 15 225 18 228 
rect 15 228 18 231 
rect 15 231 18 234 
rect 15 234 18 237 
rect 15 237 18 240 
rect 15 240 18 243 
rect 15 243 18 246 
rect 15 246 18 249 
rect 15 249 18 252 
rect 15 252 18 255 
rect 15 255 18 258 
rect 15 258 18 261 
rect 15 261 18 264 
rect 15 264 18 267 
rect 15 267 18 270 
rect 15 270 18 273 
rect 15 273 18 276 
rect 15 276 18 279 
rect 15 279 18 282 
rect 15 282 18 285 
rect 15 285 18 288 
rect 15 288 18 291 
rect 15 291 18 294 
rect 15 294 18 297 
rect 15 297 18 300 
rect 15 300 18 303 
rect 15 303 18 306 
rect 15 306 18 309 
rect 15 309 18 312 
rect 15 312 18 315 
rect 15 315 18 318 
rect 15 318 18 321 
rect 15 321 18 324 
rect 15 324 18 327 
rect 15 327 18 330 
rect 15 330 18 333 
rect 15 333 18 336 
rect 15 336 18 339 
rect 15 339 18 342 
rect 15 342 18 345 
rect 15 345 18 348 
rect 15 348 18 351 
rect 15 351 18 354 
rect 15 354 18 357 
rect 15 357 18 360 
rect 15 360 18 363 
rect 15 363 18 366 
rect 15 366 18 369 
rect 15 369 18 372 
rect 15 372 18 375 
rect 15 375 18 378 
rect 15 378 18 381 
rect 15 381 18 384 
rect 15 384 18 387 
rect 15 387 18 390 
rect 15 390 18 393 
rect 15 393 18 396 
rect 15 396 18 399 
rect 15 399 18 402 
rect 15 402 18 405 
rect 15 405 18 408 
rect 15 408 18 411 
rect 15 411 18 414 
rect 15 414 18 417 
rect 15 417 18 420 
rect 15 420 18 423 
rect 15 423 18 426 
rect 15 426 18 429 
rect 15 429 18 432 
rect 15 432 18 435 
rect 15 435 18 438 
rect 15 438 18 441 
rect 15 441 18 444 
rect 15 444 18 447 
rect 15 447 18 450 
rect 15 450 18 453 
rect 15 453 18 456 
rect 15 456 18 459 
rect 15 459 18 462 
rect 15 462 18 465 
rect 15 465 18 468 
rect 15 468 18 471 
rect 15 471 18 474 
rect 15 474 18 477 
rect 15 477 18 480 
rect 15 480 18 483 
rect 15 483 18 486 
rect 15 486 18 489 
rect 15 489 18 492 
rect 15 492 18 495 
rect 15 495 18 498 
rect 15 498 18 501 
rect 15 501 18 504 
rect 15 504 18 507 
rect 15 507 18 510 
rect 18 0 21 3 
rect 18 3 21 6 
rect 18 6 21 9 
rect 18 9 21 12 
rect 18 12 21 15 
rect 18 15 21 18 
rect 18 18 21 21 
rect 18 21 21 24 
rect 18 24 21 27 
rect 18 27 21 30 
rect 18 30 21 33 
rect 18 33 21 36 
rect 18 36 21 39 
rect 18 39 21 42 
rect 18 42 21 45 
rect 18 45 21 48 
rect 18 48 21 51 
rect 18 51 21 54 
rect 18 54 21 57 
rect 18 57 21 60 
rect 18 60 21 63 
rect 18 63 21 66 
rect 18 66 21 69 
rect 18 69 21 72 
rect 18 72 21 75 
rect 18 75 21 78 
rect 18 78 21 81 
rect 18 81 21 84 
rect 18 84 21 87 
rect 18 87 21 90 
rect 18 90 21 93 
rect 18 93 21 96 
rect 18 96 21 99 
rect 18 99 21 102 
rect 18 102 21 105 
rect 18 105 21 108 
rect 18 108 21 111 
rect 18 111 21 114 
rect 18 114 21 117 
rect 18 117 21 120 
rect 18 120 21 123 
rect 18 123 21 126 
rect 18 126 21 129 
rect 18 129 21 132 
rect 18 132 21 135 
rect 18 135 21 138 
rect 18 138 21 141 
rect 18 141 21 144 
rect 18 144 21 147 
rect 18 147 21 150 
rect 18 150 21 153 
rect 18 153 21 156 
rect 18 156 21 159 
rect 18 159 21 162 
rect 18 162 21 165 
rect 18 165 21 168 
rect 18 168 21 171 
rect 18 171 21 174 
rect 18 174 21 177 
rect 18 177 21 180 
rect 18 180 21 183 
rect 18 183 21 186 
rect 18 186 21 189 
rect 18 189 21 192 
rect 18 192 21 195 
rect 18 195 21 198 
rect 18 198 21 201 
rect 18 201 21 204 
rect 18 204 21 207 
rect 18 207 21 210 
rect 18 210 21 213 
rect 18 213 21 216 
rect 18 216 21 219 
rect 18 219 21 222 
rect 18 222 21 225 
rect 18 225 21 228 
rect 18 228 21 231 
rect 18 231 21 234 
rect 18 234 21 237 
rect 18 237 21 240 
rect 18 240 21 243 
rect 18 243 21 246 
rect 18 246 21 249 
rect 18 249 21 252 
rect 18 252 21 255 
rect 18 255 21 258 
rect 18 258 21 261 
rect 18 261 21 264 
rect 18 264 21 267 
rect 18 267 21 270 
rect 18 270 21 273 
rect 18 273 21 276 
rect 18 276 21 279 
rect 18 279 21 282 
rect 18 282 21 285 
rect 18 285 21 288 
rect 18 288 21 291 
rect 18 291 21 294 
rect 18 294 21 297 
rect 18 297 21 300 
rect 18 300 21 303 
rect 18 303 21 306 
rect 18 306 21 309 
rect 18 309 21 312 
rect 18 312 21 315 
rect 18 315 21 318 
rect 18 318 21 321 
rect 18 321 21 324 
rect 18 324 21 327 
rect 18 327 21 330 
rect 18 330 21 333 
rect 18 333 21 336 
rect 18 336 21 339 
rect 18 339 21 342 
rect 18 342 21 345 
rect 18 345 21 348 
rect 18 348 21 351 
rect 18 351 21 354 
rect 18 354 21 357 
rect 18 357 21 360 
rect 18 360 21 363 
rect 18 363 21 366 
rect 18 366 21 369 
rect 18 369 21 372 
rect 18 372 21 375 
rect 18 375 21 378 
rect 18 378 21 381 
rect 18 381 21 384 
rect 18 384 21 387 
rect 18 387 21 390 
rect 18 390 21 393 
rect 18 393 21 396 
rect 18 396 21 399 
rect 18 399 21 402 
rect 18 402 21 405 
rect 18 405 21 408 
rect 18 408 21 411 
rect 18 411 21 414 
rect 18 414 21 417 
rect 18 417 21 420 
rect 18 420 21 423 
rect 18 423 21 426 
rect 18 426 21 429 
rect 18 429 21 432 
rect 18 432 21 435 
rect 18 435 21 438 
rect 18 438 21 441 
rect 18 441 21 444 
rect 18 444 21 447 
rect 18 447 21 450 
rect 18 450 21 453 
rect 18 453 21 456 
rect 18 456 21 459 
rect 18 459 21 462 
rect 18 462 21 465 
rect 18 465 21 468 
rect 18 468 21 471 
rect 18 471 21 474 
rect 18 474 21 477 
rect 18 477 21 480 
rect 18 480 21 483 
rect 18 483 21 486 
rect 18 486 21 489 
rect 18 489 21 492 
rect 18 492 21 495 
rect 18 495 21 498 
rect 18 498 21 501 
rect 18 501 21 504 
rect 18 504 21 507 
rect 18 507 21 510 
rect 21 0 24 3 
rect 21 3 24 6 
rect 21 6 24 9 
rect 21 9 24 12 
rect 21 12 24 15 
rect 21 15 24 18 
rect 21 18 24 21 
rect 21 21 24 24 
rect 21 24 24 27 
rect 21 27 24 30 
rect 21 30 24 33 
rect 21 33 24 36 
rect 21 36 24 39 
rect 21 39 24 42 
rect 21 42 24 45 
rect 21 45 24 48 
rect 21 48 24 51 
rect 21 51 24 54 
rect 21 54 24 57 
rect 21 57 24 60 
rect 21 60 24 63 
rect 21 63 24 66 
rect 21 66 24 69 
rect 21 69 24 72 
rect 21 72 24 75 
rect 21 75 24 78 
rect 21 78 24 81 
rect 21 81 24 84 
rect 21 84 24 87 
rect 21 87 24 90 
rect 21 90 24 93 
rect 21 93 24 96 
rect 21 96 24 99 
rect 21 99 24 102 
rect 21 102 24 105 
rect 21 105 24 108 
rect 21 108 24 111 
rect 21 111 24 114 
rect 21 114 24 117 
rect 21 117 24 120 
rect 21 120 24 123 
rect 21 123 24 126 
rect 21 126 24 129 
rect 21 129 24 132 
rect 21 132 24 135 
rect 21 135 24 138 
rect 21 138 24 141 
rect 21 141 24 144 
rect 21 144 24 147 
rect 21 147 24 150 
rect 21 150 24 153 
rect 21 153 24 156 
rect 21 156 24 159 
rect 21 159 24 162 
rect 21 162 24 165 
rect 21 165 24 168 
rect 21 168 24 171 
rect 21 171 24 174 
rect 21 174 24 177 
rect 21 177 24 180 
rect 21 180 24 183 
rect 21 183 24 186 
rect 21 186 24 189 
rect 21 189 24 192 
rect 21 192 24 195 
rect 21 195 24 198 
rect 21 198 24 201 
rect 21 201 24 204 
rect 21 204 24 207 
rect 21 207 24 210 
rect 21 210 24 213 
rect 21 213 24 216 
rect 21 216 24 219 
rect 21 219 24 222 
rect 21 222 24 225 
rect 21 225 24 228 
rect 21 228 24 231 
rect 21 231 24 234 
rect 21 234 24 237 
rect 21 237 24 240 
rect 21 240 24 243 
rect 21 243 24 246 
rect 21 246 24 249 
rect 21 249 24 252 
rect 21 252 24 255 
rect 21 255 24 258 
rect 21 258 24 261 
rect 21 261 24 264 
rect 21 264 24 267 
rect 21 267 24 270 
rect 21 270 24 273 
rect 21 273 24 276 
rect 21 276 24 279 
rect 21 279 24 282 
rect 21 282 24 285 
rect 21 285 24 288 
rect 21 288 24 291 
rect 21 291 24 294 
rect 21 294 24 297 
rect 21 297 24 300 
rect 21 300 24 303 
rect 21 303 24 306 
rect 21 306 24 309 
rect 21 309 24 312 
rect 21 312 24 315 
rect 21 315 24 318 
rect 21 318 24 321 
rect 21 321 24 324 
rect 21 324 24 327 
rect 21 327 24 330 
rect 21 330 24 333 
rect 21 333 24 336 
rect 21 336 24 339 
rect 21 339 24 342 
rect 21 342 24 345 
rect 21 345 24 348 
rect 21 348 24 351 
rect 21 351 24 354 
rect 21 354 24 357 
rect 21 357 24 360 
rect 21 360 24 363 
rect 21 363 24 366 
rect 21 366 24 369 
rect 21 369 24 372 
rect 21 372 24 375 
rect 21 375 24 378 
rect 21 378 24 381 
rect 21 381 24 384 
rect 21 384 24 387 
rect 21 387 24 390 
rect 21 390 24 393 
rect 21 393 24 396 
rect 21 396 24 399 
rect 21 399 24 402 
rect 21 402 24 405 
rect 21 405 24 408 
rect 21 408 24 411 
rect 21 411 24 414 
rect 21 414 24 417 
rect 21 417 24 420 
rect 21 420 24 423 
rect 21 423 24 426 
rect 21 426 24 429 
rect 21 429 24 432 
rect 21 432 24 435 
rect 21 435 24 438 
rect 21 438 24 441 
rect 21 441 24 444 
rect 21 444 24 447 
rect 21 447 24 450 
rect 21 450 24 453 
rect 21 453 24 456 
rect 21 456 24 459 
rect 21 459 24 462 
rect 21 462 24 465 
rect 21 465 24 468 
rect 21 468 24 471 
rect 21 471 24 474 
rect 21 474 24 477 
rect 21 477 24 480 
rect 21 480 24 483 
rect 21 483 24 486 
rect 21 486 24 489 
rect 21 489 24 492 
rect 21 492 24 495 
rect 21 495 24 498 
rect 21 498 24 501 
rect 21 501 24 504 
rect 21 504 24 507 
rect 21 507 24 510 
rect 24 0 27 3 
rect 24 3 27 6 
rect 24 6 27 9 
rect 24 9 27 12 
rect 24 12 27 15 
rect 24 15 27 18 
rect 24 18 27 21 
rect 24 21 27 24 
rect 24 24 27 27 
rect 24 27 27 30 
rect 24 30 27 33 
rect 24 33 27 36 
rect 24 36 27 39 
rect 24 39 27 42 
rect 24 42 27 45 
rect 24 45 27 48 
rect 24 48 27 51 
rect 24 51 27 54 
rect 24 54 27 57 
rect 24 57 27 60 
rect 24 60 27 63 
rect 24 63 27 66 
rect 24 66 27 69 
rect 24 69 27 72 
rect 24 72 27 75 
rect 24 75 27 78 
rect 24 78 27 81 
rect 24 81 27 84 
rect 24 84 27 87 
rect 24 87 27 90 
rect 24 90 27 93 
rect 24 93 27 96 
rect 24 96 27 99 
rect 24 99 27 102 
rect 24 102 27 105 
rect 24 105 27 108 
rect 24 108 27 111 
rect 24 111 27 114 
rect 24 114 27 117 
rect 24 117 27 120 
rect 24 120 27 123 
rect 24 123 27 126 
rect 24 126 27 129 
rect 24 129 27 132 
rect 24 132 27 135 
rect 24 135 27 138 
rect 24 138 27 141 
rect 24 141 27 144 
rect 24 144 27 147 
rect 24 147 27 150 
rect 24 150 27 153 
rect 24 153 27 156 
rect 24 156 27 159 
rect 24 159 27 162 
rect 24 162 27 165 
rect 24 165 27 168 
rect 24 168 27 171 
rect 24 171 27 174 
rect 24 174 27 177 
rect 24 177 27 180 
rect 24 180 27 183 
rect 24 183 27 186 
rect 24 186 27 189 
rect 24 189 27 192 
rect 24 192 27 195 
rect 24 195 27 198 
rect 24 198 27 201 
rect 24 201 27 204 
rect 24 204 27 207 
rect 24 207 27 210 
rect 24 210 27 213 
rect 24 213 27 216 
rect 24 216 27 219 
rect 24 219 27 222 
rect 24 222 27 225 
rect 24 225 27 228 
rect 24 228 27 231 
rect 24 231 27 234 
rect 24 234 27 237 
rect 24 237 27 240 
rect 24 240 27 243 
rect 24 243 27 246 
rect 24 246 27 249 
rect 24 249 27 252 
rect 24 252 27 255 
rect 24 255 27 258 
rect 24 258 27 261 
rect 24 261 27 264 
rect 24 264 27 267 
rect 24 267 27 270 
rect 24 270 27 273 
rect 24 273 27 276 
rect 24 276 27 279 
rect 24 279 27 282 
rect 24 282 27 285 
rect 24 285 27 288 
rect 24 288 27 291 
rect 24 291 27 294 
rect 24 294 27 297 
rect 24 297 27 300 
rect 24 300 27 303 
rect 24 303 27 306 
rect 24 306 27 309 
rect 24 309 27 312 
rect 24 312 27 315 
rect 24 315 27 318 
rect 24 318 27 321 
rect 24 321 27 324 
rect 24 324 27 327 
rect 24 327 27 330 
rect 24 330 27 333 
rect 24 333 27 336 
rect 24 336 27 339 
rect 24 339 27 342 
rect 24 342 27 345 
rect 24 345 27 348 
rect 24 348 27 351 
rect 24 351 27 354 
rect 24 354 27 357 
rect 24 357 27 360 
rect 24 360 27 363 
rect 24 363 27 366 
rect 24 366 27 369 
rect 24 369 27 372 
rect 24 372 27 375 
rect 24 375 27 378 
rect 24 378 27 381 
rect 24 381 27 384 
rect 24 384 27 387 
rect 24 387 27 390 
rect 24 390 27 393 
rect 24 393 27 396 
rect 24 396 27 399 
rect 24 399 27 402 
rect 24 402 27 405 
rect 24 405 27 408 
rect 24 408 27 411 
rect 24 411 27 414 
rect 24 414 27 417 
rect 24 417 27 420 
rect 24 420 27 423 
rect 24 423 27 426 
rect 24 426 27 429 
rect 24 429 27 432 
rect 24 432 27 435 
rect 24 435 27 438 
rect 24 438 27 441 
rect 24 441 27 444 
rect 24 444 27 447 
rect 24 447 27 450 
rect 24 450 27 453 
rect 24 453 27 456 
rect 24 456 27 459 
rect 24 459 27 462 
rect 24 462 27 465 
rect 24 465 27 468 
rect 24 468 27 471 
rect 24 471 27 474 
rect 24 474 27 477 
rect 24 477 27 480 
rect 24 480 27 483 
rect 24 483 27 486 
rect 24 486 27 489 
rect 24 489 27 492 
rect 24 492 27 495 
rect 24 495 27 498 
rect 24 498 27 501 
rect 24 501 27 504 
rect 24 504 27 507 
rect 24 507 27 510 
rect 27 0 30 3 
rect 27 3 30 6 
rect 27 6 30 9 
rect 27 9 30 12 
rect 27 12 30 15 
rect 27 15 30 18 
rect 27 18 30 21 
rect 27 21 30 24 
rect 27 24 30 27 
rect 27 27 30 30 
rect 27 30 30 33 
rect 27 33 30 36 
rect 27 36 30 39 
rect 27 39 30 42 
rect 27 42 30 45 
rect 27 45 30 48 
rect 27 48 30 51 
rect 27 51 30 54 
rect 27 54 30 57 
rect 27 57 30 60 
rect 27 60 30 63 
rect 27 63 30 66 
rect 27 66 30 69 
rect 27 69 30 72 
rect 27 72 30 75 
rect 27 75 30 78 
rect 27 78 30 81 
rect 27 81 30 84 
rect 27 84 30 87 
rect 27 87 30 90 
rect 27 90 30 93 
rect 27 93 30 96 
rect 27 96 30 99 
rect 27 99 30 102 
rect 27 102 30 105 
rect 27 105 30 108 
rect 27 108 30 111 
rect 27 111 30 114 
rect 27 114 30 117 
rect 27 117 30 120 
rect 27 120 30 123 
rect 27 123 30 126 
rect 27 126 30 129 
rect 27 129 30 132 
rect 27 132 30 135 
rect 27 135 30 138 
rect 27 138 30 141 
rect 27 141 30 144 
rect 27 144 30 147 
rect 27 147 30 150 
rect 27 150 30 153 
rect 27 153 30 156 
rect 27 156 30 159 
rect 27 159 30 162 
rect 27 162 30 165 
rect 27 165 30 168 
rect 27 168 30 171 
rect 27 171 30 174 
rect 27 174 30 177 
rect 27 177 30 180 
rect 27 180 30 183 
rect 27 183 30 186 
rect 27 186 30 189 
rect 27 189 30 192 
rect 27 192 30 195 
rect 27 195 30 198 
rect 27 198 30 201 
rect 27 201 30 204 
rect 27 204 30 207 
rect 27 207 30 210 
rect 27 210 30 213 
rect 27 213 30 216 
rect 27 216 30 219 
rect 27 219 30 222 
rect 27 222 30 225 
rect 27 225 30 228 
rect 27 228 30 231 
rect 27 231 30 234 
rect 27 234 30 237 
rect 27 237 30 240 
rect 27 240 30 243 
rect 27 243 30 246 
rect 27 246 30 249 
rect 27 249 30 252 
rect 27 252 30 255 
rect 27 255 30 258 
rect 27 258 30 261 
rect 27 261 30 264 
rect 27 264 30 267 
rect 27 267 30 270 
rect 27 270 30 273 
rect 27 273 30 276 
rect 27 276 30 279 
rect 27 279 30 282 
rect 27 282 30 285 
rect 27 285 30 288 
rect 27 288 30 291 
rect 27 291 30 294 
rect 27 294 30 297 
rect 27 297 30 300 
rect 27 300 30 303 
rect 27 303 30 306 
rect 27 306 30 309 
rect 27 309 30 312 
rect 27 312 30 315 
rect 27 315 30 318 
rect 27 318 30 321 
rect 27 321 30 324 
rect 27 324 30 327 
rect 27 327 30 330 
rect 27 330 30 333 
rect 27 333 30 336 
rect 27 336 30 339 
rect 27 339 30 342 
rect 27 342 30 345 
rect 27 345 30 348 
rect 27 348 30 351 
rect 27 351 30 354 
rect 27 354 30 357 
rect 27 357 30 360 
rect 27 360 30 363 
rect 27 363 30 366 
rect 27 366 30 369 
rect 27 369 30 372 
rect 27 372 30 375 
rect 27 375 30 378 
rect 27 378 30 381 
rect 27 381 30 384 
rect 27 384 30 387 
rect 27 387 30 390 
rect 27 390 30 393 
rect 27 393 30 396 
rect 27 396 30 399 
rect 27 399 30 402 
rect 27 402 30 405 
rect 27 405 30 408 
rect 27 408 30 411 
rect 27 411 30 414 
rect 27 414 30 417 
rect 27 417 30 420 
rect 27 420 30 423 
rect 27 423 30 426 
rect 27 426 30 429 
rect 27 429 30 432 
rect 27 432 30 435 
rect 27 435 30 438 
rect 27 438 30 441 
rect 27 441 30 444 
rect 27 444 30 447 
rect 27 447 30 450 
rect 27 450 30 453 
rect 27 453 30 456 
rect 27 456 30 459 
rect 27 459 30 462 
rect 27 462 30 465 
rect 27 465 30 468 
rect 27 468 30 471 
rect 27 471 30 474 
rect 27 474 30 477 
rect 27 477 30 480 
rect 27 480 30 483 
rect 27 483 30 486 
rect 27 486 30 489 
rect 27 489 30 492 
rect 27 492 30 495 
rect 27 495 30 498 
rect 27 498 30 501 
rect 27 501 30 504 
rect 27 504 30 507 
rect 27 507 30 510 
rect 30 0 33 3 
rect 30 3 33 6 
rect 30 6 33 9 
rect 30 9 33 12 
rect 30 12 33 15 
rect 30 15 33 18 
rect 30 18 33 21 
rect 30 21 33 24 
rect 30 24 33 27 
rect 30 27 33 30 
rect 30 30 33 33 
rect 30 33 33 36 
rect 30 36 33 39 
rect 30 39 33 42 
rect 30 42 33 45 
rect 30 45 33 48 
rect 30 48 33 51 
rect 30 51 33 54 
rect 30 54 33 57 
rect 30 57 33 60 
rect 30 60 33 63 
rect 30 63 33 66 
rect 30 66 33 69 
rect 30 69 33 72 
rect 30 72 33 75 
rect 30 75 33 78 
rect 30 78 33 81 
rect 30 81 33 84 
rect 30 84 33 87 
rect 30 87 33 90 
rect 30 90 33 93 
rect 30 93 33 96 
rect 30 96 33 99 
rect 30 99 33 102 
rect 30 102 33 105 
rect 30 105 33 108 
rect 30 108 33 111 
rect 30 111 33 114 
rect 30 114 33 117 
rect 30 117 33 120 
rect 30 120 33 123 
rect 30 123 33 126 
rect 30 126 33 129 
rect 30 129 33 132 
rect 30 132 33 135 
rect 30 135 33 138 
rect 30 138 33 141 
rect 30 141 33 144 
rect 30 144 33 147 
rect 30 147 33 150 
rect 30 150 33 153 
rect 30 153 33 156 
rect 30 156 33 159 
rect 30 159 33 162 
rect 30 162 33 165 
rect 30 165 33 168 
rect 30 168 33 171 
rect 30 171 33 174 
rect 30 174 33 177 
rect 30 177 33 180 
rect 30 180 33 183 
rect 30 183 33 186 
rect 30 186 33 189 
rect 30 189 33 192 
rect 30 192 33 195 
rect 30 195 33 198 
rect 30 198 33 201 
rect 30 201 33 204 
rect 30 204 33 207 
rect 30 207 33 210 
rect 30 210 33 213 
rect 30 213 33 216 
rect 30 216 33 219 
rect 30 219 33 222 
rect 30 222 33 225 
rect 30 225 33 228 
rect 30 228 33 231 
rect 30 231 33 234 
rect 30 234 33 237 
rect 30 237 33 240 
rect 30 240 33 243 
rect 30 243 33 246 
rect 30 246 33 249 
rect 30 249 33 252 
rect 30 252 33 255 
rect 30 255 33 258 
rect 30 258 33 261 
rect 30 261 33 264 
rect 30 264 33 267 
rect 30 267 33 270 
rect 30 270 33 273 
rect 30 273 33 276 
rect 30 276 33 279 
rect 30 279 33 282 
rect 30 282 33 285 
rect 30 285 33 288 
rect 30 288 33 291 
rect 30 291 33 294 
rect 30 294 33 297 
rect 30 297 33 300 
rect 30 300 33 303 
rect 30 303 33 306 
rect 30 306 33 309 
rect 30 309 33 312 
rect 30 312 33 315 
rect 30 315 33 318 
rect 30 318 33 321 
rect 30 321 33 324 
rect 30 324 33 327 
rect 30 327 33 330 
rect 30 330 33 333 
rect 30 333 33 336 
rect 30 336 33 339 
rect 30 339 33 342 
rect 30 342 33 345 
rect 30 345 33 348 
rect 30 348 33 351 
rect 30 351 33 354 
rect 30 354 33 357 
rect 30 357 33 360 
rect 30 360 33 363 
rect 30 363 33 366 
rect 30 366 33 369 
rect 30 369 33 372 
rect 30 372 33 375 
rect 30 375 33 378 
rect 30 378 33 381 
rect 30 381 33 384 
rect 30 384 33 387 
rect 30 387 33 390 
rect 30 390 33 393 
rect 30 393 33 396 
rect 30 396 33 399 
rect 30 399 33 402 
rect 30 402 33 405 
rect 30 405 33 408 
rect 30 408 33 411 
rect 30 411 33 414 
rect 30 414 33 417 
rect 30 417 33 420 
rect 30 420 33 423 
rect 30 423 33 426 
rect 30 426 33 429 
rect 30 429 33 432 
rect 30 432 33 435 
rect 30 435 33 438 
rect 30 438 33 441 
rect 30 441 33 444 
rect 30 444 33 447 
rect 30 447 33 450 
rect 30 450 33 453 
rect 30 453 33 456 
rect 30 456 33 459 
rect 30 459 33 462 
rect 30 462 33 465 
rect 30 465 33 468 
rect 30 468 33 471 
rect 30 471 33 474 
rect 30 474 33 477 
rect 30 477 33 480 
rect 30 480 33 483 
rect 30 483 33 486 
rect 30 486 33 489 
rect 30 489 33 492 
rect 30 492 33 495 
rect 30 495 33 498 
rect 30 498 33 501 
rect 30 501 33 504 
rect 30 504 33 507 
rect 30 507 33 510 
rect 33 0 36 3 
rect 33 3 36 6 
rect 33 6 36 9 
rect 33 9 36 12 
rect 33 12 36 15 
rect 33 15 36 18 
rect 33 18 36 21 
rect 33 21 36 24 
rect 33 24 36 27 
rect 33 27 36 30 
rect 33 30 36 33 
rect 33 33 36 36 
rect 33 36 36 39 
rect 33 39 36 42 
rect 33 42 36 45 
rect 33 45 36 48 
rect 33 48 36 51 
rect 33 51 36 54 
rect 33 54 36 57 
rect 33 57 36 60 
rect 33 60 36 63 
rect 33 63 36 66 
rect 33 66 36 69 
rect 33 69 36 72 
rect 33 72 36 75 
rect 33 75 36 78 
rect 33 78 36 81 
rect 33 81 36 84 
rect 33 84 36 87 
rect 33 87 36 90 
rect 33 90 36 93 
rect 33 93 36 96 
rect 33 96 36 99 
rect 33 99 36 102 
rect 33 102 36 105 
rect 33 105 36 108 
rect 33 108 36 111 
rect 33 111 36 114 
rect 33 114 36 117 
rect 33 117 36 120 
rect 33 120 36 123 
rect 33 123 36 126 
rect 33 126 36 129 
rect 33 129 36 132 
rect 33 132 36 135 
rect 33 135 36 138 
rect 33 138 36 141 
rect 33 141 36 144 
rect 33 144 36 147 
rect 33 147 36 150 
rect 33 150 36 153 
rect 33 153 36 156 
rect 33 156 36 159 
rect 33 159 36 162 
rect 33 162 36 165 
rect 33 165 36 168 
rect 33 168 36 171 
rect 33 171 36 174 
rect 33 174 36 177 
rect 33 177 36 180 
rect 33 180 36 183 
rect 33 183 36 186 
rect 33 186 36 189 
rect 33 189 36 192 
rect 33 192 36 195 
rect 33 195 36 198 
rect 33 198 36 201 
rect 33 201 36 204 
rect 33 204 36 207 
rect 33 207 36 210 
rect 33 210 36 213 
rect 33 213 36 216 
rect 33 216 36 219 
rect 33 219 36 222 
rect 33 222 36 225 
rect 33 225 36 228 
rect 33 228 36 231 
rect 33 231 36 234 
rect 33 234 36 237 
rect 33 237 36 240 
rect 33 240 36 243 
rect 33 243 36 246 
rect 33 246 36 249 
rect 33 249 36 252 
rect 33 252 36 255 
rect 33 255 36 258 
rect 33 258 36 261 
rect 33 261 36 264 
rect 33 264 36 267 
rect 33 267 36 270 
rect 33 270 36 273 
rect 33 273 36 276 
rect 33 276 36 279 
rect 33 279 36 282 
rect 33 282 36 285 
rect 33 285 36 288 
rect 33 288 36 291 
rect 33 291 36 294 
rect 33 294 36 297 
rect 33 297 36 300 
rect 33 300 36 303 
rect 33 303 36 306 
rect 33 306 36 309 
rect 33 309 36 312 
rect 33 312 36 315 
rect 33 315 36 318 
rect 33 318 36 321 
rect 33 321 36 324 
rect 33 324 36 327 
rect 33 327 36 330 
rect 33 330 36 333 
rect 33 333 36 336 
rect 33 336 36 339 
rect 33 339 36 342 
rect 33 342 36 345 
rect 33 345 36 348 
rect 33 348 36 351 
rect 33 351 36 354 
rect 33 354 36 357 
rect 33 357 36 360 
rect 33 360 36 363 
rect 33 363 36 366 
rect 33 366 36 369 
rect 33 369 36 372 
rect 33 372 36 375 
rect 33 375 36 378 
rect 33 378 36 381 
rect 33 381 36 384 
rect 33 384 36 387 
rect 33 387 36 390 
rect 33 390 36 393 
rect 33 393 36 396 
rect 33 396 36 399 
rect 33 399 36 402 
rect 33 402 36 405 
rect 33 405 36 408 
rect 33 408 36 411 
rect 33 411 36 414 
rect 33 414 36 417 
rect 33 417 36 420 
rect 33 420 36 423 
rect 33 423 36 426 
rect 33 426 36 429 
rect 33 429 36 432 
rect 33 432 36 435 
rect 33 435 36 438 
rect 33 438 36 441 
rect 33 441 36 444 
rect 33 444 36 447 
rect 33 447 36 450 
rect 33 450 36 453 
rect 33 453 36 456 
rect 33 456 36 459 
rect 33 459 36 462 
rect 33 462 36 465 
rect 33 465 36 468 
rect 33 468 36 471 
rect 33 471 36 474 
rect 33 474 36 477 
rect 33 477 36 480 
rect 33 480 36 483 
rect 33 483 36 486 
rect 33 486 36 489 
rect 33 489 36 492 
rect 33 492 36 495 
rect 33 495 36 498 
rect 33 498 36 501 
rect 33 501 36 504 
rect 33 504 36 507 
rect 33 507 36 510 
rect 36 0 39 3 
rect 36 3 39 6 
rect 36 6 39 9 
rect 36 9 39 12 
rect 36 12 39 15 
rect 36 15 39 18 
rect 36 18 39 21 
rect 36 21 39 24 
rect 36 24 39 27 
rect 36 27 39 30 
rect 36 30 39 33 
rect 36 33 39 36 
rect 36 36 39 39 
rect 36 39 39 42 
rect 36 42 39 45 
rect 36 45 39 48 
rect 36 48 39 51 
rect 36 51 39 54 
rect 36 54 39 57 
rect 36 57 39 60 
rect 36 60 39 63 
rect 36 63 39 66 
rect 36 66 39 69 
rect 36 69 39 72 
rect 36 72 39 75 
rect 36 75 39 78 
rect 36 78 39 81 
rect 36 81 39 84 
rect 36 84 39 87 
rect 36 87 39 90 
rect 36 90 39 93 
rect 36 93 39 96 
rect 36 96 39 99 
rect 36 99 39 102 
rect 36 102 39 105 
rect 36 105 39 108 
rect 36 108 39 111 
rect 36 111 39 114 
rect 36 114 39 117 
rect 36 117 39 120 
rect 36 120 39 123 
rect 36 123 39 126 
rect 36 126 39 129 
rect 36 129 39 132 
rect 36 132 39 135 
rect 36 135 39 138 
rect 36 138 39 141 
rect 36 141 39 144 
rect 36 144 39 147 
rect 36 147 39 150 
rect 36 150 39 153 
rect 36 153 39 156 
rect 36 156 39 159 
rect 36 159 39 162 
rect 36 162 39 165 
rect 36 165 39 168 
rect 36 168 39 171 
rect 36 171 39 174 
rect 36 174 39 177 
rect 36 177 39 180 
rect 36 180 39 183 
rect 36 183 39 186 
rect 36 186 39 189 
rect 36 189 39 192 
rect 36 192 39 195 
rect 36 195 39 198 
rect 36 198 39 201 
rect 36 201 39 204 
rect 36 204 39 207 
rect 36 207 39 210 
rect 36 210 39 213 
rect 36 213 39 216 
rect 36 216 39 219 
rect 36 219 39 222 
rect 36 222 39 225 
rect 36 225 39 228 
rect 36 228 39 231 
rect 36 231 39 234 
rect 36 234 39 237 
rect 36 237 39 240 
rect 36 240 39 243 
rect 36 243 39 246 
rect 36 246 39 249 
rect 36 249 39 252 
rect 36 252 39 255 
rect 36 255 39 258 
rect 36 258 39 261 
rect 36 261 39 264 
rect 36 264 39 267 
rect 36 267 39 270 
rect 36 270 39 273 
rect 36 273 39 276 
rect 36 276 39 279 
rect 36 279 39 282 
rect 36 282 39 285 
rect 36 285 39 288 
rect 36 288 39 291 
rect 36 291 39 294 
rect 36 294 39 297 
rect 36 297 39 300 
rect 36 300 39 303 
rect 36 303 39 306 
rect 36 306 39 309 
rect 36 309 39 312 
rect 36 312 39 315 
rect 36 315 39 318 
rect 36 318 39 321 
rect 36 321 39 324 
rect 36 324 39 327 
rect 36 327 39 330 
rect 36 330 39 333 
rect 36 333 39 336 
rect 36 336 39 339 
rect 36 339 39 342 
rect 36 342 39 345 
rect 36 345 39 348 
rect 36 348 39 351 
rect 36 351 39 354 
rect 36 354 39 357 
rect 36 357 39 360 
rect 36 360 39 363 
rect 36 363 39 366 
rect 36 366 39 369 
rect 36 369 39 372 
rect 36 372 39 375 
rect 36 375 39 378 
rect 36 378 39 381 
rect 36 381 39 384 
rect 36 384 39 387 
rect 36 387 39 390 
rect 36 390 39 393 
rect 36 393 39 396 
rect 36 396 39 399 
rect 36 399 39 402 
rect 36 402 39 405 
rect 36 405 39 408 
rect 36 408 39 411 
rect 36 411 39 414 
rect 36 414 39 417 
rect 36 417 39 420 
rect 36 420 39 423 
rect 36 423 39 426 
rect 36 426 39 429 
rect 36 429 39 432 
rect 36 432 39 435 
rect 36 435 39 438 
rect 36 438 39 441 
rect 36 441 39 444 
rect 36 444 39 447 
rect 36 447 39 450 
rect 36 450 39 453 
rect 36 453 39 456 
rect 36 456 39 459 
rect 36 459 39 462 
rect 36 462 39 465 
rect 36 465 39 468 
rect 36 468 39 471 
rect 36 471 39 474 
rect 36 474 39 477 
rect 36 477 39 480 
rect 36 480 39 483 
rect 36 483 39 486 
rect 36 486 39 489 
rect 36 489 39 492 
rect 36 492 39 495 
rect 36 495 39 498 
rect 36 498 39 501 
rect 36 501 39 504 
rect 36 504 39 507 
rect 36 507 39 510 
rect 39 0 42 3 
rect 39 3 42 6 
rect 39 6 42 9 
rect 39 9 42 12 
rect 39 12 42 15 
rect 39 15 42 18 
rect 39 18 42 21 
rect 39 21 42 24 
rect 39 24 42 27 
rect 39 27 42 30 
rect 39 30 42 33 
rect 39 33 42 36 
rect 39 36 42 39 
rect 39 39 42 42 
rect 39 42 42 45 
rect 39 45 42 48 
rect 39 48 42 51 
rect 39 51 42 54 
rect 39 54 42 57 
rect 39 57 42 60 
rect 39 60 42 63 
rect 39 63 42 66 
rect 39 66 42 69 
rect 39 69 42 72 
rect 39 72 42 75 
rect 39 75 42 78 
rect 39 78 42 81 
rect 39 81 42 84 
rect 39 84 42 87 
rect 39 87 42 90 
rect 39 90 42 93 
rect 39 93 42 96 
rect 39 96 42 99 
rect 39 99 42 102 
rect 39 102 42 105 
rect 39 105 42 108 
rect 39 108 42 111 
rect 39 111 42 114 
rect 39 114 42 117 
rect 39 117 42 120 
rect 39 120 42 123 
rect 39 123 42 126 
rect 39 126 42 129 
rect 39 129 42 132 
rect 39 132 42 135 
rect 39 135 42 138 
rect 39 138 42 141 
rect 39 141 42 144 
rect 39 144 42 147 
rect 39 147 42 150 
rect 39 150 42 153 
rect 39 153 42 156 
rect 39 156 42 159 
rect 39 159 42 162 
rect 39 162 42 165 
rect 39 165 42 168 
rect 39 168 42 171 
rect 39 171 42 174 
rect 39 174 42 177 
rect 39 177 42 180 
rect 39 180 42 183 
rect 39 183 42 186 
rect 39 186 42 189 
rect 39 189 42 192 
rect 39 192 42 195 
rect 39 195 42 198 
rect 39 198 42 201 
rect 39 201 42 204 
rect 39 204 42 207 
rect 39 207 42 210 
rect 39 210 42 213 
rect 39 213 42 216 
rect 39 216 42 219 
rect 39 219 42 222 
rect 39 222 42 225 
rect 39 225 42 228 
rect 39 228 42 231 
rect 39 231 42 234 
rect 39 234 42 237 
rect 39 237 42 240 
rect 39 240 42 243 
rect 39 243 42 246 
rect 39 246 42 249 
rect 39 249 42 252 
rect 39 252 42 255 
rect 39 255 42 258 
rect 39 258 42 261 
rect 39 261 42 264 
rect 39 264 42 267 
rect 39 267 42 270 
rect 39 270 42 273 
rect 39 273 42 276 
rect 39 276 42 279 
rect 39 279 42 282 
rect 39 282 42 285 
rect 39 285 42 288 
rect 39 288 42 291 
rect 39 291 42 294 
rect 39 294 42 297 
rect 39 297 42 300 
rect 39 300 42 303 
rect 39 303 42 306 
rect 39 306 42 309 
rect 39 309 42 312 
rect 39 312 42 315 
rect 39 315 42 318 
rect 39 318 42 321 
rect 39 321 42 324 
rect 39 324 42 327 
rect 39 327 42 330 
rect 39 330 42 333 
rect 39 333 42 336 
rect 39 336 42 339 
rect 39 339 42 342 
rect 39 342 42 345 
rect 39 345 42 348 
rect 39 348 42 351 
rect 39 351 42 354 
rect 39 354 42 357 
rect 39 357 42 360 
rect 39 360 42 363 
rect 39 363 42 366 
rect 39 366 42 369 
rect 39 369 42 372 
rect 39 372 42 375 
rect 39 375 42 378 
rect 39 378 42 381 
rect 39 381 42 384 
rect 39 384 42 387 
rect 39 387 42 390 
rect 39 390 42 393 
rect 39 393 42 396 
rect 39 396 42 399 
rect 39 399 42 402 
rect 39 402 42 405 
rect 39 405 42 408 
rect 39 408 42 411 
rect 39 411 42 414 
rect 39 414 42 417 
rect 39 417 42 420 
rect 39 420 42 423 
rect 39 423 42 426 
rect 39 426 42 429 
rect 39 429 42 432 
rect 39 432 42 435 
rect 39 435 42 438 
rect 39 438 42 441 
rect 39 441 42 444 
rect 39 444 42 447 
rect 39 447 42 450 
rect 39 450 42 453 
rect 39 453 42 456 
rect 39 456 42 459 
rect 39 459 42 462 
rect 39 462 42 465 
rect 39 465 42 468 
rect 39 468 42 471 
rect 39 471 42 474 
rect 39 474 42 477 
rect 39 477 42 480 
rect 39 480 42 483 
rect 39 483 42 486 
rect 39 486 42 489 
rect 39 489 42 492 
rect 39 492 42 495 
rect 39 495 42 498 
rect 39 498 42 501 
rect 39 501 42 504 
rect 39 504 42 507 
rect 39 507 42 510 
rect 42 0 45 3 
rect 42 3 45 6 
rect 42 6 45 9 
rect 42 9 45 12 
rect 42 12 45 15 
rect 42 15 45 18 
rect 42 18 45 21 
rect 42 21 45 24 
rect 42 24 45 27 
rect 42 27 45 30 
rect 42 30 45 33 
rect 42 33 45 36 
rect 42 36 45 39 
rect 42 39 45 42 
rect 42 42 45 45 
rect 42 45 45 48 
rect 42 48 45 51 
rect 42 51 45 54 
rect 42 54 45 57 
rect 42 57 45 60 
rect 42 60 45 63 
rect 42 63 45 66 
rect 42 66 45 69 
rect 42 69 45 72 
rect 42 72 45 75 
rect 42 75 45 78 
rect 42 78 45 81 
rect 42 81 45 84 
rect 42 84 45 87 
rect 42 87 45 90 
rect 42 90 45 93 
rect 42 93 45 96 
rect 42 96 45 99 
rect 42 99 45 102 
rect 42 102 45 105 
rect 42 105 45 108 
rect 42 108 45 111 
rect 42 111 45 114 
rect 42 114 45 117 
rect 42 117 45 120 
rect 42 120 45 123 
rect 42 123 45 126 
rect 42 126 45 129 
rect 42 129 45 132 
rect 42 132 45 135 
rect 42 135 45 138 
rect 42 138 45 141 
rect 42 141 45 144 
rect 42 144 45 147 
rect 42 147 45 150 
rect 42 150 45 153 
rect 42 153 45 156 
rect 42 156 45 159 
rect 42 159 45 162 
rect 42 162 45 165 
rect 42 165 45 168 
rect 42 168 45 171 
rect 42 171 45 174 
rect 42 174 45 177 
rect 42 177 45 180 
rect 42 180 45 183 
rect 42 183 45 186 
rect 42 186 45 189 
rect 42 189 45 192 
rect 42 192 45 195 
rect 42 195 45 198 
rect 42 198 45 201 
rect 42 201 45 204 
rect 42 204 45 207 
rect 42 207 45 210 
rect 42 210 45 213 
rect 42 213 45 216 
rect 42 216 45 219 
rect 42 219 45 222 
rect 42 222 45 225 
rect 42 225 45 228 
rect 42 228 45 231 
rect 42 231 45 234 
rect 42 234 45 237 
rect 42 237 45 240 
rect 42 240 45 243 
rect 42 243 45 246 
rect 42 246 45 249 
rect 42 249 45 252 
rect 42 252 45 255 
rect 42 255 45 258 
rect 42 258 45 261 
rect 42 261 45 264 
rect 42 264 45 267 
rect 42 267 45 270 
rect 42 270 45 273 
rect 42 273 45 276 
rect 42 276 45 279 
rect 42 279 45 282 
rect 42 282 45 285 
rect 42 285 45 288 
rect 42 288 45 291 
rect 42 291 45 294 
rect 42 294 45 297 
rect 42 297 45 300 
rect 42 300 45 303 
rect 42 303 45 306 
rect 42 306 45 309 
rect 42 309 45 312 
rect 42 312 45 315 
rect 42 315 45 318 
rect 42 318 45 321 
rect 42 321 45 324 
rect 42 324 45 327 
rect 42 327 45 330 
rect 42 330 45 333 
rect 42 333 45 336 
rect 42 336 45 339 
rect 42 339 45 342 
rect 42 342 45 345 
rect 42 345 45 348 
rect 42 348 45 351 
rect 42 351 45 354 
rect 42 354 45 357 
rect 42 357 45 360 
rect 42 360 45 363 
rect 42 363 45 366 
rect 42 366 45 369 
rect 42 369 45 372 
rect 42 372 45 375 
rect 42 375 45 378 
rect 42 378 45 381 
rect 42 381 45 384 
rect 42 384 45 387 
rect 42 387 45 390 
rect 42 390 45 393 
rect 42 393 45 396 
rect 42 396 45 399 
rect 42 399 45 402 
rect 42 402 45 405 
rect 42 405 45 408 
rect 42 408 45 411 
rect 42 411 45 414 
rect 42 414 45 417 
rect 42 417 45 420 
rect 42 420 45 423 
rect 42 423 45 426 
rect 42 426 45 429 
rect 42 429 45 432 
rect 42 432 45 435 
rect 42 435 45 438 
rect 42 438 45 441 
rect 42 441 45 444 
rect 42 444 45 447 
rect 42 447 45 450 
rect 42 450 45 453 
rect 42 453 45 456 
rect 42 456 45 459 
rect 42 459 45 462 
rect 42 462 45 465 
rect 42 465 45 468 
rect 42 468 45 471 
rect 42 471 45 474 
rect 42 474 45 477 
rect 42 477 45 480 
rect 42 480 45 483 
rect 42 483 45 486 
rect 42 486 45 489 
rect 42 489 45 492 
rect 42 492 45 495 
rect 42 495 45 498 
rect 42 498 45 501 
rect 42 501 45 504 
rect 42 504 45 507 
rect 42 507 45 510 
rect 45 0 48 3 
rect 45 3 48 6 
rect 45 6 48 9 
rect 45 9 48 12 
rect 45 12 48 15 
rect 45 15 48 18 
rect 45 18 48 21 
rect 45 21 48 24 
rect 45 24 48 27 
rect 45 27 48 30 
rect 45 30 48 33 
rect 45 33 48 36 
rect 45 36 48 39 
rect 45 39 48 42 
rect 45 42 48 45 
rect 45 45 48 48 
rect 45 48 48 51 
rect 45 51 48 54 
rect 45 54 48 57 
rect 45 57 48 60 
rect 45 60 48 63 
rect 45 63 48 66 
rect 45 66 48 69 
rect 45 69 48 72 
rect 45 72 48 75 
rect 45 75 48 78 
rect 45 78 48 81 
rect 45 81 48 84 
rect 45 84 48 87 
rect 45 87 48 90 
rect 45 90 48 93 
rect 45 93 48 96 
rect 45 96 48 99 
rect 45 99 48 102 
rect 45 102 48 105 
rect 45 105 48 108 
rect 45 108 48 111 
rect 45 111 48 114 
rect 45 114 48 117 
rect 45 117 48 120 
rect 45 120 48 123 
rect 45 123 48 126 
rect 45 126 48 129 
rect 45 129 48 132 
rect 45 132 48 135 
rect 45 135 48 138 
rect 45 138 48 141 
rect 45 141 48 144 
rect 45 144 48 147 
rect 45 147 48 150 
rect 45 150 48 153 
rect 45 153 48 156 
rect 45 156 48 159 
rect 45 159 48 162 
rect 45 162 48 165 
rect 45 165 48 168 
rect 45 168 48 171 
rect 45 171 48 174 
rect 45 174 48 177 
rect 45 177 48 180 
rect 45 180 48 183 
rect 45 183 48 186 
rect 45 186 48 189 
rect 45 189 48 192 
rect 45 192 48 195 
rect 45 195 48 198 
rect 45 198 48 201 
rect 45 201 48 204 
rect 45 204 48 207 
rect 45 207 48 210 
rect 45 210 48 213 
rect 45 213 48 216 
rect 45 216 48 219 
rect 45 219 48 222 
rect 45 222 48 225 
rect 45 225 48 228 
rect 45 228 48 231 
rect 45 231 48 234 
rect 45 234 48 237 
rect 45 237 48 240 
rect 45 240 48 243 
rect 45 243 48 246 
rect 45 246 48 249 
rect 45 249 48 252 
rect 45 252 48 255 
rect 45 255 48 258 
rect 45 258 48 261 
rect 45 261 48 264 
rect 45 264 48 267 
rect 45 267 48 270 
rect 45 270 48 273 
rect 45 273 48 276 
rect 45 276 48 279 
rect 45 279 48 282 
rect 45 282 48 285 
rect 45 285 48 288 
rect 45 288 48 291 
rect 45 291 48 294 
rect 45 294 48 297 
rect 45 297 48 300 
rect 45 300 48 303 
rect 45 303 48 306 
rect 45 306 48 309 
rect 45 309 48 312 
rect 45 312 48 315 
rect 45 315 48 318 
rect 45 318 48 321 
rect 45 321 48 324 
rect 45 324 48 327 
rect 45 327 48 330 
rect 45 330 48 333 
rect 45 333 48 336 
rect 45 336 48 339 
rect 45 339 48 342 
rect 45 342 48 345 
rect 45 345 48 348 
rect 45 348 48 351 
rect 45 351 48 354 
rect 45 354 48 357 
rect 45 357 48 360 
rect 45 360 48 363 
rect 45 363 48 366 
rect 45 366 48 369 
rect 45 369 48 372 
rect 45 372 48 375 
rect 45 375 48 378 
rect 45 378 48 381 
rect 45 381 48 384 
rect 45 384 48 387 
rect 45 387 48 390 
rect 45 390 48 393 
rect 45 393 48 396 
rect 45 396 48 399 
rect 45 399 48 402 
rect 45 402 48 405 
rect 45 405 48 408 
rect 45 408 48 411 
rect 45 411 48 414 
rect 45 414 48 417 
rect 45 417 48 420 
rect 45 420 48 423 
rect 45 423 48 426 
rect 45 426 48 429 
rect 45 429 48 432 
rect 45 432 48 435 
rect 45 435 48 438 
rect 45 438 48 441 
rect 45 441 48 444 
rect 45 444 48 447 
rect 45 447 48 450 
rect 45 450 48 453 
rect 45 453 48 456 
rect 45 456 48 459 
rect 45 459 48 462 
rect 45 462 48 465 
rect 45 465 48 468 
rect 45 468 48 471 
rect 45 471 48 474 
rect 45 474 48 477 
rect 45 477 48 480 
rect 45 480 48 483 
rect 45 483 48 486 
rect 45 486 48 489 
rect 45 489 48 492 
rect 45 492 48 495 
rect 45 495 48 498 
rect 45 498 48 501 
rect 45 501 48 504 
rect 45 504 48 507 
rect 45 507 48 510 
rect 48 0 51 3 
rect 48 3 51 6 
rect 48 6 51 9 
rect 48 9 51 12 
rect 48 12 51 15 
rect 48 15 51 18 
rect 48 18 51 21 
rect 48 21 51 24 
rect 48 24 51 27 
rect 48 27 51 30 
rect 48 30 51 33 
rect 48 33 51 36 
rect 48 36 51 39 
rect 48 39 51 42 
rect 48 42 51 45 
rect 48 45 51 48 
rect 48 48 51 51 
rect 48 51 51 54 
rect 48 54 51 57 
rect 48 57 51 60 
rect 48 60 51 63 
rect 48 63 51 66 
rect 48 66 51 69 
rect 48 69 51 72 
rect 48 72 51 75 
rect 48 75 51 78 
rect 48 78 51 81 
rect 48 81 51 84 
rect 48 84 51 87 
rect 48 87 51 90 
rect 48 90 51 93 
rect 48 93 51 96 
rect 48 96 51 99 
rect 48 99 51 102 
rect 48 102 51 105 
rect 48 105 51 108 
rect 48 108 51 111 
rect 48 111 51 114 
rect 48 114 51 117 
rect 48 117 51 120 
rect 48 120 51 123 
rect 48 123 51 126 
rect 48 126 51 129 
rect 48 129 51 132 
rect 48 132 51 135 
rect 48 135 51 138 
rect 48 138 51 141 
rect 48 141 51 144 
rect 48 144 51 147 
rect 48 147 51 150 
rect 48 150 51 153 
rect 48 153 51 156 
rect 48 156 51 159 
rect 48 159 51 162 
rect 48 162 51 165 
rect 48 165 51 168 
rect 48 168 51 171 
rect 48 171 51 174 
rect 48 174 51 177 
rect 48 177 51 180 
rect 48 180 51 183 
rect 48 183 51 186 
rect 48 186 51 189 
rect 48 189 51 192 
rect 48 192 51 195 
rect 48 195 51 198 
rect 48 198 51 201 
rect 48 201 51 204 
rect 48 204 51 207 
rect 48 207 51 210 
rect 48 210 51 213 
rect 48 213 51 216 
rect 48 216 51 219 
rect 48 219 51 222 
rect 48 222 51 225 
rect 48 225 51 228 
rect 48 228 51 231 
rect 48 231 51 234 
rect 48 234 51 237 
rect 48 237 51 240 
rect 48 240 51 243 
rect 48 243 51 246 
rect 48 246 51 249 
rect 48 249 51 252 
rect 48 252 51 255 
rect 48 255 51 258 
rect 48 258 51 261 
rect 48 261 51 264 
rect 48 264 51 267 
rect 48 267 51 270 
rect 48 270 51 273 
rect 48 273 51 276 
rect 48 276 51 279 
rect 48 279 51 282 
rect 48 282 51 285 
rect 48 285 51 288 
rect 48 288 51 291 
rect 48 291 51 294 
rect 48 294 51 297 
rect 48 297 51 300 
rect 48 300 51 303 
rect 48 303 51 306 
rect 48 306 51 309 
rect 48 309 51 312 
rect 48 312 51 315 
rect 48 315 51 318 
rect 48 318 51 321 
rect 48 321 51 324 
rect 48 324 51 327 
rect 48 327 51 330 
rect 48 330 51 333 
rect 48 333 51 336 
rect 48 336 51 339 
rect 48 339 51 342 
rect 48 342 51 345 
rect 48 345 51 348 
rect 48 348 51 351 
rect 48 351 51 354 
rect 48 354 51 357 
rect 48 357 51 360 
rect 48 360 51 363 
rect 48 363 51 366 
rect 48 366 51 369 
rect 48 369 51 372 
rect 48 372 51 375 
rect 48 375 51 378 
rect 48 378 51 381 
rect 48 381 51 384 
rect 48 384 51 387 
rect 48 387 51 390 
rect 48 390 51 393 
rect 48 393 51 396 
rect 48 396 51 399 
rect 48 399 51 402 
rect 48 402 51 405 
rect 48 405 51 408 
rect 48 408 51 411 
rect 48 411 51 414 
rect 48 414 51 417 
rect 48 417 51 420 
rect 48 420 51 423 
rect 48 423 51 426 
rect 48 426 51 429 
rect 48 429 51 432 
rect 48 432 51 435 
rect 48 435 51 438 
rect 48 438 51 441 
rect 48 441 51 444 
rect 48 444 51 447 
rect 48 447 51 450 
rect 48 450 51 453 
rect 48 453 51 456 
rect 48 456 51 459 
rect 48 459 51 462 
rect 48 462 51 465 
rect 48 465 51 468 
rect 48 468 51 471 
rect 48 471 51 474 
rect 48 474 51 477 
rect 48 477 51 480 
rect 48 480 51 483 
rect 48 483 51 486 
rect 48 486 51 489 
rect 48 489 51 492 
rect 48 492 51 495 
rect 48 495 51 498 
rect 48 498 51 501 
rect 48 501 51 504 
rect 48 504 51 507 
rect 48 507 51 510 
rect 51 0 54 3 
rect 51 3 54 6 
rect 51 6 54 9 
rect 51 9 54 12 
rect 51 12 54 15 
rect 51 15 54 18 
rect 51 18 54 21 
rect 51 21 54 24 
rect 51 24 54 27 
rect 51 27 54 30 
rect 51 30 54 33 
rect 51 33 54 36 
rect 51 36 54 39 
rect 51 39 54 42 
rect 51 42 54 45 
rect 51 45 54 48 
rect 51 48 54 51 
rect 51 51 54 54 
rect 51 54 54 57 
rect 51 57 54 60 
rect 51 60 54 63 
rect 51 63 54 66 
rect 51 66 54 69 
rect 51 69 54 72 
rect 51 72 54 75 
rect 51 75 54 78 
rect 51 78 54 81 
rect 51 81 54 84 
rect 51 84 54 87 
rect 51 87 54 90 
rect 51 90 54 93 
rect 51 93 54 96 
rect 51 96 54 99 
rect 51 99 54 102 
rect 51 102 54 105 
rect 51 105 54 108 
rect 51 108 54 111 
rect 51 111 54 114 
rect 51 114 54 117 
rect 51 117 54 120 
rect 51 120 54 123 
rect 51 123 54 126 
rect 51 126 54 129 
rect 51 129 54 132 
rect 51 132 54 135 
rect 51 135 54 138 
rect 51 138 54 141 
rect 51 141 54 144 
rect 51 144 54 147 
rect 51 147 54 150 
rect 51 150 54 153 
rect 51 153 54 156 
rect 51 156 54 159 
rect 51 159 54 162 
rect 51 162 54 165 
rect 51 165 54 168 
rect 51 168 54 171 
rect 51 171 54 174 
rect 51 174 54 177 
rect 51 177 54 180 
rect 51 180 54 183 
rect 51 183 54 186 
rect 51 186 54 189 
rect 51 189 54 192 
rect 51 192 54 195 
rect 51 195 54 198 
rect 51 198 54 201 
rect 51 201 54 204 
rect 51 204 54 207 
rect 51 207 54 210 
rect 51 210 54 213 
rect 51 213 54 216 
rect 51 216 54 219 
rect 51 219 54 222 
rect 51 222 54 225 
rect 51 225 54 228 
rect 51 228 54 231 
rect 51 231 54 234 
rect 51 234 54 237 
rect 51 237 54 240 
rect 51 240 54 243 
rect 51 243 54 246 
rect 51 246 54 249 
rect 51 249 54 252 
rect 51 252 54 255 
rect 51 255 54 258 
rect 51 258 54 261 
rect 51 261 54 264 
rect 51 264 54 267 
rect 51 267 54 270 
rect 51 270 54 273 
rect 51 273 54 276 
rect 51 276 54 279 
rect 51 279 54 282 
rect 51 282 54 285 
rect 51 285 54 288 
rect 51 288 54 291 
rect 51 291 54 294 
rect 51 294 54 297 
rect 51 297 54 300 
rect 51 300 54 303 
rect 51 303 54 306 
rect 51 306 54 309 
rect 51 309 54 312 
rect 51 312 54 315 
rect 51 315 54 318 
rect 51 318 54 321 
rect 51 321 54 324 
rect 51 324 54 327 
rect 51 327 54 330 
rect 51 330 54 333 
rect 51 333 54 336 
rect 51 336 54 339 
rect 51 339 54 342 
rect 51 342 54 345 
rect 51 345 54 348 
rect 51 348 54 351 
rect 51 351 54 354 
rect 51 354 54 357 
rect 51 357 54 360 
rect 51 360 54 363 
rect 51 363 54 366 
rect 51 366 54 369 
rect 51 369 54 372 
rect 51 372 54 375 
rect 51 375 54 378 
rect 51 378 54 381 
rect 51 381 54 384 
rect 51 384 54 387 
rect 51 387 54 390 
rect 51 390 54 393 
rect 51 393 54 396 
rect 51 396 54 399 
rect 51 399 54 402 
rect 51 402 54 405 
rect 51 405 54 408 
rect 51 408 54 411 
rect 51 411 54 414 
rect 51 414 54 417 
rect 51 417 54 420 
rect 51 420 54 423 
rect 51 423 54 426 
rect 51 426 54 429 
rect 51 429 54 432 
rect 51 432 54 435 
rect 51 435 54 438 
rect 51 438 54 441 
rect 51 441 54 444 
rect 51 444 54 447 
rect 51 447 54 450 
rect 51 450 54 453 
rect 51 453 54 456 
rect 51 456 54 459 
rect 51 459 54 462 
rect 51 462 54 465 
rect 51 465 54 468 
rect 51 468 54 471 
rect 51 471 54 474 
rect 51 474 54 477 
rect 51 477 54 480 
rect 51 480 54 483 
rect 51 483 54 486 
rect 51 486 54 489 
rect 51 489 54 492 
rect 51 492 54 495 
rect 51 495 54 498 
rect 51 498 54 501 
rect 51 501 54 504 
rect 51 504 54 507 
rect 51 507 54 510 
rect 54 0 57 3 
rect 54 3 57 6 
rect 54 6 57 9 
rect 54 9 57 12 
rect 54 12 57 15 
rect 54 15 57 18 
rect 54 18 57 21 
rect 54 21 57 24 
rect 54 24 57 27 
rect 54 27 57 30 
rect 54 30 57 33 
rect 54 33 57 36 
rect 54 36 57 39 
rect 54 39 57 42 
rect 54 42 57 45 
rect 54 45 57 48 
rect 54 48 57 51 
rect 54 51 57 54 
rect 54 54 57 57 
rect 54 57 57 60 
rect 54 60 57 63 
rect 54 63 57 66 
rect 54 66 57 69 
rect 54 69 57 72 
rect 54 72 57 75 
rect 54 75 57 78 
rect 54 78 57 81 
rect 54 81 57 84 
rect 54 84 57 87 
rect 54 87 57 90 
rect 54 90 57 93 
rect 54 93 57 96 
rect 54 96 57 99 
rect 54 99 57 102 
rect 54 102 57 105 
rect 54 105 57 108 
rect 54 108 57 111 
rect 54 111 57 114 
rect 54 114 57 117 
rect 54 117 57 120 
rect 54 120 57 123 
rect 54 123 57 126 
rect 54 126 57 129 
rect 54 129 57 132 
rect 54 132 57 135 
rect 54 135 57 138 
rect 54 138 57 141 
rect 54 141 57 144 
rect 54 144 57 147 
rect 54 147 57 150 
rect 54 150 57 153 
rect 54 153 57 156 
rect 54 156 57 159 
rect 54 159 57 162 
rect 54 162 57 165 
rect 54 165 57 168 
rect 54 168 57 171 
rect 54 171 57 174 
rect 54 174 57 177 
rect 54 177 57 180 
rect 54 180 57 183 
rect 54 183 57 186 
rect 54 186 57 189 
rect 54 189 57 192 
rect 54 192 57 195 
rect 54 195 57 198 
rect 54 198 57 201 
rect 54 201 57 204 
rect 54 204 57 207 
rect 54 207 57 210 
rect 54 210 57 213 
rect 54 213 57 216 
rect 54 216 57 219 
rect 54 219 57 222 
rect 54 222 57 225 
rect 54 225 57 228 
rect 54 228 57 231 
rect 54 231 57 234 
rect 54 234 57 237 
rect 54 237 57 240 
rect 54 240 57 243 
rect 54 243 57 246 
rect 54 246 57 249 
rect 54 249 57 252 
rect 54 252 57 255 
rect 54 255 57 258 
rect 54 258 57 261 
rect 54 261 57 264 
rect 54 264 57 267 
rect 54 267 57 270 
rect 54 270 57 273 
rect 54 273 57 276 
rect 54 276 57 279 
rect 54 279 57 282 
rect 54 282 57 285 
rect 54 285 57 288 
rect 54 288 57 291 
rect 54 291 57 294 
rect 54 294 57 297 
rect 54 297 57 300 
rect 54 300 57 303 
rect 54 303 57 306 
rect 54 306 57 309 
rect 54 309 57 312 
rect 54 312 57 315 
rect 54 315 57 318 
rect 54 318 57 321 
rect 54 321 57 324 
rect 54 324 57 327 
rect 54 327 57 330 
rect 54 330 57 333 
rect 54 333 57 336 
rect 54 336 57 339 
rect 54 339 57 342 
rect 54 342 57 345 
rect 54 345 57 348 
rect 54 348 57 351 
rect 54 351 57 354 
rect 54 354 57 357 
rect 54 357 57 360 
rect 54 360 57 363 
rect 54 363 57 366 
rect 54 366 57 369 
rect 54 369 57 372 
rect 54 372 57 375 
rect 54 375 57 378 
rect 54 378 57 381 
rect 54 381 57 384 
rect 54 384 57 387 
rect 54 387 57 390 
rect 54 390 57 393 
rect 54 393 57 396 
rect 54 396 57 399 
rect 54 399 57 402 
rect 54 402 57 405 
rect 54 405 57 408 
rect 54 408 57 411 
rect 54 411 57 414 
rect 54 414 57 417 
rect 54 417 57 420 
rect 54 420 57 423 
rect 54 423 57 426 
rect 54 426 57 429 
rect 54 429 57 432 
rect 54 432 57 435 
rect 54 435 57 438 
rect 54 438 57 441 
rect 54 441 57 444 
rect 54 444 57 447 
rect 54 447 57 450 
rect 54 450 57 453 
rect 54 453 57 456 
rect 54 456 57 459 
rect 54 459 57 462 
rect 54 462 57 465 
rect 54 465 57 468 
rect 54 468 57 471 
rect 54 471 57 474 
rect 54 474 57 477 
rect 54 477 57 480 
rect 54 480 57 483 
rect 54 483 57 486 
rect 54 486 57 489 
rect 54 489 57 492 
rect 54 492 57 495 
rect 54 495 57 498 
rect 54 498 57 501 
rect 54 501 57 504 
rect 54 504 57 507 
rect 54 507 57 510 
rect 57 0 60 3 
rect 57 3 60 6 
rect 57 6 60 9 
rect 57 9 60 12 
rect 57 12 60 15 
rect 57 15 60 18 
rect 57 18 60 21 
rect 57 21 60 24 
rect 57 24 60 27 
rect 57 27 60 30 
rect 57 30 60 33 
rect 57 33 60 36 
rect 57 36 60 39 
rect 57 39 60 42 
rect 57 42 60 45 
rect 57 45 60 48 
rect 57 48 60 51 
rect 57 51 60 54 
rect 57 54 60 57 
rect 57 57 60 60 
rect 57 60 60 63 
rect 57 63 60 66 
rect 57 66 60 69 
rect 57 69 60 72 
rect 57 72 60 75 
rect 57 75 60 78 
rect 57 78 60 81 
rect 57 81 60 84 
rect 57 84 60 87 
rect 57 87 60 90 
rect 57 90 60 93 
rect 57 93 60 96 
rect 57 96 60 99 
rect 57 99 60 102 
rect 57 102 60 105 
rect 57 105 60 108 
rect 57 108 60 111 
rect 57 111 60 114 
rect 57 114 60 117 
rect 57 117 60 120 
rect 57 120 60 123 
rect 57 123 60 126 
rect 57 126 60 129 
rect 57 129 60 132 
rect 57 132 60 135 
rect 57 135 60 138 
rect 57 138 60 141 
rect 57 141 60 144 
rect 57 144 60 147 
rect 57 147 60 150 
rect 57 150 60 153 
rect 57 153 60 156 
rect 57 156 60 159 
rect 57 159 60 162 
rect 57 162 60 165 
rect 57 165 60 168 
rect 57 168 60 171 
rect 57 171 60 174 
rect 57 174 60 177 
rect 57 177 60 180 
rect 57 180 60 183 
rect 57 183 60 186 
rect 57 186 60 189 
rect 57 189 60 192 
rect 57 192 60 195 
rect 57 195 60 198 
rect 57 198 60 201 
rect 57 201 60 204 
rect 57 204 60 207 
rect 57 207 60 210 
rect 57 210 60 213 
rect 57 213 60 216 
rect 57 216 60 219 
rect 57 219 60 222 
rect 57 222 60 225 
rect 57 225 60 228 
rect 57 228 60 231 
rect 57 231 60 234 
rect 57 234 60 237 
rect 57 237 60 240 
rect 57 240 60 243 
rect 57 243 60 246 
rect 57 246 60 249 
rect 57 249 60 252 
rect 57 252 60 255 
rect 57 255 60 258 
rect 57 258 60 261 
rect 57 261 60 264 
rect 57 264 60 267 
rect 57 267 60 270 
rect 57 270 60 273 
rect 57 273 60 276 
rect 57 276 60 279 
rect 57 279 60 282 
rect 57 282 60 285 
rect 57 285 60 288 
rect 57 288 60 291 
rect 57 291 60 294 
rect 57 294 60 297 
rect 57 297 60 300 
rect 57 300 60 303 
rect 57 303 60 306 
rect 57 306 60 309 
rect 57 309 60 312 
rect 57 312 60 315 
rect 57 315 60 318 
rect 57 318 60 321 
rect 57 321 60 324 
rect 57 324 60 327 
rect 57 327 60 330 
rect 57 330 60 333 
rect 57 333 60 336 
rect 57 336 60 339 
rect 57 339 60 342 
rect 57 342 60 345 
rect 57 345 60 348 
rect 57 348 60 351 
rect 57 351 60 354 
rect 57 354 60 357 
rect 57 357 60 360 
rect 57 360 60 363 
rect 57 363 60 366 
rect 57 366 60 369 
rect 57 369 60 372 
rect 57 372 60 375 
rect 57 375 60 378 
rect 57 378 60 381 
rect 57 381 60 384 
rect 57 384 60 387 
rect 57 387 60 390 
rect 57 390 60 393 
rect 57 393 60 396 
rect 57 396 60 399 
rect 57 399 60 402 
rect 57 402 60 405 
rect 57 405 60 408 
rect 57 408 60 411 
rect 57 411 60 414 
rect 57 414 60 417 
rect 57 417 60 420 
rect 57 420 60 423 
rect 57 423 60 426 
rect 57 426 60 429 
rect 57 429 60 432 
rect 57 432 60 435 
rect 57 435 60 438 
rect 57 438 60 441 
rect 57 441 60 444 
rect 57 444 60 447 
rect 57 447 60 450 
rect 57 450 60 453 
rect 57 453 60 456 
rect 57 456 60 459 
rect 57 459 60 462 
rect 57 462 60 465 
rect 57 465 60 468 
rect 57 468 60 471 
rect 57 471 60 474 
rect 57 474 60 477 
rect 57 477 60 480 
rect 57 480 60 483 
rect 57 483 60 486 
rect 57 486 60 489 
rect 57 489 60 492 
rect 57 492 60 495 
rect 57 495 60 498 
rect 57 498 60 501 
rect 57 501 60 504 
rect 57 504 60 507 
rect 57 507 60 510 
rect 60 0 63 3 
rect 60 3 63 6 
rect 60 6 63 9 
rect 60 9 63 12 
rect 60 12 63 15 
rect 60 15 63 18 
rect 60 18 63 21 
rect 60 21 63 24 
rect 60 24 63 27 
rect 60 27 63 30 
rect 60 30 63 33 
rect 60 33 63 36 
rect 60 36 63 39 
rect 60 39 63 42 
rect 60 42 63 45 
rect 60 45 63 48 
rect 60 48 63 51 
rect 60 51 63 54 
rect 60 54 63 57 
rect 60 57 63 60 
rect 60 60 63 63 
rect 60 63 63 66 
rect 60 66 63 69 
rect 60 69 63 72 
rect 60 72 63 75 
rect 60 75 63 78 
rect 60 78 63 81 
rect 60 81 63 84 
rect 60 84 63 87 
rect 60 87 63 90 
rect 60 90 63 93 
rect 60 93 63 96 
rect 60 96 63 99 
rect 60 99 63 102 
rect 60 102 63 105 
rect 60 105 63 108 
rect 60 108 63 111 
rect 60 111 63 114 
rect 60 114 63 117 
rect 60 117 63 120 
rect 60 120 63 123 
rect 60 123 63 126 
rect 60 126 63 129 
rect 60 129 63 132 
rect 60 132 63 135 
rect 60 135 63 138 
rect 60 138 63 141 
rect 60 141 63 144 
rect 60 144 63 147 
rect 60 147 63 150 
rect 60 150 63 153 
rect 60 153 63 156 
rect 60 156 63 159 
rect 60 159 63 162 
rect 60 162 63 165 
rect 60 165 63 168 
rect 60 168 63 171 
rect 60 171 63 174 
rect 60 174 63 177 
rect 60 177 63 180 
rect 60 180 63 183 
rect 60 183 63 186 
rect 60 186 63 189 
rect 60 189 63 192 
rect 60 192 63 195 
rect 60 195 63 198 
rect 60 198 63 201 
rect 60 201 63 204 
rect 60 204 63 207 
rect 60 207 63 210 
rect 60 210 63 213 
rect 60 213 63 216 
rect 60 216 63 219 
rect 60 219 63 222 
rect 60 222 63 225 
rect 60 225 63 228 
rect 60 228 63 231 
rect 60 231 63 234 
rect 60 234 63 237 
rect 60 237 63 240 
rect 60 240 63 243 
rect 60 243 63 246 
rect 60 246 63 249 
rect 60 249 63 252 
rect 60 252 63 255 
rect 60 255 63 258 
rect 60 258 63 261 
rect 60 261 63 264 
rect 60 264 63 267 
rect 60 267 63 270 
rect 60 270 63 273 
rect 60 273 63 276 
rect 60 276 63 279 
rect 60 279 63 282 
rect 60 282 63 285 
rect 60 285 63 288 
rect 60 288 63 291 
rect 60 291 63 294 
rect 60 294 63 297 
rect 60 297 63 300 
rect 60 300 63 303 
rect 60 303 63 306 
rect 60 306 63 309 
rect 60 309 63 312 
rect 60 312 63 315 
rect 60 315 63 318 
rect 60 318 63 321 
rect 60 321 63 324 
rect 60 324 63 327 
rect 60 327 63 330 
rect 60 330 63 333 
rect 60 333 63 336 
rect 60 336 63 339 
rect 60 339 63 342 
rect 60 342 63 345 
rect 60 345 63 348 
rect 60 348 63 351 
rect 60 351 63 354 
rect 60 354 63 357 
rect 60 357 63 360 
rect 60 360 63 363 
rect 60 363 63 366 
rect 60 366 63 369 
rect 60 369 63 372 
rect 60 372 63 375 
rect 60 375 63 378 
rect 60 378 63 381 
rect 60 381 63 384 
rect 60 384 63 387 
rect 60 387 63 390 
rect 60 390 63 393 
rect 60 393 63 396 
rect 60 396 63 399 
rect 60 399 63 402 
rect 60 402 63 405 
rect 60 405 63 408 
rect 60 408 63 411 
rect 60 411 63 414 
rect 60 414 63 417 
rect 60 417 63 420 
rect 60 420 63 423 
rect 60 423 63 426 
rect 60 426 63 429 
rect 60 429 63 432 
rect 60 432 63 435 
rect 60 435 63 438 
rect 60 438 63 441 
rect 60 441 63 444 
rect 60 444 63 447 
rect 60 447 63 450 
rect 60 450 63 453 
rect 60 453 63 456 
rect 60 456 63 459 
rect 60 459 63 462 
rect 60 462 63 465 
rect 60 465 63 468 
rect 60 468 63 471 
rect 60 471 63 474 
rect 60 474 63 477 
rect 60 477 63 480 
rect 60 480 63 483 
rect 60 483 63 486 
rect 60 486 63 489 
rect 60 489 63 492 
rect 60 492 63 495 
rect 60 495 63 498 
rect 60 498 63 501 
rect 60 501 63 504 
rect 60 504 63 507 
rect 60 507 63 510 
rect 63 0 66 3 
rect 63 3 66 6 
rect 63 6 66 9 
rect 63 9 66 12 
rect 63 12 66 15 
rect 63 15 66 18 
rect 63 18 66 21 
rect 63 21 66 24 
rect 63 24 66 27 
rect 63 27 66 30 
rect 63 30 66 33 
rect 63 33 66 36 
rect 63 36 66 39 
rect 63 39 66 42 
rect 63 42 66 45 
rect 63 45 66 48 
rect 63 48 66 51 
rect 63 51 66 54 
rect 63 54 66 57 
rect 63 57 66 60 
rect 63 60 66 63 
rect 63 63 66 66 
rect 63 66 66 69 
rect 63 69 66 72 
rect 63 72 66 75 
rect 63 75 66 78 
rect 63 78 66 81 
rect 63 81 66 84 
rect 63 84 66 87 
rect 63 87 66 90 
rect 63 90 66 93 
rect 63 93 66 96 
rect 63 96 66 99 
rect 63 99 66 102 
rect 63 102 66 105 
rect 63 105 66 108 
rect 63 108 66 111 
rect 63 111 66 114 
rect 63 114 66 117 
rect 63 117 66 120 
rect 63 120 66 123 
rect 63 123 66 126 
rect 63 126 66 129 
rect 63 129 66 132 
rect 63 132 66 135 
rect 63 135 66 138 
rect 63 138 66 141 
rect 63 141 66 144 
rect 63 144 66 147 
rect 63 147 66 150 
rect 63 150 66 153 
rect 63 153 66 156 
rect 63 156 66 159 
rect 63 159 66 162 
rect 63 162 66 165 
rect 63 165 66 168 
rect 63 168 66 171 
rect 63 171 66 174 
rect 63 174 66 177 
rect 63 177 66 180 
rect 63 180 66 183 
rect 63 183 66 186 
rect 63 186 66 189 
rect 63 189 66 192 
rect 63 192 66 195 
rect 63 195 66 198 
rect 63 198 66 201 
rect 63 201 66 204 
rect 63 204 66 207 
rect 63 207 66 210 
rect 63 210 66 213 
rect 63 213 66 216 
rect 63 216 66 219 
rect 63 219 66 222 
rect 63 222 66 225 
rect 63 225 66 228 
rect 63 228 66 231 
rect 63 231 66 234 
rect 63 234 66 237 
rect 63 237 66 240 
rect 63 240 66 243 
rect 63 243 66 246 
rect 63 246 66 249 
rect 63 249 66 252 
rect 63 252 66 255 
rect 63 255 66 258 
rect 63 258 66 261 
rect 63 261 66 264 
rect 63 264 66 267 
rect 63 267 66 270 
rect 63 270 66 273 
rect 63 273 66 276 
rect 63 276 66 279 
rect 63 279 66 282 
rect 63 282 66 285 
rect 63 285 66 288 
rect 63 288 66 291 
rect 63 291 66 294 
rect 63 294 66 297 
rect 63 297 66 300 
rect 63 300 66 303 
rect 63 303 66 306 
rect 63 306 66 309 
rect 63 309 66 312 
rect 63 312 66 315 
rect 63 315 66 318 
rect 63 318 66 321 
rect 63 321 66 324 
rect 63 324 66 327 
rect 63 327 66 330 
rect 63 330 66 333 
rect 63 333 66 336 
rect 63 336 66 339 
rect 63 339 66 342 
rect 63 342 66 345 
rect 63 345 66 348 
rect 63 348 66 351 
rect 63 351 66 354 
rect 63 354 66 357 
rect 63 357 66 360 
rect 63 360 66 363 
rect 63 363 66 366 
rect 63 366 66 369 
rect 63 369 66 372 
rect 63 372 66 375 
rect 63 375 66 378 
rect 63 378 66 381 
rect 63 381 66 384 
rect 63 384 66 387 
rect 63 387 66 390 
rect 63 390 66 393 
rect 63 393 66 396 
rect 63 396 66 399 
rect 63 399 66 402 
rect 63 402 66 405 
rect 63 405 66 408 
rect 63 408 66 411 
rect 63 411 66 414 
rect 63 414 66 417 
rect 63 417 66 420 
rect 63 420 66 423 
rect 63 423 66 426 
rect 63 426 66 429 
rect 63 429 66 432 
rect 63 432 66 435 
rect 63 435 66 438 
rect 63 438 66 441 
rect 63 441 66 444 
rect 63 444 66 447 
rect 63 447 66 450 
rect 63 450 66 453 
rect 63 453 66 456 
rect 63 456 66 459 
rect 63 459 66 462 
rect 63 462 66 465 
rect 63 465 66 468 
rect 63 468 66 471 
rect 63 471 66 474 
rect 63 474 66 477 
rect 63 477 66 480 
rect 63 480 66 483 
rect 63 483 66 486 
rect 63 486 66 489 
rect 63 489 66 492 
rect 63 492 66 495 
rect 63 495 66 498 
rect 63 498 66 501 
rect 63 501 66 504 
rect 63 504 66 507 
rect 63 507 66 510 
rect 66 0 69 3 
rect 66 3 69 6 
rect 66 6 69 9 
rect 66 9 69 12 
rect 66 12 69 15 
rect 66 15 69 18 
rect 66 18 69 21 
rect 66 21 69 24 
rect 66 24 69 27 
rect 66 27 69 30 
rect 66 30 69 33 
rect 66 33 69 36 
rect 66 36 69 39 
rect 66 39 69 42 
rect 66 42 69 45 
rect 66 45 69 48 
rect 66 48 69 51 
rect 66 51 69 54 
rect 66 54 69 57 
rect 66 57 69 60 
rect 66 60 69 63 
rect 66 63 69 66 
rect 66 66 69 69 
rect 66 69 69 72 
rect 66 72 69 75 
rect 66 75 69 78 
rect 66 78 69 81 
rect 66 81 69 84 
rect 66 84 69 87 
rect 66 87 69 90 
rect 66 90 69 93 
rect 66 93 69 96 
rect 66 96 69 99 
rect 66 99 69 102 
rect 66 102 69 105 
rect 66 105 69 108 
rect 66 108 69 111 
rect 66 111 69 114 
rect 66 114 69 117 
rect 66 117 69 120 
rect 66 120 69 123 
rect 66 123 69 126 
rect 66 126 69 129 
rect 66 129 69 132 
rect 66 132 69 135 
rect 66 135 69 138 
rect 66 138 69 141 
rect 66 141 69 144 
rect 66 144 69 147 
rect 66 147 69 150 
rect 66 150 69 153 
rect 66 153 69 156 
rect 66 156 69 159 
rect 66 159 69 162 
rect 66 162 69 165 
rect 66 165 69 168 
rect 66 168 69 171 
rect 66 171 69 174 
rect 66 174 69 177 
rect 66 177 69 180 
rect 66 180 69 183 
rect 66 183 69 186 
rect 66 186 69 189 
rect 66 189 69 192 
rect 66 192 69 195 
rect 66 195 69 198 
rect 66 198 69 201 
rect 66 201 69 204 
rect 66 204 69 207 
rect 66 207 69 210 
rect 66 210 69 213 
rect 66 213 69 216 
rect 66 216 69 219 
rect 66 219 69 222 
rect 66 222 69 225 
rect 66 225 69 228 
rect 66 228 69 231 
rect 66 231 69 234 
rect 66 234 69 237 
rect 66 237 69 240 
rect 66 240 69 243 
rect 66 243 69 246 
rect 66 246 69 249 
rect 66 249 69 252 
rect 66 252 69 255 
rect 66 255 69 258 
rect 66 258 69 261 
rect 66 261 69 264 
rect 66 264 69 267 
rect 66 267 69 270 
rect 66 270 69 273 
rect 66 273 69 276 
rect 66 276 69 279 
rect 66 279 69 282 
rect 66 282 69 285 
rect 66 285 69 288 
rect 66 288 69 291 
rect 66 291 69 294 
rect 66 294 69 297 
rect 66 297 69 300 
rect 66 300 69 303 
rect 66 303 69 306 
rect 66 306 69 309 
rect 66 309 69 312 
rect 66 312 69 315 
rect 66 315 69 318 
rect 66 318 69 321 
rect 66 321 69 324 
rect 66 324 69 327 
rect 66 327 69 330 
rect 66 330 69 333 
rect 66 333 69 336 
rect 66 336 69 339 
rect 66 339 69 342 
rect 66 342 69 345 
rect 66 345 69 348 
rect 66 348 69 351 
rect 66 351 69 354 
rect 66 354 69 357 
rect 66 357 69 360 
rect 66 360 69 363 
rect 66 363 69 366 
rect 66 366 69 369 
rect 66 369 69 372 
rect 66 372 69 375 
rect 66 375 69 378 
rect 66 378 69 381 
rect 66 381 69 384 
rect 66 384 69 387 
rect 66 387 69 390 
rect 66 390 69 393 
rect 66 393 69 396 
rect 66 396 69 399 
rect 66 399 69 402 
rect 66 402 69 405 
rect 66 405 69 408 
rect 66 408 69 411 
rect 66 411 69 414 
rect 66 414 69 417 
rect 66 417 69 420 
rect 66 420 69 423 
rect 66 423 69 426 
rect 66 426 69 429 
rect 66 429 69 432 
rect 66 432 69 435 
rect 66 435 69 438 
rect 66 438 69 441 
rect 66 441 69 444 
rect 66 444 69 447 
rect 66 447 69 450 
rect 66 450 69 453 
rect 66 453 69 456 
rect 66 456 69 459 
rect 66 459 69 462 
rect 66 462 69 465 
rect 66 465 69 468 
rect 66 468 69 471 
rect 66 471 69 474 
rect 66 474 69 477 
rect 66 477 69 480 
rect 66 480 69 483 
rect 66 483 69 486 
rect 66 486 69 489 
rect 66 489 69 492 
rect 66 492 69 495 
rect 66 495 69 498 
rect 66 498 69 501 
rect 66 501 69 504 
rect 66 504 69 507 
rect 66 507 69 510 
rect 69 0 72 3 
rect 69 3 72 6 
rect 69 6 72 9 
rect 69 9 72 12 
rect 69 12 72 15 
rect 69 15 72 18 
rect 69 18 72 21 
rect 69 21 72 24 
rect 69 24 72 27 
rect 69 27 72 30 
rect 69 30 72 33 
rect 69 33 72 36 
rect 69 36 72 39 
rect 69 39 72 42 
rect 69 42 72 45 
rect 69 45 72 48 
rect 69 48 72 51 
rect 69 51 72 54 
rect 69 54 72 57 
rect 69 57 72 60 
rect 69 60 72 63 
rect 69 63 72 66 
rect 69 66 72 69 
rect 69 69 72 72 
rect 69 72 72 75 
rect 69 75 72 78 
rect 69 78 72 81 
rect 69 81 72 84 
rect 69 84 72 87 
rect 69 87 72 90 
rect 69 90 72 93 
rect 69 93 72 96 
rect 69 96 72 99 
rect 69 99 72 102 
rect 69 102 72 105 
rect 69 105 72 108 
rect 69 108 72 111 
rect 69 111 72 114 
rect 69 114 72 117 
rect 69 117 72 120 
rect 69 120 72 123 
rect 69 123 72 126 
rect 69 126 72 129 
rect 69 129 72 132 
rect 69 132 72 135 
rect 69 135 72 138 
rect 69 138 72 141 
rect 69 141 72 144 
rect 69 144 72 147 
rect 69 147 72 150 
rect 69 150 72 153 
rect 69 153 72 156 
rect 69 156 72 159 
rect 69 159 72 162 
rect 69 162 72 165 
rect 69 165 72 168 
rect 69 168 72 171 
rect 69 171 72 174 
rect 69 174 72 177 
rect 69 177 72 180 
rect 69 180 72 183 
rect 69 183 72 186 
rect 69 186 72 189 
rect 69 189 72 192 
rect 69 192 72 195 
rect 69 195 72 198 
rect 69 198 72 201 
rect 69 201 72 204 
rect 69 204 72 207 
rect 69 207 72 210 
rect 69 210 72 213 
rect 69 213 72 216 
rect 69 216 72 219 
rect 69 219 72 222 
rect 69 222 72 225 
rect 69 225 72 228 
rect 69 228 72 231 
rect 69 231 72 234 
rect 69 234 72 237 
rect 69 237 72 240 
rect 69 240 72 243 
rect 69 243 72 246 
rect 69 246 72 249 
rect 69 249 72 252 
rect 69 252 72 255 
rect 69 255 72 258 
rect 69 258 72 261 
rect 69 261 72 264 
rect 69 264 72 267 
rect 69 267 72 270 
rect 69 270 72 273 
rect 69 273 72 276 
rect 69 276 72 279 
rect 69 279 72 282 
rect 69 282 72 285 
rect 69 285 72 288 
rect 69 288 72 291 
rect 69 291 72 294 
rect 69 294 72 297 
rect 69 297 72 300 
rect 69 300 72 303 
rect 69 303 72 306 
rect 69 306 72 309 
rect 69 309 72 312 
rect 69 312 72 315 
rect 69 315 72 318 
rect 69 318 72 321 
rect 69 321 72 324 
rect 69 324 72 327 
rect 69 327 72 330 
rect 69 330 72 333 
rect 69 333 72 336 
rect 69 336 72 339 
rect 69 339 72 342 
rect 69 342 72 345 
rect 69 345 72 348 
rect 69 348 72 351 
rect 69 351 72 354 
rect 69 354 72 357 
rect 69 357 72 360 
rect 69 360 72 363 
rect 69 363 72 366 
rect 69 366 72 369 
rect 69 369 72 372 
rect 69 372 72 375 
rect 69 375 72 378 
rect 69 378 72 381 
rect 69 381 72 384 
rect 69 384 72 387 
rect 69 387 72 390 
rect 69 390 72 393 
rect 69 393 72 396 
rect 69 396 72 399 
rect 69 399 72 402 
rect 69 402 72 405 
rect 69 405 72 408 
rect 69 408 72 411 
rect 69 411 72 414 
rect 69 414 72 417 
rect 69 417 72 420 
rect 69 420 72 423 
rect 69 423 72 426 
rect 69 426 72 429 
rect 69 429 72 432 
rect 69 432 72 435 
rect 69 435 72 438 
rect 69 438 72 441 
rect 69 441 72 444 
rect 69 444 72 447 
rect 69 447 72 450 
rect 69 450 72 453 
rect 69 453 72 456 
rect 69 456 72 459 
rect 69 459 72 462 
rect 69 462 72 465 
rect 69 465 72 468 
rect 69 468 72 471 
rect 69 471 72 474 
rect 69 474 72 477 
rect 69 477 72 480 
rect 69 480 72 483 
rect 69 483 72 486 
rect 69 486 72 489 
rect 69 489 72 492 
rect 69 492 72 495 
rect 69 495 72 498 
rect 69 498 72 501 
rect 69 501 72 504 
rect 69 504 72 507 
rect 69 507 72 510 
rect 72 0 75 3 
rect 72 3 75 6 
rect 72 6 75 9 
rect 72 9 75 12 
rect 72 12 75 15 
rect 72 15 75 18 
rect 72 18 75 21 
rect 72 21 75 24 
rect 72 24 75 27 
rect 72 27 75 30 
rect 72 30 75 33 
rect 72 33 75 36 
rect 72 36 75 39 
rect 72 39 75 42 
rect 72 42 75 45 
rect 72 45 75 48 
rect 72 48 75 51 
rect 72 51 75 54 
rect 72 54 75 57 
rect 72 57 75 60 
rect 72 60 75 63 
rect 72 63 75 66 
rect 72 66 75 69 
rect 72 69 75 72 
rect 72 72 75 75 
rect 72 75 75 78 
rect 72 78 75 81 
rect 72 81 75 84 
rect 72 84 75 87 
rect 72 87 75 90 
rect 72 90 75 93 
rect 72 93 75 96 
rect 72 96 75 99 
rect 72 99 75 102 
rect 72 102 75 105 
rect 72 105 75 108 
rect 72 108 75 111 
rect 72 111 75 114 
rect 72 114 75 117 
rect 72 117 75 120 
rect 72 120 75 123 
rect 72 123 75 126 
rect 72 126 75 129 
rect 72 129 75 132 
rect 72 132 75 135 
rect 72 135 75 138 
rect 72 138 75 141 
rect 72 141 75 144 
rect 72 144 75 147 
rect 72 147 75 150 
rect 72 150 75 153 
rect 72 153 75 156 
rect 72 156 75 159 
rect 72 159 75 162 
rect 72 162 75 165 
rect 72 165 75 168 
rect 72 168 75 171 
rect 72 171 75 174 
rect 72 174 75 177 
rect 72 177 75 180 
rect 72 180 75 183 
rect 72 183 75 186 
rect 72 186 75 189 
rect 72 189 75 192 
rect 72 192 75 195 
rect 72 195 75 198 
rect 72 198 75 201 
rect 72 201 75 204 
rect 72 204 75 207 
rect 72 207 75 210 
rect 72 210 75 213 
rect 72 213 75 216 
rect 72 216 75 219 
rect 72 219 75 222 
rect 72 222 75 225 
rect 72 225 75 228 
rect 72 228 75 231 
rect 72 231 75 234 
rect 72 234 75 237 
rect 72 237 75 240 
rect 72 240 75 243 
rect 72 243 75 246 
rect 72 246 75 249 
rect 72 249 75 252 
rect 72 252 75 255 
rect 72 255 75 258 
rect 72 258 75 261 
rect 72 261 75 264 
rect 72 264 75 267 
rect 72 267 75 270 
rect 72 270 75 273 
rect 72 273 75 276 
rect 72 276 75 279 
rect 72 279 75 282 
rect 72 282 75 285 
rect 72 285 75 288 
rect 72 288 75 291 
rect 72 291 75 294 
rect 72 294 75 297 
rect 72 297 75 300 
rect 72 300 75 303 
rect 72 303 75 306 
rect 72 306 75 309 
rect 72 309 75 312 
rect 72 312 75 315 
rect 72 315 75 318 
rect 72 318 75 321 
rect 72 321 75 324 
rect 72 324 75 327 
rect 72 327 75 330 
rect 72 330 75 333 
rect 72 333 75 336 
rect 72 336 75 339 
rect 72 339 75 342 
rect 72 342 75 345 
rect 72 345 75 348 
rect 72 348 75 351 
rect 72 351 75 354 
rect 72 354 75 357 
rect 72 357 75 360 
rect 72 360 75 363 
rect 72 363 75 366 
rect 72 366 75 369 
rect 72 369 75 372 
rect 72 372 75 375 
rect 72 375 75 378 
rect 72 378 75 381 
rect 72 381 75 384 
rect 72 384 75 387 
rect 72 387 75 390 
rect 72 390 75 393 
rect 72 393 75 396 
rect 72 396 75 399 
rect 72 399 75 402 
rect 72 402 75 405 
rect 72 405 75 408 
rect 72 408 75 411 
rect 72 411 75 414 
rect 72 414 75 417 
rect 72 417 75 420 
rect 72 420 75 423 
rect 72 423 75 426 
rect 72 426 75 429 
rect 72 429 75 432 
rect 72 432 75 435 
rect 72 435 75 438 
rect 72 438 75 441 
rect 72 441 75 444 
rect 72 444 75 447 
rect 72 447 75 450 
rect 72 450 75 453 
rect 72 453 75 456 
rect 72 456 75 459 
rect 72 459 75 462 
rect 72 462 75 465 
rect 72 465 75 468 
rect 72 468 75 471 
rect 72 471 75 474 
rect 72 474 75 477 
rect 72 477 75 480 
rect 72 480 75 483 
rect 72 483 75 486 
rect 72 486 75 489 
rect 72 489 75 492 
rect 72 492 75 495 
rect 72 495 75 498 
rect 72 498 75 501 
rect 72 501 75 504 
rect 72 504 75 507 
rect 72 507 75 510 
rect 75 0 78 3 
rect 75 3 78 6 
rect 75 6 78 9 
rect 75 9 78 12 
rect 75 12 78 15 
rect 75 15 78 18 
rect 75 18 78 21 
rect 75 21 78 24 
rect 75 24 78 27 
rect 75 27 78 30 
rect 75 30 78 33 
rect 75 33 78 36 
rect 75 36 78 39 
rect 75 39 78 42 
rect 75 42 78 45 
rect 75 45 78 48 
rect 75 48 78 51 
rect 75 51 78 54 
rect 75 54 78 57 
rect 75 57 78 60 
rect 75 60 78 63 
rect 75 63 78 66 
rect 75 66 78 69 
rect 75 69 78 72 
rect 75 72 78 75 
rect 75 75 78 78 
rect 75 78 78 81 
rect 75 81 78 84 
rect 75 84 78 87 
rect 75 87 78 90 
rect 75 90 78 93 
rect 75 93 78 96 
rect 75 96 78 99 
rect 75 99 78 102 
rect 75 102 78 105 
rect 75 105 78 108 
rect 75 108 78 111 
rect 75 111 78 114 
rect 75 114 78 117 
rect 75 117 78 120 
rect 75 120 78 123 
rect 75 123 78 126 
rect 75 126 78 129 
rect 75 129 78 132 
rect 75 132 78 135 
rect 75 135 78 138 
rect 75 138 78 141 
rect 75 141 78 144 
rect 75 144 78 147 
rect 75 147 78 150 
rect 75 150 78 153 
rect 75 153 78 156 
rect 75 156 78 159 
rect 75 159 78 162 
rect 75 162 78 165 
rect 75 165 78 168 
rect 75 168 78 171 
rect 75 171 78 174 
rect 75 174 78 177 
rect 75 177 78 180 
rect 75 180 78 183 
rect 75 183 78 186 
rect 75 186 78 189 
rect 75 189 78 192 
rect 75 192 78 195 
rect 75 195 78 198 
rect 75 198 78 201 
rect 75 201 78 204 
rect 75 204 78 207 
rect 75 207 78 210 
rect 75 210 78 213 
rect 75 213 78 216 
rect 75 216 78 219 
rect 75 219 78 222 
rect 75 222 78 225 
rect 75 225 78 228 
rect 75 228 78 231 
rect 75 231 78 234 
rect 75 234 78 237 
rect 75 237 78 240 
rect 75 240 78 243 
rect 75 243 78 246 
rect 75 246 78 249 
rect 75 249 78 252 
rect 75 252 78 255 
rect 75 255 78 258 
rect 75 258 78 261 
rect 75 261 78 264 
rect 75 264 78 267 
rect 75 267 78 270 
rect 75 270 78 273 
rect 75 273 78 276 
rect 75 276 78 279 
rect 75 279 78 282 
rect 75 282 78 285 
rect 75 285 78 288 
rect 75 288 78 291 
rect 75 291 78 294 
rect 75 294 78 297 
rect 75 297 78 300 
rect 75 300 78 303 
rect 75 303 78 306 
rect 75 306 78 309 
rect 75 309 78 312 
rect 75 312 78 315 
rect 75 315 78 318 
rect 75 318 78 321 
rect 75 321 78 324 
rect 75 324 78 327 
rect 75 327 78 330 
rect 75 330 78 333 
rect 75 333 78 336 
rect 75 336 78 339 
rect 75 339 78 342 
rect 75 342 78 345 
rect 75 345 78 348 
rect 75 348 78 351 
rect 75 351 78 354 
rect 75 354 78 357 
rect 75 357 78 360 
rect 75 360 78 363 
rect 75 363 78 366 
rect 75 366 78 369 
rect 75 369 78 372 
rect 75 372 78 375 
rect 75 375 78 378 
rect 75 378 78 381 
rect 75 381 78 384 
rect 75 384 78 387 
rect 75 387 78 390 
rect 75 390 78 393 
rect 75 393 78 396 
rect 75 396 78 399 
rect 75 399 78 402 
rect 75 402 78 405 
rect 75 405 78 408 
rect 75 408 78 411 
rect 75 411 78 414 
rect 75 414 78 417 
rect 75 417 78 420 
rect 75 420 78 423 
rect 75 423 78 426 
rect 75 426 78 429 
rect 75 429 78 432 
rect 75 432 78 435 
rect 75 435 78 438 
rect 75 438 78 441 
rect 75 441 78 444 
rect 75 444 78 447 
rect 75 447 78 450 
rect 75 450 78 453 
rect 75 453 78 456 
rect 75 456 78 459 
rect 75 459 78 462 
rect 75 462 78 465 
rect 75 465 78 468 
rect 75 468 78 471 
rect 75 471 78 474 
rect 75 474 78 477 
rect 75 477 78 480 
rect 75 480 78 483 
rect 75 483 78 486 
rect 75 486 78 489 
rect 75 489 78 492 
rect 75 492 78 495 
rect 75 495 78 498 
rect 75 498 78 501 
rect 75 501 78 504 
rect 75 504 78 507 
rect 75 507 78 510 
rect 78 0 81 3 
rect 78 3 81 6 
rect 78 6 81 9 
rect 78 9 81 12 
rect 78 12 81 15 
rect 78 15 81 18 
rect 78 18 81 21 
rect 78 21 81 24 
rect 78 24 81 27 
rect 78 27 81 30 
rect 78 30 81 33 
rect 78 33 81 36 
rect 78 36 81 39 
rect 78 39 81 42 
rect 78 42 81 45 
rect 78 45 81 48 
rect 78 48 81 51 
rect 78 51 81 54 
rect 78 54 81 57 
rect 78 57 81 60 
rect 78 60 81 63 
rect 78 63 81 66 
rect 78 66 81 69 
rect 78 69 81 72 
rect 78 72 81 75 
rect 78 75 81 78 
rect 78 78 81 81 
rect 78 81 81 84 
rect 78 84 81 87 
rect 78 87 81 90 
rect 78 90 81 93 
rect 78 93 81 96 
rect 78 96 81 99 
rect 78 99 81 102 
rect 78 102 81 105 
rect 78 105 81 108 
rect 78 108 81 111 
rect 78 111 81 114 
rect 78 114 81 117 
rect 78 117 81 120 
rect 78 120 81 123 
rect 78 123 81 126 
rect 78 126 81 129 
rect 78 129 81 132 
rect 78 132 81 135 
rect 78 135 81 138 
rect 78 138 81 141 
rect 78 141 81 144 
rect 78 144 81 147 
rect 78 147 81 150 
rect 78 150 81 153 
rect 78 153 81 156 
rect 78 156 81 159 
rect 78 159 81 162 
rect 78 162 81 165 
rect 78 165 81 168 
rect 78 168 81 171 
rect 78 171 81 174 
rect 78 174 81 177 
rect 78 177 81 180 
rect 78 180 81 183 
rect 78 183 81 186 
rect 78 186 81 189 
rect 78 189 81 192 
rect 78 192 81 195 
rect 78 195 81 198 
rect 78 198 81 201 
rect 78 201 81 204 
rect 78 204 81 207 
rect 78 207 81 210 
rect 78 210 81 213 
rect 78 213 81 216 
rect 78 216 81 219 
rect 78 219 81 222 
rect 78 222 81 225 
rect 78 225 81 228 
rect 78 228 81 231 
rect 78 231 81 234 
rect 78 234 81 237 
rect 78 237 81 240 
rect 78 240 81 243 
rect 78 243 81 246 
rect 78 246 81 249 
rect 78 249 81 252 
rect 78 252 81 255 
rect 78 255 81 258 
rect 78 258 81 261 
rect 78 261 81 264 
rect 78 264 81 267 
rect 78 267 81 270 
rect 78 270 81 273 
rect 78 273 81 276 
rect 78 276 81 279 
rect 78 279 81 282 
rect 78 282 81 285 
rect 78 285 81 288 
rect 78 288 81 291 
rect 78 291 81 294 
rect 78 294 81 297 
rect 78 297 81 300 
rect 78 300 81 303 
rect 78 303 81 306 
rect 78 306 81 309 
rect 78 309 81 312 
rect 78 312 81 315 
rect 78 315 81 318 
rect 78 318 81 321 
rect 78 321 81 324 
rect 78 324 81 327 
rect 78 327 81 330 
rect 78 330 81 333 
rect 78 333 81 336 
rect 78 336 81 339 
rect 78 339 81 342 
rect 78 342 81 345 
rect 78 345 81 348 
rect 78 348 81 351 
rect 78 351 81 354 
rect 78 354 81 357 
rect 78 357 81 360 
rect 78 360 81 363 
rect 78 363 81 366 
rect 78 366 81 369 
rect 78 369 81 372 
rect 78 372 81 375 
rect 78 375 81 378 
rect 78 378 81 381 
rect 78 381 81 384 
rect 78 384 81 387 
rect 78 387 81 390 
rect 78 390 81 393 
rect 78 393 81 396 
rect 78 396 81 399 
rect 78 399 81 402 
rect 78 402 81 405 
rect 78 405 81 408 
rect 78 408 81 411 
rect 78 411 81 414 
rect 78 414 81 417 
rect 78 417 81 420 
rect 78 420 81 423 
rect 78 423 81 426 
rect 78 426 81 429 
rect 78 429 81 432 
rect 78 432 81 435 
rect 78 435 81 438 
rect 78 438 81 441 
rect 78 441 81 444 
rect 78 444 81 447 
rect 78 447 81 450 
rect 78 450 81 453 
rect 78 453 81 456 
rect 78 456 81 459 
rect 78 459 81 462 
rect 78 462 81 465 
rect 78 465 81 468 
rect 78 468 81 471 
rect 78 471 81 474 
rect 78 474 81 477 
rect 78 477 81 480 
rect 78 480 81 483 
rect 78 483 81 486 
rect 78 486 81 489 
rect 78 489 81 492 
rect 78 492 81 495 
rect 78 495 81 498 
rect 78 498 81 501 
rect 78 501 81 504 
rect 78 504 81 507 
rect 78 507 81 510 
rect 81 0 84 3 
rect 81 3 84 6 
rect 81 6 84 9 
rect 81 9 84 12 
rect 81 12 84 15 
rect 81 15 84 18 
rect 81 18 84 21 
rect 81 21 84 24 
rect 81 24 84 27 
rect 81 27 84 30 
rect 81 30 84 33 
rect 81 33 84 36 
rect 81 36 84 39 
rect 81 39 84 42 
rect 81 42 84 45 
rect 81 45 84 48 
rect 81 48 84 51 
rect 81 51 84 54 
rect 81 54 84 57 
rect 81 57 84 60 
rect 81 60 84 63 
rect 81 63 84 66 
rect 81 66 84 69 
rect 81 69 84 72 
rect 81 72 84 75 
rect 81 75 84 78 
rect 81 78 84 81 
rect 81 81 84 84 
rect 81 84 84 87 
rect 81 87 84 90 
rect 81 90 84 93 
rect 81 93 84 96 
rect 81 96 84 99 
rect 81 99 84 102 
rect 81 102 84 105 
rect 81 105 84 108 
rect 81 108 84 111 
rect 81 111 84 114 
rect 81 114 84 117 
rect 81 117 84 120 
rect 81 120 84 123 
rect 81 123 84 126 
rect 81 126 84 129 
rect 81 129 84 132 
rect 81 132 84 135 
rect 81 135 84 138 
rect 81 138 84 141 
rect 81 141 84 144 
rect 81 144 84 147 
rect 81 147 84 150 
rect 81 150 84 153 
rect 81 153 84 156 
rect 81 156 84 159 
rect 81 159 84 162 
rect 81 162 84 165 
rect 81 165 84 168 
rect 81 168 84 171 
rect 81 171 84 174 
rect 81 174 84 177 
rect 81 177 84 180 
rect 81 180 84 183 
rect 81 183 84 186 
rect 81 186 84 189 
rect 81 189 84 192 
rect 81 192 84 195 
rect 81 195 84 198 
rect 81 198 84 201 
rect 81 201 84 204 
rect 81 204 84 207 
rect 81 207 84 210 
rect 81 210 84 213 
rect 81 213 84 216 
rect 81 216 84 219 
rect 81 219 84 222 
rect 81 222 84 225 
rect 81 225 84 228 
rect 81 228 84 231 
rect 81 231 84 234 
rect 81 234 84 237 
rect 81 237 84 240 
rect 81 240 84 243 
rect 81 243 84 246 
rect 81 246 84 249 
rect 81 249 84 252 
rect 81 252 84 255 
rect 81 255 84 258 
rect 81 258 84 261 
rect 81 261 84 264 
rect 81 264 84 267 
rect 81 267 84 270 
rect 81 270 84 273 
rect 81 273 84 276 
rect 81 276 84 279 
rect 81 279 84 282 
rect 81 282 84 285 
rect 81 285 84 288 
rect 81 288 84 291 
rect 81 291 84 294 
rect 81 294 84 297 
rect 81 297 84 300 
rect 81 300 84 303 
rect 81 303 84 306 
rect 81 306 84 309 
rect 81 309 84 312 
rect 81 312 84 315 
rect 81 315 84 318 
rect 81 318 84 321 
rect 81 321 84 324 
rect 81 324 84 327 
rect 81 327 84 330 
rect 81 330 84 333 
rect 81 333 84 336 
rect 81 336 84 339 
rect 81 339 84 342 
rect 81 342 84 345 
rect 81 345 84 348 
rect 81 348 84 351 
rect 81 351 84 354 
rect 81 354 84 357 
rect 81 357 84 360 
rect 81 360 84 363 
rect 81 363 84 366 
rect 81 366 84 369 
rect 81 369 84 372 
rect 81 372 84 375 
rect 81 375 84 378 
rect 81 378 84 381 
rect 81 381 84 384 
rect 81 384 84 387 
rect 81 387 84 390 
rect 81 390 84 393 
rect 81 393 84 396 
rect 81 396 84 399 
rect 81 399 84 402 
rect 81 402 84 405 
rect 81 405 84 408 
rect 81 408 84 411 
rect 81 411 84 414 
rect 81 414 84 417 
rect 81 417 84 420 
rect 81 420 84 423 
rect 81 423 84 426 
rect 81 426 84 429 
rect 81 429 84 432 
rect 81 432 84 435 
rect 81 435 84 438 
rect 81 438 84 441 
rect 81 441 84 444 
rect 81 444 84 447 
rect 81 447 84 450 
rect 81 450 84 453 
rect 81 453 84 456 
rect 81 456 84 459 
rect 81 459 84 462 
rect 81 462 84 465 
rect 81 465 84 468 
rect 81 468 84 471 
rect 81 471 84 474 
rect 81 474 84 477 
rect 81 477 84 480 
rect 81 480 84 483 
rect 81 483 84 486 
rect 81 486 84 489 
rect 81 489 84 492 
rect 81 492 84 495 
rect 81 495 84 498 
rect 81 498 84 501 
rect 81 501 84 504 
rect 81 504 84 507 
rect 81 507 84 510 
rect 84 0 87 3 
rect 84 3 87 6 
rect 84 6 87 9 
rect 84 9 87 12 
rect 84 12 87 15 
rect 84 15 87 18 
rect 84 18 87 21 
rect 84 21 87 24 
rect 84 24 87 27 
rect 84 27 87 30 
rect 84 30 87 33 
rect 84 33 87 36 
rect 84 36 87 39 
rect 84 39 87 42 
rect 84 42 87 45 
rect 84 45 87 48 
rect 84 48 87 51 
rect 84 51 87 54 
rect 84 54 87 57 
rect 84 57 87 60 
rect 84 60 87 63 
rect 84 63 87 66 
rect 84 66 87 69 
rect 84 69 87 72 
rect 84 72 87 75 
rect 84 75 87 78 
rect 84 78 87 81 
rect 84 81 87 84 
rect 84 84 87 87 
rect 84 87 87 90 
rect 84 90 87 93 
rect 84 93 87 96 
rect 84 96 87 99 
rect 84 99 87 102 
rect 84 102 87 105 
rect 84 105 87 108 
rect 84 108 87 111 
rect 84 111 87 114 
rect 84 114 87 117 
rect 84 117 87 120 
rect 84 120 87 123 
rect 84 123 87 126 
rect 84 126 87 129 
rect 84 129 87 132 
rect 84 132 87 135 
rect 84 135 87 138 
rect 84 138 87 141 
rect 84 141 87 144 
rect 84 144 87 147 
rect 84 147 87 150 
rect 84 150 87 153 
rect 84 153 87 156 
rect 84 156 87 159 
rect 84 159 87 162 
rect 84 162 87 165 
rect 84 165 87 168 
rect 84 168 87 171 
rect 84 171 87 174 
rect 84 174 87 177 
rect 84 177 87 180 
rect 84 180 87 183 
rect 84 183 87 186 
rect 84 186 87 189 
rect 84 189 87 192 
rect 84 192 87 195 
rect 84 195 87 198 
rect 84 198 87 201 
rect 84 201 87 204 
rect 84 204 87 207 
rect 84 207 87 210 
rect 84 210 87 213 
rect 84 213 87 216 
rect 84 216 87 219 
rect 84 219 87 222 
rect 84 222 87 225 
rect 84 225 87 228 
rect 84 228 87 231 
rect 84 231 87 234 
rect 84 234 87 237 
rect 84 237 87 240 
rect 84 240 87 243 
rect 84 243 87 246 
rect 84 246 87 249 
rect 84 249 87 252 
rect 84 252 87 255 
rect 84 255 87 258 
rect 84 258 87 261 
rect 84 261 87 264 
rect 84 264 87 267 
rect 84 267 87 270 
rect 84 270 87 273 
rect 84 273 87 276 
rect 84 276 87 279 
rect 84 279 87 282 
rect 84 282 87 285 
rect 84 285 87 288 
rect 84 288 87 291 
rect 84 291 87 294 
rect 84 294 87 297 
rect 84 297 87 300 
rect 84 300 87 303 
rect 84 303 87 306 
rect 84 306 87 309 
rect 84 309 87 312 
rect 84 312 87 315 
rect 84 315 87 318 
rect 84 318 87 321 
rect 84 321 87 324 
rect 84 324 87 327 
rect 84 327 87 330 
rect 84 330 87 333 
rect 84 333 87 336 
rect 84 336 87 339 
rect 84 339 87 342 
rect 84 342 87 345 
rect 84 345 87 348 
rect 84 348 87 351 
rect 84 351 87 354 
rect 84 354 87 357 
rect 84 357 87 360 
rect 84 360 87 363 
rect 84 363 87 366 
rect 84 366 87 369 
rect 84 369 87 372 
rect 84 372 87 375 
rect 84 375 87 378 
rect 84 378 87 381 
rect 84 381 87 384 
rect 84 384 87 387 
rect 84 387 87 390 
rect 84 390 87 393 
rect 84 393 87 396 
rect 84 396 87 399 
rect 84 399 87 402 
rect 84 402 87 405 
rect 84 405 87 408 
rect 84 408 87 411 
rect 84 411 87 414 
rect 84 414 87 417 
rect 84 417 87 420 
rect 84 420 87 423 
rect 84 423 87 426 
rect 84 426 87 429 
rect 84 429 87 432 
rect 84 432 87 435 
rect 84 435 87 438 
rect 84 438 87 441 
rect 84 441 87 444 
rect 84 444 87 447 
rect 84 447 87 450 
rect 84 450 87 453 
rect 84 453 87 456 
rect 84 456 87 459 
rect 84 459 87 462 
rect 84 462 87 465 
rect 84 465 87 468 
rect 84 468 87 471 
rect 84 471 87 474 
rect 84 474 87 477 
rect 84 477 87 480 
rect 84 480 87 483 
rect 84 483 87 486 
rect 84 486 87 489 
rect 84 489 87 492 
rect 84 492 87 495 
rect 84 495 87 498 
rect 84 498 87 501 
rect 84 501 87 504 
rect 84 504 87 507 
rect 84 507 87 510 
rect 87 0 90 3 
rect 87 3 90 6 
rect 87 6 90 9 
rect 87 9 90 12 
rect 87 12 90 15 
rect 87 15 90 18 
rect 87 18 90 21 
rect 87 21 90 24 
rect 87 24 90 27 
rect 87 27 90 30 
rect 87 30 90 33 
rect 87 33 90 36 
rect 87 36 90 39 
rect 87 39 90 42 
rect 87 42 90 45 
rect 87 45 90 48 
rect 87 48 90 51 
rect 87 51 90 54 
rect 87 54 90 57 
rect 87 57 90 60 
rect 87 60 90 63 
rect 87 63 90 66 
rect 87 66 90 69 
rect 87 69 90 72 
rect 87 72 90 75 
rect 87 75 90 78 
rect 87 78 90 81 
rect 87 81 90 84 
rect 87 84 90 87 
rect 87 87 90 90 
rect 87 90 90 93 
rect 87 93 90 96 
rect 87 96 90 99 
rect 87 99 90 102 
rect 87 102 90 105 
rect 87 105 90 108 
rect 87 108 90 111 
rect 87 111 90 114 
rect 87 114 90 117 
rect 87 117 90 120 
rect 87 120 90 123 
rect 87 123 90 126 
rect 87 126 90 129 
rect 87 129 90 132 
rect 87 132 90 135 
rect 87 135 90 138 
rect 87 138 90 141 
rect 87 141 90 144 
rect 87 144 90 147 
rect 87 147 90 150 
rect 87 150 90 153 
rect 87 153 90 156 
rect 87 156 90 159 
rect 87 159 90 162 
rect 87 162 90 165 
rect 87 165 90 168 
rect 87 168 90 171 
rect 87 171 90 174 
rect 87 174 90 177 
rect 87 177 90 180 
rect 87 180 90 183 
rect 87 183 90 186 
rect 87 186 90 189 
rect 87 189 90 192 
rect 87 192 90 195 
rect 87 195 90 198 
rect 87 198 90 201 
rect 87 201 90 204 
rect 87 204 90 207 
rect 87 207 90 210 
rect 87 210 90 213 
rect 87 213 90 216 
rect 87 216 90 219 
rect 87 219 90 222 
rect 87 222 90 225 
rect 87 225 90 228 
rect 87 228 90 231 
rect 87 231 90 234 
rect 87 234 90 237 
rect 87 237 90 240 
rect 87 240 90 243 
rect 87 243 90 246 
rect 87 246 90 249 
rect 87 249 90 252 
rect 87 252 90 255 
rect 87 255 90 258 
rect 87 258 90 261 
rect 87 261 90 264 
rect 87 264 90 267 
rect 87 267 90 270 
rect 87 270 90 273 
rect 87 273 90 276 
rect 87 276 90 279 
rect 87 279 90 282 
rect 87 282 90 285 
rect 87 285 90 288 
rect 87 288 90 291 
rect 87 291 90 294 
rect 87 294 90 297 
rect 87 297 90 300 
rect 87 300 90 303 
rect 87 303 90 306 
rect 87 306 90 309 
rect 87 309 90 312 
rect 87 312 90 315 
rect 87 315 90 318 
rect 87 318 90 321 
rect 87 321 90 324 
rect 87 324 90 327 
rect 87 327 90 330 
rect 87 330 90 333 
rect 87 333 90 336 
rect 87 336 90 339 
rect 87 339 90 342 
rect 87 342 90 345 
rect 87 345 90 348 
rect 87 348 90 351 
rect 87 351 90 354 
rect 87 354 90 357 
rect 87 357 90 360 
rect 87 360 90 363 
rect 87 363 90 366 
rect 87 366 90 369 
rect 87 369 90 372 
rect 87 372 90 375 
rect 87 375 90 378 
rect 87 378 90 381 
rect 87 381 90 384 
rect 87 384 90 387 
rect 87 387 90 390 
rect 87 390 90 393 
rect 87 393 90 396 
rect 87 396 90 399 
rect 87 399 90 402 
rect 87 402 90 405 
rect 87 405 90 408 
rect 87 408 90 411 
rect 87 411 90 414 
rect 87 414 90 417 
rect 87 417 90 420 
rect 87 420 90 423 
rect 87 423 90 426 
rect 87 426 90 429 
rect 87 429 90 432 
rect 87 432 90 435 
rect 87 435 90 438 
rect 87 438 90 441 
rect 87 441 90 444 
rect 87 444 90 447 
rect 87 447 90 450 
rect 87 450 90 453 
rect 87 453 90 456 
rect 87 456 90 459 
rect 87 459 90 462 
rect 87 462 90 465 
rect 87 465 90 468 
rect 87 468 90 471 
rect 87 471 90 474 
rect 87 474 90 477 
rect 87 477 90 480 
rect 87 480 90 483 
rect 87 483 90 486 
rect 87 486 90 489 
rect 87 489 90 492 
rect 87 492 90 495 
rect 87 495 90 498 
rect 87 498 90 501 
rect 87 501 90 504 
rect 87 504 90 507 
rect 87 507 90 510 
rect 90 0 93 3 
rect 90 3 93 6 
rect 90 6 93 9 
rect 90 9 93 12 
rect 90 12 93 15 
rect 90 15 93 18 
rect 90 18 93 21 
rect 90 21 93 24 
rect 90 24 93 27 
rect 90 27 93 30 
rect 90 30 93 33 
rect 90 33 93 36 
rect 90 36 93 39 
rect 90 39 93 42 
rect 90 42 93 45 
rect 90 45 93 48 
rect 90 48 93 51 
rect 90 51 93 54 
rect 90 54 93 57 
rect 90 57 93 60 
rect 90 60 93 63 
rect 90 63 93 66 
rect 90 66 93 69 
rect 90 69 93 72 
rect 90 72 93 75 
rect 90 75 93 78 
rect 90 78 93 81 
rect 90 81 93 84 
rect 90 84 93 87 
rect 90 87 93 90 
rect 90 90 93 93 
rect 90 93 93 96 
rect 90 96 93 99 
rect 90 99 93 102 
rect 90 102 93 105 
rect 90 105 93 108 
rect 90 108 93 111 
rect 90 111 93 114 
rect 90 114 93 117 
rect 90 117 93 120 
rect 90 120 93 123 
rect 90 123 93 126 
rect 90 126 93 129 
rect 90 129 93 132 
rect 90 132 93 135 
rect 90 135 93 138 
rect 90 138 93 141 
rect 90 141 93 144 
rect 90 144 93 147 
rect 90 147 93 150 
rect 90 150 93 153 
rect 90 153 93 156 
rect 90 156 93 159 
rect 90 159 93 162 
rect 90 162 93 165 
rect 90 165 93 168 
rect 90 168 93 171 
rect 90 171 93 174 
rect 90 174 93 177 
rect 90 177 93 180 
rect 90 180 93 183 
rect 90 183 93 186 
rect 90 186 93 189 
rect 90 189 93 192 
rect 90 192 93 195 
rect 90 195 93 198 
rect 90 198 93 201 
rect 90 201 93 204 
rect 90 204 93 207 
rect 90 207 93 210 
rect 90 210 93 213 
rect 90 213 93 216 
rect 90 216 93 219 
rect 90 219 93 222 
rect 90 222 93 225 
rect 90 225 93 228 
rect 90 228 93 231 
rect 90 231 93 234 
rect 90 234 93 237 
rect 90 237 93 240 
rect 90 240 93 243 
rect 90 243 93 246 
rect 90 246 93 249 
rect 90 249 93 252 
rect 90 252 93 255 
rect 90 255 93 258 
rect 90 258 93 261 
rect 90 261 93 264 
rect 90 264 93 267 
rect 90 267 93 270 
rect 90 270 93 273 
rect 90 273 93 276 
rect 90 276 93 279 
rect 90 279 93 282 
rect 90 282 93 285 
rect 90 285 93 288 
rect 90 288 93 291 
rect 90 291 93 294 
rect 90 294 93 297 
rect 90 297 93 300 
rect 90 300 93 303 
rect 90 303 93 306 
rect 90 306 93 309 
rect 90 309 93 312 
rect 90 312 93 315 
rect 90 315 93 318 
rect 90 318 93 321 
rect 90 321 93 324 
rect 90 324 93 327 
rect 90 327 93 330 
rect 90 330 93 333 
rect 90 333 93 336 
rect 90 336 93 339 
rect 90 339 93 342 
rect 90 342 93 345 
rect 90 345 93 348 
rect 90 348 93 351 
rect 90 351 93 354 
rect 90 354 93 357 
rect 90 357 93 360 
rect 90 360 93 363 
rect 90 363 93 366 
rect 90 366 93 369 
rect 90 369 93 372 
rect 90 372 93 375 
rect 90 375 93 378 
rect 90 378 93 381 
rect 90 381 93 384 
rect 90 384 93 387 
rect 90 387 93 390 
rect 90 390 93 393 
rect 90 393 93 396 
rect 90 396 93 399 
rect 90 399 93 402 
rect 90 402 93 405 
rect 90 405 93 408 
rect 90 408 93 411 
rect 90 411 93 414 
rect 90 414 93 417 
rect 90 417 93 420 
rect 90 420 93 423 
rect 90 423 93 426 
rect 90 426 93 429 
rect 90 429 93 432 
rect 90 432 93 435 
rect 90 435 93 438 
rect 90 438 93 441 
rect 90 441 93 444 
rect 90 444 93 447 
rect 90 447 93 450 
rect 90 450 93 453 
rect 90 453 93 456 
rect 90 456 93 459 
rect 90 459 93 462 
rect 90 462 93 465 
rect 90 465 93 468 
rect 90 468 93 471 
rect 90 471 93 474 
rect 90 474 93 477 
rect 90 477 93 480 
rect 90 480 93 483 
rect 90 483 93 486 
rect 90 486 93 489 
rect 90 489 93 492 
rect 90 492 93 495 
rect 90 495 93 498 
rect 90 498 93 501 
rect 90 501 93 504 
rect 90 504 93 507 
rect 90 507 93 510 
rect 93 0 96 3 
rect 93 3 96 6 
rect 93 6 96 9 
rect 93 9 96 12 
rect 93 12 96 15 
rect 93 15 96 18 
rect 93 18 96 21 
rect 93 21 96 24 
rect 93 24 96 27 
rect 93 27 96 30 
rect 93 30 96 33 
rect 93 33 96 36 
rect 93 36 96 39 
rect 93 39 96 42 
rect 93 42 96 45 
rect 93 45 96 48 
rect 93 48 96 51 
rect 93 51 96 54 
rect 93 54 96 57 
rect 93 57 96 60 
rect 93 60 96 63 
rect 93 63 96 66 
rect 93 66 96 69 
rect 93 69 96 72 
rect 93 72 96 75 
rect 93 75 96 78 
rect 93 78 96 81 
rect 93 81 96 84 
rect 93 84 96 87 
rect 93 87 96 90 
rect 93 90 96 93 
rect 93 93 96 96 
rect 93 96 96 99 
rect 93 99 96 102 
rect 93 102 96 105 
rect 93 105 96 108 
rect 93 108 96 111 
rect 93 111 96 114 
rect 93 114 96 117 
rect 93 117 96 120 
rect 93 120 96 123 
rect 93 123 96 126 
rect 93 126 96 129 
rect 93 129 96 132 
rect 93 132 96 135 
rect 93 135 96 138 
rect 93 138 96 141 
rect 93 141 96 144 
rect 93 144 96 147 
rect 93 147 96 150 
rect 93 150 96 153 
rect 93 153 96 156 
rect 93 156 96 159 
rect 93 159 96 162 
rect 93 162 96 165 
rect 93 165 96 168 
rect 93 168 96 171 
rect 93 171 96 174 
rect 93 174 96 177 
rect 93 177 96 180 
rect 93 180 96 183 
rect 93 183 96 186 
rect 93 186 96 189 
rect 93 189 96 192 
rect 93 192 96 195 
rect 93 195 96 198 
rect 93 198 96 201 
rect 93 201 96 204 
rect 93 204 96 207 
rect 93 207 96 210 
rect 93 210 96 213 
rect 93 213 96 216 
rect 93 216 96 219 
rect 93 219 96 222 
rect 93 222 96 225 
rect 93 225 96 228 
rect 93 228 96 231 
rect 93 231 96 234 
rect 93 234 96 237 
rect 93 237 96 240 
rect 93 240 96 243 
rect 93 243 96 246 
rect 93 246 96 249 
rect 93 249 96 252 
rect 93 252 96 255 
rect 93 255 96 258 
rect 93 258 96 261 
rect 93 261 96 264 
rect 93 264 96 267 
rect 93 267 96 270 
rect 93 270 96 273 
rect 93 273 96 276 
rect 93 276 96 279 
rect 93 279 96 282 
rect 93 282 96 285 
rect 93 285 96 288 
rect 93 288 96 291 
rect 93 291 96 294 
rect 93 294 96 297 
rect 93 297 96 300 
rect 93 300 96 303 
rect 93 303 96 306 
rect 93 306 96 309 
rect 93 309 96 312 
rect 93 312 96 315 
rect 93 315 96 318 
rect 93 318 96 321 
rect 93 321 96 324 
rect 93 324 96 327 
rect 93 327 96 330 
rect 93 330 96 333 
rect 93 333 96 336 
rect 93 336 96 339 
rect 93 339 96 342 
rect 93 342 96 345 
rect 93 345 96 348 
rect 93 348 96 351 
rect 93 351 96 354 
rect 93 354 96 357 
rect 93 357 96 360 
rect 93 360 96 363 
rect 93 363 96 366 
rect 93 366 96 369 
rect 93 369 96 372 
rect 93 372 96 375 
rect 93 375 96 378 
rect 93 378 96 381 
rect 93 381 96 384 
rect 93 384 96 387 
rect 93 387 96 390 
rect 93 390 96 393 
rect 93 393 96 396 
rect 93 396 96 399 
rect 93 399 96 402 
rect 93 402 96 405 
rect 93 405 96 408 
rect 93 408 96 411 
rect 93 411 96 414 
rect 93 414 96 417 
rect 93 417 96 420 
rect 93 420 96 423 
rect 93 423 96 426 
rect 93 426 96 429 
rect 93 429 96 432 
rect 93 432 96 435 
rect 93 435 96 438 
rect 93 438 96 441 
rect 93 441 96 444 
rect 93 444 96 447 
rect 93 447 96 450 
rect 93 450 96 453 
rect 93 453 96 456 
rect 93 456 96 459 
rect 93 459 96 462 
rect 93 462 96 465 
rect 93 465 96 468 
rect 93 468 96 471 
rect 93 471 96 474 
rect 93 474 96 477 
rect 93 477 96 480 
rect 93 480 96 483 
rect 93 483 96 486 
rect 93 486 96 489 
rect 93 489 96 492 
rect 93 492 96 495 
rect 93 495 96 498 
rect 93 498 96 501 
rect 93 501 96 504 
rect 93 504 96 507 
rect 93 507 96 510 
rect 96 0 99 3 
rect 96 3 99 6 
rect 96 6 99 9 
rect 96 9 99 12 
rect 96 12 99 15 
rect 96 15 99 18 
rect 96 18 99 21 
rect 96 21 99 24 
rect 96 24 99 27 
rect 96 27 99 30 
rect 96 30 99 33 
rect 96 33 99 36 
rect 96 36 99 39 
rect 96 39 99 42 
rect 96 42 99 45 
rect 96 45 99 48 
rect 96 48 99 51 
rect 96 51 99 54 
rect 96 54 99 57 
rect 96 57 99 60 
rect 96 60 99 63 
rect 96 63 99 66 
rect 96 66 99 69 
rect 96 69 99 72 
rect 96 72 99 75 
rect 96 75 99 78 
rect 96 78 99 81 
rect 96 81 99 84 
rect 96 84 99 87 
rect 96 87 99 90 
rect 96 90 99 93 
rect 96 93 99 96 
rect 96 96 99 99 
rect 96 99 99 102 
rect 96 102 99 105 
rect 96 105 99 108 
rect 96 108 99 111 
rect 96 111 99 114 
rect 96 114 99 117 
rect 96 117 99 120 
rect 96 120 99 123 
rect 96 123 99 126 
rect 96 126 99 129 
rect 96 129 99 132 
rect 96 132 99 135 
rect 96 135 99 138 
rect 96 138 99 141 
rect 96 141 99 144 
rect 96 144 99 147 
rect 96 147 99 150 
rect 96 150 99 153 
rect 96 153 99 156 
rect 96 156 99 159 
rect 96 159 99 162 
rect 96 162 99 165 
rect 96 165 99 168 
rect 96 168 99 171 
rect 96 171 99 174 
rect 96 174 99 177 
rect 96 177 99 180 
rect 96 180 99 183 
rect 96 183 99 186 
rect 96 186 99 189 
rect 96 189 99 192 
rect 96 192 99 195 
rect 96 195 99 198 
rect 96 198 99 201 
rect 96 201 99 204 
rect 96 204 99 207 
rect 96 207 99 210 
rect 96 210 99 213 
rect 96 213 99 216 
rect 96 216 99 219 
rect 96 219 99 222 
rect 96 222 99 225 
rect 96 225 99 228 
rect 96 228 99 231 
rect 96 231 99 234 
rect 96 234 99 237 
rect 96 237 99 240 
rect 96 240 99 243 
rect 96 243 99 246 
rect 96 246 99 249 
rect 96 249 99 252 
rect 96 252 99 255 
rect 96 255 99 258 
rect 96 258 99 261 
rect 96 261 99 264 
rect 96 264 99 267 
rect 96 267 99 270 
rect 96 270 99 273 
rect 96 273 99 276 
rect 96 276 99 279 
rect 96 279 99 282 
rect 96 282 99 285 
rect 96 285 99 288 
rect 96 288 99 291 
rect 96 291 99 294 
rect 96 294 99 297 
rect 96 297 99 300 
rect 96 300 99 303 
rect 96 303 99 306 
rect 96 306 99 309 
rect 96 309 99 312 
rect 96 312 99 315 
rect 96 315 99 318 
rect 96 318 99 321 
rect 96 321 99 324 
rect 96 324 99 327 
rect 96 327 99 330 
rect 96 330 99 333 
rect 96 333 99 336 
rect 96 336 99 339 
rect 96 339 99 342 
rect 96 342 99 345 
rect 96 345 99 348 
rect 96 348 99 351 
rect 96 351 99 354 
rect 96 354 99 357 
rect 96 357 99 360 
rect 96 360 99 363 
rect 96 363 99 366 
rect 96 366 99 369 
rect 96 369 99 372 
rect 96 372 99 375 
rect 96 375 99 378 
rect 96 378 99 381 
rect 96 381 99 384 
rect 96 384 99 387 
rect 96 387 99 390 
rect 96 390 99 393 
rect 96 393 99 396 
rect 96 396 99 399 
rect 96 399 99 402 
rect 96 402 99 405 
rect 96 405 99 408 
rect 96 408 99 411 
rect 96 411 99 414 
rect 96 414 99 417 
rect 96 417 99 420 
rect 96 420 99 423 
rect 96 423 99 426 
rect 96 426 99 429 
rect 96 429 99 432 
rect 96 432 99 435 
rect 96 435 99 438 
rect 96 438 99 441 
rect 96 441 99 444 
rect 96 444 99 447 
rect 96 447 99 450 
rect 96 450 99 453 
rect 96 453 99 456 
rect 96 456 99 459 
rect 96 459 99 462 
rect 96 462 99 465 
rect 96 465 99 468 
rect 96 468 99 471 
rect 96 471 99 474 
rect 96 474 99 477 
rect 96 477 99 480 
rect 96 480 99 483 
rect 96 483 99 486 
rect 96 486 99 489 
rect 96 489 99 492 
rect 96 492 99 495 
rect 96 495 99 498 
rect 96 498 99 501 
rect 96 501 99 504 
rect 96 504 99 507 
rect 96 507 99 510 
rect 99 0 102 3 
rect 99 3 102 6 
rect 99 6 102 9 
rect 99 9 102 12 
rect 99 12 102 15 
rect 99 15 102 18 
rect 99 18 102 21 
rect 99 21 102 24 
rect 99 24 102 27 
rect 99 27 102 30 
rect 99 30 102 33 
rect 99 33 102 36 
rect 99 36 102 39 
rect 99 39 102 42 
rect 99 42 102 45 
rect 99 45 102 48 
rect 99 48 102 51 
rect 99 51 102 54 
rect 99 54 102 57 
rect 99 57 102 60 
rect 99 60 102 63 
rect 99 63 102 66 
rect 99 66 102 69 
rect 99 69 102 72 
rect 99 72 102 75 
rect 99 75 102 78 
rect 99 78 102 81 
rect 99 81 102 84 
rect 99 84 102 87 
rect 99 87 102 90 
rect 99 90 102 93 
rect 99 93 102 96 
rect 99 96 102 99 
rect 99 99 102 102 
rect 99 102 102 105 
rect 99 105 102 108 
rect 99 108 102 111 
rect 99 111 102 114 
rect 99 114 102 117 
rect 99 117 102 120 
rect 99 120 102 123 
rect 99 123 102 126 
rect 99 126 102 129 
rect 99 129 102 132 
rect 99 132 102 135 
rect 99 135 102 138 
rect 99 138 102 141 
rect 99 141 102 144 
rect 99 144 102 147 
rect 99 147 102 150 
rect 99 150 102 153 
rect 99 153 102 156 
rect 99 156 102 159 
rect 99 159 102 162 
rect 99 162 102 165 
rect 99 165 102 168 
rect 99 168 102 171 
rect 99 171 102 174 
rect 99 174 102 177 
rect 99 177 102 180 
rect 99 180 102 183 
rect 99 183 102 186 
rect 99 186 102 189 
rect 99 189 102 192 
rect 99 192 102 195 
rect 99 195 102 198 
rect 99 198 102 201 
rect 99 201 102 204 
rect 99 204 102 207 
rect 99 207 102 210 
rect 99 210 102 213 
rect 99 213 102 216 
rect 99 216 102 219 
rect 99 219 102 222 
rect 99 222 102 225 
rect 99 225 102 228 
rect 99 228 102 231 
rect 99 231 102 234 
rect 99 234 102 237 
rect 99 237 102 240 
rect 99 240 102 243 
rect 99 243 102 246 
rect 99 246 102 249 
rect 99 249 102 252 
rect 99 252 102 255 
rect 99 255 102 258 
rect 99 258 102 261 
rect 99 261 102 264 
rect 99 264 102 267 
rect 99 267 102 270 
rect 99 270 102 273 
rect 99 273 102 276 
rect 99 276 102 279 
rect 99 279 102 282 
rect 99 282 102 285 
rect 99 285 102 288 
rect 99 288 102 291 
rect 99 291 102 294 
rect 99 294 102 297 
rect 99 297 102 300 
rect 99 300 102 303 
rect 99 303 102 306 
rect 99 306 102 309 
rect 99 309 102 312 
rect 99 312 102 315 
rect 99 315 102 318 
rect 99 318 102 321 
rect 99 321 102 324 
rect 99 324 102 327 
rect 99 327 102 330 
rect 99 330 102 333 
rect 99 333 102 336 
rect 99 336 102 339 
rect 99 339 102 342 
rect 99 342 102 345 
rect 99 345 102 348 
rect 99 348 102 351 
rect 99 351 102 354 
rect 99 354 102 357 
rect 99 357 102 360 
rect 99 360 102 363 
rect 99 363 102 366 
rect 99 366 102 369 
rect 99 369 102 372 
rect 99 372 102 375 
rect 99 375 102 378 
rect 99 378 102 381 
rect 99 381 102 384 
rect 99 384 102 387 
rect 99 387 102 390 
rect 99 390 102 393 
rect 99 393 102 396 
rect 99 396 102 399 
rect 99 399 102 402 
rect 99 402 102 405 
rect 99 405 102 408 
rect 99 408 102 411 
rect 99 411 102 414 
rect 99 414 102 417 
rect 99 417 102 420 
rect 99 420 102 423 
rect 99 423 102 426 
rect 99 426 102 429 
rect 99 429 102 432 
rect 99 432 102 435 
rect 99 435 102 438 
rect 99 438 102 441 
rect 99 441 102 444 
rect 99 444 102 447 
rect 99 447 102 450 
rect 99 450 102 453 
rect 99 453 102 456 
rect 99 456 102 459 
rect 99 459 102 462 
rect 99 462 102 465 
rect 99 465 102 468 
rect 99 468 102 471 
rect 99 471 102 474 
rect 99 474 102 477 
rect 99 477 102 480 
rect 99 480 102 483 
rect 99 483 102 486 
rect 99 486 102 489 
rect 99 489 102 492 
rect 99 492 102 495 
rect 99 495 102 498 
rect 99 498 102 501 
rect 99 501 102 504 
rect 99 504 102 507 
rect 99 507 102 510 
rect 102 0 105 3 
rect 102 3 105 6 
rect 102 6 105 9 
rect 102 9 105 12 
rect 102 12 105 15 
rect 102 15 105 18 
rect 102 18 105 21 
rect 102 21 105 24 
rect 102 24 105 27 
rect 102 27 105 30 
rect 102 30 105 33 
rect 102 33 105 36 
rect 102 36 105 39 
rect 102 39 105 42 
rect 102 42 105 45 
rect 102 45 105 48 
rect 102 48 105 51 
rect 102 51 105 54 
rect 102 54 105 57 
rect 102 57 105 60 
rect 102 60 105 63 
rect 102 63 105 66 
rect 102 66 105 69 
rect 102 69 105 72 
rect 102 72 105 75 
rect 102 75 105 78 
rect 102 78 105 81 
rect 102 81 105 84 
rect 102 84 105 87 
rect 102 87 105 90 
rect 102 90 105 93 
rect 102 93 105 96 
rect 102 96 105 99 
rect 102 99 105 102 
rect 102 102 105 105 
rect 102 105 105 108 
rect 102 108 105 111 
rect 102 111 105 114 
rect 102 114 105 117 
rect 102 117 105 120 
rect 102 120 105 123 
rect 102 123 105 126 
rect 102 126 105 129 
rect 102 129 105 132 
rect 102 132 105 135 
rect 102 135 105 138 
rect 102 138 105 141 
rect 102 141 105 144 
rect 102 144 105 147 
rect 102 147 105 150 
rect 102 150 105 153 
rect 102 153 105 156 
rect 102 156 105 159 
rect 102 159 105 162 
rect 102 162 105 165 
rect 102 165 105 168 
rect 102 168 105 171 
rect 102 171 105 174 
rect 102 174 105 177 
rect 102 177 105 180 
rect 102 180 105 183 
rect 102 183 105 186 
rect 102 186 105 189 
rect 102 189 105 192 
rect 102 192 105 195 
rect 102 195 105 198 
rect 102 198 105 201 
rect 102 201 105 204 
rect 102 204 105 207 
rect 102 207 105 210 
rect 102 210 105 213 
rect 102 213 105 216 
rect 102 216 105 219 
rect 102 219 105 222 
rect 102 222 105 225 
rect 102 225 105 228 
rect 102 228 105 231 
rect 102 231 105 234 
rect 102 234 105 237 
rect 102 237 105 240 
rect 102 240 105 243 
rect 102 243 105 246 
rect 102 246 105 249 
rect 102 249 105 252 
rect 102 252 105 255 
rect 102 255 105 258 
rect 102 258 105 261 
rect 102 261 105 264 
rect 102 264 105 267 
rect 102 267 105 270 
rect 102 270 105 273 
rect 102 273 105 276 
rect 102 276 105 279 
rect 102 279 105 282 
rect 102 282 105 285 
rect 102 285 105 288 
rect 102 288 105 291 
rect 102 291 105 294 
rect 102 294 105 297 
rect 102 297 105 300 
rect 102 300 105 303 
rect 102 303 105 306 
rect 102 306 105 309 
rect 102 309 105 312 
rect 102 312 105 315 
rect 102 315 105 318 
rect 102 318 105 321 
rect 102 321 105 324 
rect 102 324 105 327 
rect 102 327 105 330 
rect 102 330 105 333 
rect 102 333 105 336 
rect 102 336 105 339 
rect 102 339 105 342 
rect 102 342 105 345 
rect 102 345 105 348 
rect 102 348 105 351 
rect 102 351 105 354 
rect 102 354 105 357 
rect 102 357 105 360 
rect 102 360 105 363 
rect 102 363 105 366 
rect 102 366 105 369 
rect 102 369 105 372 
rect 102 372 105 375 
rect 102 375 105 378 
rect 102 378 105 381 
rect 102 381 105 384 
rect 102 384 105 387 
rect 102 387 105 390 
rect 102 390 105 393 
rect 102 393 105 396 
rect 102 396 105 399 
rect 102 399 105 402 
rect 102 402 105 405 
rect 102 405 105 408 
rect 102 408 105 411 
rect 102 411 105 414 
rect 102 414 105 417 
rect 102 417 105 420 
rect 102 420 105 423 
rect 102 423 105 426 
rect 102 426 105 429 
rect 102 429 105 432 
rect 102 432 105 435 
rect 102 435 105 438 
rect 102 438 105 441 
rect 102 441 105 444 
rect 102 444 105 447 
rect 102 447 105 450 
rect 102 450 105 453 
rect 102 453 105 456 
rect 102 456 105 459 
rect 102 459 105 462 
rect 102 462 105 465 
rect 102 465 105 468 
rect 102 468 105 471 
rect 102 471 105 474 
rect 102 474 105 477 
rect 102 477 105 480 
rect 102 480 105 483 
rect 102 483 105 486 
rect 102 486 105 489 
rect 102 489 105 492 
rect 102 492 105 495 
rect 102 495 105 498 
rect 102 498 105 501 
rect 102 501 105 504 
rect 102 504 105 507 
rect 102 507 105 510 
rect 105 0 108 3 
rect 105 3 108 6 
rect 105 6 108 9 
rect 105 9 108 12 
rect 105 12 108 15 
rect 105 15 108 18 
rect 105 18 108 21 
rect 105 21 108 24 
rect 105 24 108 27 
rect 105 27 108 30 
rect 105 30 108 33 
rect 105 33 108 36 
rect 105 36 108 39 
rect 105 39 108 42 
rect 105 42 108 45 
rect 105 45 108 48 
rect 105 48 108 51 
rect 105 51 108 54 
rect 105 54 108 57 
rect 105 57 108 60 
rect 105 60 108 63 
rect 105 63 108 66 
rect 105 66 108 69 
rect 105 69 108 72 
rect 105 72 108 75 
rect 105 75 108 78 
rect 105 78 108 81 
rect 105 81 108 84 
rect 105 84 108 87 
rect 105 87 108 90 
rect 105 90 108 93 
rect 105 93 108 96 
rect 105 96 108 99 
rect 105 99 108 102 
rect 105 102 108 105 
rect 105 105 108 108 
rect 105 108 108 111 
rect 105 111 108 114 
rect 105 114 108 117 
rect 105 117 108 120 
rect 105 120 108 123 
rect 105 123 108 126 
rect 105 126 108 129 
rect 105 129 108 132 
rect 105 132 108 135 
rect 105 135 108 138 
rect 105 138 108 141 
rect 105 141 108 144 
rect 105 144 108 147 
rect 105 147 108 150 
rect 105 150 108 153 
rect 105 153 108 156 
rect 105 156 108 159 
rect 105 159 108 162 
rect 105 162 108 165 
rect 105 165 108 168 
rect 105 168 108 171 
rect 105 171 108 174 
rect 105 174 108 177 
rect 105 177 108 180 
rect 105 180 108 183 
rect 105 183 108 186 
rect 105 186 108 189 
rect 105 189 108 192 
rect 105 192 108 195 
rect 105 195 108 198 
rect 105 198 108 201 
rect 105 201 108 204 
rect 105 204 108 207 
rect 105 207 108 210 
rect 105 210 108 213 
rect 105 213 108 216 
rect 105 216 108 219 
rect 105 219 108 222 
rect 105 222 108 225 
rect 105 225 108 228 
rect 105 228 108 231 
rect 105 231 108 234 
rect 105 234 108 237 
rect 105 237 108 240 
rect 105 240 108 243 
rect 105 243 108 246 
rect 105 246 108 249 
rect 105 249 108 252 
rect 105 252 108 255 
rect 105 255 108 258 
rect 105 258 108 261 
rect 105 261 108 264 
rect 105 264 108 267 
rect 105 267 108 270 
rect 105 270 108 273 
rect 105 273 108 276 
rect 105 276 108 279 
rect 105 279 108 282 
rect 105 282 108 285 
rect 105 285 108 288 
rect 105 288 108 291 
rect 105 291 108 294 
rect 105 294 108 297 
rect 105 297 108 300 
rect 105 300 108 303 
rect 105 303 108 306 
rect 105 306 108 309 
rect 105 309 108 312 
rect 105 312 108 315 
rect 105 315 108 318 
rect 105 318 108 321 
rect 105 321 108 324 
rect 105 324 108 327 
rect 105 327 108 330 
rect 105 330 108 333 
rect 105 333 108 336 
rect 105 336 108 339 
rect 105 339 108 342 
rect 105 342 108 345 
rect 105 345 108 348 
rect 105 348 108 351 
rect 105 351 108 354 
rect 105 354 108 357 
rect 105 357 108 360 
rect 105 360 108 363 
rect 105 363 108 366 
rect 105 366 108 369 
rect 105 369 108 372 
rect 105 372 108 375 
rect 105 375 108 378 
rect 105 378 108 381 
rect 105 381 108 384 
rect 105 384 108 387 
rect 105 387 108 390 
rect 105 390 108 393 
rect 105 393 108 396 
rect 105 396 108 399 
rect 105 399 108 402 
rect 105 402 108 405 
rect 105 405 108 408 
rect 105 408 108 411 
rect 105 411 108 414 
rect 105 414 108 417 
rect 105 417 108 420 
rect 105 420 108 423 
rect 105 423 108 426 
rect 105 426 108 429 
rect 105 429 108 432 
rect 105 432 108 435 
rect 105 435 108 438 
rect 105 438 108 441 
rect 105 441 108 444 
rect 105 444 108 447 
rect 105 447 108 450 
rect 105 450 108 453 
rect 105 453 108 456 
rect 105 456 108 459 
rect 105 459 108 462 
rect 105 462 108 465 
rect 105 465 108 468 
rect 105 468 108 471 
rect 105 471 108 474 
rect 105 474 108 477 
rect 105 477 108 480 
rect 105 480 108 483 
rect 105 483 108 486 
rect 105 486 108 489 
rect 105 489 108 492 
rect 105 492 108 495 
rect 105 495 108 498 
rect 105 498 108 501 
rect 105 501 108 504 
rect 105 504 108 507 
rect 105 507 108 510 
rect 108 0 111 3 
rect 108 3 111 6 
rect 108 6 111 9 
rect 108 9 111 12 
rect 108 12 111 15 
rect 108 15 111 18 
rect 108 18 111 21 
rect 108 21 111 24 
rect 108 24 111 27 
rect 108 27 111 30 
rect 108 30 111 33 
rect 108 33 111 36 
rect 108 36 111 39 
rect 108 39 111 42 
rect 108 42 111 45 
rect 108 45 111 48 
rect 108 48 111 51 
rect 108 51 111 54 
rect 108 54 111 57 
rect 108 57 111 60 
rect 108 60 111 63 
rect 108 63 111 66 
rect 108 66 111 69 
rect 108 69 111 72 
rect 108 72 111 75 
rect 108 75 111 78 
rect 108 78 111 81 
rect 108 81 111 84 
rect 108 84 111 87 
rect 108 87 111 90 
rect 108 90 111 93 
rect 108 93 111 96 
rect 108 96 111 99 
rect 108 99 111 102 
rect 108 102 111 105 
rect 108 105 111 108 
rect 108 108 111 111 
rect 108 111 111 114 
rect 108 114 111 117 
rect 108 117 111 120 
rect 108 120 111 123 
rect 108 123 111 126 
rect 108 126 111 129 
rect 108 129 111 132 
rect 108 132 111 135 
rect 108 135 111 138 
rect 108 138 111 141 
rect 108 141 111 144 
rect 108 144 111 147 
rect 108 147 111 150 
rect 108 150 111 153 
rect 108 153 111 156 
rect 108 156 111 159 
rect 108 159 111 162 
rect 108 162 111 165 
rect 108 165 111 168 
rect 108 168 111 171 
rect 108 171 111 174 
rect 108 174 111 177 
rect 108 177 111 180 
rect 108 180 111 183 
rect 108 183 111 186 
rect 108 186 111 189 
rect 108 189 111 192 
rect 108 192 111 195 
rect 108 195 111 198 
rect 108 198 111 201 
rect 108 201 111 204 
rect 108 204 111 207 
rect 108 207 111 210 
rect 108 210 111 213 
rect 108 213 111 216 
rect 108 216 111 219 
rect 108 219 111 222 
rect 108 222 111 225 
rect 108 225 111 228 
rect 108 228 111 231 
rect 108 231 111 234 
rect 108 234 111 237 
rect 108 237 111 240 
rect 108 240 111 243 
rect 108 243 111 246 
rect 108 246 111 249 
rect 108 249 111 252 
rect 108 252 111 255 
rect 108 255 111 258 
rect 108 258 111 261 
rect 108 261 111 264 
rect 108 264 111 267 
rect 108 267 111 270 
rect 108 270 111 273 
rect 108 273 111 276 
rect 108 276 111 279 
rect 108 279 111 282 
rect 108 282 111 285 
rect 108 285 111 288 
rect 108 288 111 291 
rect 108 291 111 294 
rect 108 294 111 297 
rect 108 297 111 300 
rect 108 300 111 303 
rect 108 303 111 306 
rect 108 306 111 309 
rect 108 309 111 312 
rect 108 312 111 315 
rect 108 315 111 318 
rect 108 318 111 321 
rect 108 321 111 324 
rect 108 324 111 327 
rect 108 327 111 330 
rect 108 330 111 333 
rect 108 333 111 336 
rect 108 336 111 339 
rect 108 339 111 342 
rect 108 342 111 345 
rect 108 345 111 348 
rect 108 348 111 351 
rect 108 351 111 354 
rect 108 354 111 357 
rect 108 357 111 360 
rect 108 360 111 363 
rect 108 363 111 366 
rect 108 366 111 369 
rect 108 369 111 372 
rect 108 372 111 375 
rect 108 375 111 378 
rect 108 378 111 381 
rect 108 381 111 384 
rect 108 384 111 387 
rect 108 387 111 390 
rect 108 390 111 393 
rect 108 393 111 396 
rect 108 396 111 399 
rect 108 399 111 402 
rect 108 402 111 405 
rect 108 405 111 408 
rect 108 408 111 411 
rect 108 411 111 414 
rect 108 414 111 417 
rect 108 417 111 420 
rect 108 420 111 423 
rect 108 423 111 426 
rect 108 426 111 429 
rect 108 429 111 432 
rect 108 432 111 435 
rect 108 435 111 438 
rect 108 438 111 441 
rect 108 441 111 444 
rect 108 444 111 447 
rect 108 447 111 450 
rect 108 450 111 453 
rect 108 453 111 456 
rect 108 456 111 459 
rect 108 459 111 462 
rect 108 462 111 465 
rect 108 465 111 468 
rect 108 468 111 471 
rect 108 471 111 474 
rect 108 474 111 477 
rect 108 477 111 480 
rect 108 480 111 483 
rect 108 483 111 486 
rect 108 486 111 489 
rect 108 489 111 492 
rect 108 492 111 495 
rect 108 495 111 498 
rect 108 498 111 501 
rect 108 501 111 504 
rect 108 504 111 507 
rect 108 507 111 510 
rect 111 0 114 3 
rect 111 3 114 6 
rect 111 6 114 9 
rect 111 9 114 12 
rect 111 12 114 15 
rect 111 15 114 18 
rect 111 18 114 21 
rect 111 21 114 24 
rect 111 24 114 27 
rect 111 27 114 30 
rect 111 30 114 33 
rect 111 33 114 36 
rect 111 36 114 39 
rect 111 39 114 42 
rect 111 42 114 45 
rect 111 45 114 48 
rect 111 48 114 51 
rect 111 51 114 54 
rect 111 54 114 57 
rect 111 57 114 60 
rect 111 60 114 63 
rect 111 63 114 66 
rect 111 66 114 69 
rect 111 69 114 72 
rect 111 72 114 75 
rect 111 75 114 78 
rect 111 78 114 81 
rect 111 81 114 84 
rect 111 84 114 87 
rect 111 87 114 90 
rect 111 90 114 93 
rect 111 93 114 96 
rect 111 96 114 99 
rect 111 99 114 102 
rect 111 102 114 105 
rect 111 105 114 108 
rect 111 108 114 111 
rect 111 111 114 114 
rect 111 114 114 117 
rect 111 117 114 120 
rect 111 120 114 123 
rect 111 123 114 126 
rect 111 126 114 129 
rect 111 129 114 132 
rect 111 132 114 135 
rect 111 135 114 138 
rect 111 138 114 141 
rect 111 141 114 144 
rect 111 144 114 147 
rect 111 147 114 150 
rect 111 150 114 153 
rect 111 153 114 156 
rect 111 156 114 159 
rect 111 159 114 162 
rect 111 162 114 165 
rect 111 165 114 168 
rect 111 168 114 171 
rect 111 171 114 174 
rect 111 174 114 177 
rect 111 177 114 180 
rect 111 180 114 183 
rect 111 183 114 186 
rect 111 186 114 189 
rect 111 189 114 192 
rect 111 192 114 195 
rect 111 195 114 198 
rect 111 198 114 201 
rect 111 201 114 204 
rect 111 204 114 207 
rect 111 207 114 210 
rect 111 210 114 213 
rect 111 213 114 216 
rect 111 216 114 219 
rect 111 219 114 222 
rect 111 222 114 225 
rect 111 225 114 228 
rect 111 228 114 231 
rect 111 231 114 234 
rect 111 234 114 237 
rect 111 237 114 240 
rect 111 240 114 243 
rect 111 243 114 246 
rect 111 246 114 249 
rect 111 249 114 252 
rect 111 252 114 255 
rect 111 255 114 258 
rect 111 258 114 261 
rect 111 261 114 264 
rect 111 264 114 267 
rect 111 267 114 270 
rect 111 270 114 273 
rect 111 273 114 276 
rect 111 276 114 279 
rect 111 279 114 282 
rect 111 282 114 285 
rect 111 285 114 288 
rect 111 288 114 291 
rect 111 291 114 294 
rect 111 294 114 297 
rect 111 297 114 300 
rect 111 300 114 303 
rect 111 303 114 306 
rect 111 306 114 309 
rect 111 309 114 312 
rect 111 312 114 315 
rect 111 315 114 318 
rect 111 318 114 321 
rect 111 321 114 324 
rect 111 324 114 327 
rect 111 327 114 330 
rect 111 330 114 333 
rect 111 333 114 336 
rect 111 336 114 339 
rect 111 339 114 342 
rect 111 342 114 345 
rect 111 345 114 348 
rect 111 348 114 351 
rect 111 351 114 354 
rect 111 354 114 357 
rect 111 357 114 360 
rect 111 360 114 363 
rect 111 363 114 366 
rect 111 366 114 369 
rect 111 369 114 372 
rect 111 372 114 375 
rect 111 375 114 378 
rect 111 378 114 381 
rect 111 381 114 384 
rect 111 384 114 387 
rect 111 387 114 390 
rect 111 390 114 393 
rect 111 393 114 396 
rect 111 396 114 399 
rect 111 399 114 402 
rect 111 402 114 405 
rect 111 405 114 408 
rect 111 408 114 411 
rect 111 411 114 414 
rect 111 414 114 417 
rect 111 417 114 420 
rect 111 420 114 423 
rect 111 423 114 426 
rect 111 426 114 429 
rect 111 429 114 432 
rect 111 432 114 435 
rect 111 435 114 438 
rect 111 438 114 441 
rect 111 441 114 444 
rect 111 444 114 447 
rect 111 447 114 450 
rect 111 450 114 453 
rect 111 453 114 456 
rect 111 456 114 459 
rect 111 459 114 462 
rect 111 462 114 465 
rect 111 465 114 468 
rect 111 468 114 471 
rect 111 471 114 474 
rect 111 474 114 477 
rect 111 477 114 480 
rect 111 480 114 483 
rect 111 483 114 486 
rect 111 486 114 489 
rect 111 489 114 492 
rect 111 492 114 495 
rect 111 495 114 498 
rect 111 498 114 501 
rect 111 501 114 504 
rect 111 504 114 507 
rect 111 507 114 510 
rect 114 0 117 3 
rect 114 3 117 6 
rect 114 6 117 9 
rect 114 9 117 12 
rect 114 12 117 15 
rect 114 15 117 18 
rect 114 18 117 21 
rect 114 21 117 24 
rect 114 24 117 27 
rect 114 27 117 30 
rect 114 30 117 33 
rect 114 33 117 36 
rect 114 36 117 39 
rect 114 39 117 42 
rect 114 42 117 45 
rect 114 45 117 48 
rect 114 48 117 51 
rect 114 51 117 54 
rect 114 54 117 57 
rect 114 57 117 60 
rect 114 60 117 63 
rect 114 63 117 66 
rect 114 66 117 69 
rect 114 69 117 72 
rect 114 72 117 75 
rect 114 75 117 78 
rect 114 78 117 81 
rect 114 81 117 84 
rect 114 84 117 87 
rect 114 87 117 90 
rect 114 90 117 93 
rect 114 93 117 96 
rect 114 96 117 99 
rect 114 99 117 102 
rect 114 102 117 105 
rect 114 105 117 108 
rect 114 108 117 111 
rect 114 111 117 114 
rect 114 114 117 117 
rect 114 117 117 120 
rect 114 120 117 123 
rect 114 123 117 126 
rect 114 126 117 129 
rect 114 129 117 132 
rect 114 132 117 135 
rect 114 135 117 138 
rect 114 138 117 141 
rect 114 141 117 144 
rect 114 144 117 147 
rect 114 147 117 150 
rect 114 150 117 153 
rect 114 153 117 156 
rect 114 156 117 159 
rect 114 159 117 162 
rect 114 162 117 165 
rect 114 165 117 168 
rect 114 168 117 171 
rect 114 171 117 174 
rect 114 174 117 177 
rect 114 177 117 180 
rect 114 180 117 183 
rect 114 183 117 186 
rect 114 186 117 189 
rect 114 189 117 192 
rect 114 192 117 195 
rect 114 195 117 198 
rect 114 198 117 201 
rect 114 201 117 204 
rect 114 204 117 207 
rect 114 207 117 210 
rect 114 210 117 213 
rect 114 213 117 216 
rect 114 216 117 219 
rect 114 219 117 222 
rect 114 222 117 225 
rect 114 225 117 228 
rect 114 228 117 231 
rect 114 231 117 234 
rect 114 234 117 237 
rect 114 237 117 240 
rect 114 240 117 243 
rect 114 243 117 246 
rect 114 246 117 249 
rect 114 249 117 252 
rect 114 252 117 255 
rect 114 255 117 258 
rect 114 258 117 261 
rect 114 261 117 264 
rect 114 264 117 267 
rect 114 267 117 270 
rect 114 270 117 273 
rect 114 273 117 276 
rect 114 276 117 279 
rect 114 279 117 282 
rect 114 282 117 285 
rect 114 285 117 288 
rect 114 288 117 291 
rect 114 291 117 294 
rect 114 294 117 297 
rect 114 297 117 300 
rect 114 300 117 303 
rect 114 303 117 306 
rect 114 306 117 309 
rect 114 309 117 312 
rect 114 312 117 315 
rect 114 315 117 318 
rect 114 318 117 321 
rect 114 321 117 324 
rect 114 324 117 327 
rect 114 327 117 330 
rect 114 330 117 333 
rect 114 333 117 336 
rect 114 336 117 339 
rect 114 339 117 342 
rect 114 342 117 345 
rect 114 345 117 348 
rect 114 348 117 351 
rect 114 351 117 354 
rect 114 354 117 357 
rect 114 357 117 360 
rect 114 360 117 363 
rect 114 363 117 366 
rect 114 366 117 369 
rect 114 369 117 372 
rect 114 372 117 375 
rect 114 375 117 378 
rect 114 378 117 381 
rect 114 381 117 384 
rect 114 384 117 387 
rect 114 387 117 390 
rect 114 390 117 393 
rect 114 393 117 396 
rect 114 396 117 399 
rect 114 399 117 402 
rect 114 402 117 405 
rect 114 405 117 408 
rect 114 408 117 411 
rect 114 411 117 414 
rect 114 414 117 417 
rect 114 417 117 420 
rect 114 420 117 423 
rect 114 423 117 426 
rect 114 426 117 429 
rect 114 429 117 432 
rect 114 432 117 435 
rect 114 435 117 438 
rect 114 438 117 441 
rect 114 441 117 444 
rect 114 444 117 447 
rect 114 447 117 450 
rect 114 450 117 453 
rect 114 453 117 456 
rect 114 456 117 459 
rect 114 459 117 462 
rect 114 462 117 465 
rect 114 465 117 468 
rect 114 468 117 471 
rect 114 471 117 474 
rect 114 474 117 477 
rect 114 477 117 480 
rect 114 480 117 483 
rect 114 483 117 486 
rect 114 486 117 489 
rect 114 489 117 492 
rect 114 492 117 495 
rect 114 495 117 498 
rect 114 498 117 501 
rect 114 501 117 504 
rect 114 504 117 507 
rect 114 507 117 510 
rect 117 0 120 3 
rect 117 3 120 6 
rect 117 6 120 9 
rect 117 9 120 12 
rect 117 12 120 15 
rect 117 15 120 18 
rect 117 18 120 21 
rect 117 21 120 24 
rect 117 24 120 27 
rect 117 27 120 30 
rect 117 30 120 33 
rect 117 33 120 36 
rect 117 36 120 39 
rect 117 39 120 42 
rect 117 42 120 45 
rect 117 45 120 48 
rect 117 48 120 51 
rect 117 51 120 54 
rect 117 54 120 57 
rect 117 57 120 60 
rect 117 60 120 63 
rect 117 63 120 66 
rect 117 66 120 69 
rect 117 69 120 72 
rect 117 72 120 75 
rect 117 75 120 78 
rect 117 78 120 81 
rect 117 81 120 84 
rect 117 84 120 87 
rect 117 87 120 90 
rect 117 90 120 93 
rect 117 93 120 96 
rect 117 96 120 99 
rect 117 99 120 102 
rect 117 102 120 105 
rect 117 105 120 108 
rect 117 108 120 111 
rect 117 111 120 114 
rect 117 114 120 117 
rect 117 117 120 120 
rect 117 120 120 123 
rect 117 123 120 126 
rect 117 126 120 129 
rect 117 129 120 132 
rect 117 132 120 135 
rect 117 135 120 138 
rect 117 138 120 141 
rect 117 141 120 144 
rect 117 144 120 147 
rect 117 147 120 150 
rect 117 150 120 153 
rect 117 153 120 156 
rect 117 156 120 159 
rect 117 159 120 162 
rect 117 162 120 165 
rect 117 165 120 168 
rect 117 168 120 171 
rect 117 171 120 174 
rect 117 174 120 177 
rect 117 177 120 180 
rect 117 180 120 183 
rect 117 183 120 186 
rect 117 186 120 189 
rect 117 189 120 192 
rect 117 192 120 195 
rect 117 195 120 198 
rect 117 198 120 201 
rect 117 201 120 204 
rect 117 204 120 207 
rect 117 207 120 210 
rect 117 210 120 213 
rect 117 213 120 216 
rect 117 216 120 219 
rect 117 219 120 222 
rect 117 222 120 225 
rect 117 225 120 228 
rect 117 228 120 231 
rect 117 231 120 234 
rect 117 234 120 237 
rect 117 237 120 240 
rect 117 240 120 243 
rect 117 243 120 246 
rect 117 246 120 249 
rect 117 249 120 252 
rect 117 252 120 255 
rect 117 255 120 258 
rect 117 258 120 261 
rect 117 261 120 264 
rect 117 264 120 267 
rect 117 267 120 270 
rect 117 270 120 273 
rect 117 273 120 276 
rect 117 276 120 279 
rect 117 279 120 282 
rect 117 282 120 285 
rect 117 285 120 288 
rect 117 288 120 291 
rect 117 291 120 294 
rect 117 294 120 297 
rect 117 297 120 300 
rect 117 300 120 303 
rect 117 303 120 306 
rect 117 306 120 309 
rect 117 309 120 312 
rect 117 312 120 315 
rect 117 315 120 318 
rect 117 318 120 321 
rect 117 321 120 324 
rect 117 324 120 327 
rect 117 327 120 330 
rect 117 330 120 333 
rect 117 333 120 336 
rect 117 336 120 339 
rect 117 339 120 342 
rect 117 342 120 345 
rect 117 345 120 348 
rect 117 348 120 351 
rect 117 351 120 354 
rect 117 354 120 357 
rect 117 357 120 360 
rect 117 360 120 363 
rect 117 363 120 366 
rect 117 366 120 369 
rect 117 369 120 372 
rect 117 372 120 375 
rect 117 375 120 378 
rect 117 378 120 381 
rect 117 381 120 384 
rect 117 384 120 387 
rect 117 387 120 390 
rect 117 390 120 393 
rect 117 393 120 396 
rect 117 396 120 399 
rect 117 399 120 402 
rect 117 402 120 405 
rect 117 405 120 408 
rect 117 408 120 411 
rect 117 411 120 414 
rect 117 414 120 417 
rect 117 417 120 420 
rect 117 420 120 423 
rect 117 423 120 426 
rect 117 426 120 429 
rect 117 429 120 432 
rect 117 432 120 435 
rect 117 435 120 438 
rect 117 438 120 441 
rect 117 441 120 444 
rect 117 444 120 447 
rect 117 447 120 450 
rect 117 450 120 453 
rect 117 453 120 456 
rect 117 456 120 459 
rect 117 459 120 462 
rect 117 462 120 465 
rect 117 465 120 468 
rect 117 468 120 471 
rect 117 471 120 474 
rect 117 474 120 477 
rect 117 477 120 480 
rect 117 480 120 483 
rect 117 483 120 486 
rect 117 486 120 489 
rect 117 489 120 492 
rect 117 492 120 495 
rect 117 495 120 498 
rect 117 498 120 501 
rect 117 501 120 504 
rect 117 504 120 507 
rect 117 507 120 510 
rect 120 0 123 3 
rect 120 3 123 6 
rect 120 6 123 9 
rect 120 9 123 12 
rect 120 12 123 15 
rect 120 15 123 18 
rect 120 18 123 21 
rect 120 21 123 24 
rect 120 24 123 27 
rect 120 27 123 30 
rect 120 30 123 33 
rect 120 33 123 36 
rect 120 36 123 39 
rect 120 39 123 42 
rect 120 42 123 45 
rect 120 45 123 48 
rect 120 48 123 51 
rect 120 51 123 54 
rect 120 54 123 57 
rect 120 57 123 60 
rect 120 60 123 63 
rect 120 63 123 66 
rect 120 66 123 69 
rect 120 69 123 72 
rect 120 72 123 75 
rect 120 75 123 78 
rect 120 78 123 81 
rect 120 81 123 84 
rect 120 84 123 87 
rect 120 87 123 90 
rect 120 90 123 93 
rect 120 93 123 96 
rect 120 96 123 99 
rect 120 99 123 102 
rect 120 102 123 105 
rect 120 105 123 108 
rect 120 108 123 111 
rect 120 111 123 114 
rect 120 114 123 117 
rect 120 117 123 120 
rect 120 120 123 123 
rect 120 123 123 126 
rect 120 126 123 129 
rect 120 129 123 132 
rect 120 132 123 135 
rect 120 135 123 138 
rect 120 138 123 141 
rect 120 141 123 144 
rect 120 144 123 147 
rect 120 147 123 150 
rect 120 150 123 153 
rect 120 153 123 156 
rect 120 156 123 159 
rect 120 159 123 162 
rect 120 162 123 165 
rect 120 165 123 168 
rect 120 168 123 171 
rect 120 171 123 174 
rect 120 174 123 177 
rect 120 177 123 180 
rect 120 180 123 183 
rect 120 183 123 186 
rect 120 186 123 189 
rect 120 189 123 192 
rect 120 192 123 195 
rect 120 195 123 198 
rect 120 198 123 201 
rect 120 201 123 204 
rect 120 204 123 207 
rect 120 207 123 210 
rect 120 210 123 213 
rect 120 213 123 216 
rect 120 216 123 219 
rect 120 219 123 222 
rect 120 222 123 225 
rect 120 225 123 228 
rect 120 228 123 231 
rect 120 231 123 234 
rect 120 234 123 237 
rect 120 237 123 240 
rect 120 240 123 243 
rect 120 243 123 246 
rect 120 246 123 249 
rect 120 249 123 252 
rect 120 252 123 255 
rect 120 255 123 258 
rect 120 258 123 261 
rect 120 261 123 264 
rect 120 264 123 267 
rect 120 267 123 270 
rect 120 270 123 273 
rect 120 273 123 276 
rect 120 276 123 279 
rect 120 279 123 282 
rect 120 282 123 285 
rect 120 285 123 288 
rect 120 288 123 291 
rect 120 291 123 294 
rect 120 294 123 297 
rect 120 297 123 300 
rect 120 300 123 303 
rect 120 303 123 306 
rect 120 306 123 309 
rect 120 309 123 312 
rect 120 312 123 315 
rect 120 315 123 318 
rect 120 318 123 321 
rect 120 321 123 324 
rect 120 324 123 327 
rect 120 327 123 330 
rect 120 330 123 333 
rect 120 333 123 336 
rect 120 336 123 339 
rect 120 339 123 342 
rect 120 342 123 345 
rect 120 345 123 348 
rect 120 348 123 351 
rect 120 351 123 354 
rect 120 354 123 357 
rect 120 357 123 360 
rect 120 360 123 363 
rect 120 363 123 366 
rect 120 366 123 369 
rect 120 369 123 372 
rect 120 372 123 375 
rect 120 375 123 378 
rect 120 378 123 381 
rect 120 381 123 384 
rect 120 384 123 387 
rect 120 387 123 390 
rect 120 390 123 393 
rect 120 393 123 396 
rect 120 396 123 399 
rect 120 399 123 402 
rect 120 402 123 405 
rect 120 405 123 408 
rect 120 408 123 411 
rect 120 411 123 414 
rect 120 414 123 417 
rect 120 417 123 420 
rect 120 420 123 423 
rect 120 423 123 426 
rect 120 426 123 429 
rect 120 429 123 432 
rect 120 432 123 435 
rect 120 435 123 438 
rect 120 438 123 441 
rect 120 441 123 444 
rect 120 444 123 447 
rect 120 447 123 450 
rect 120 450 123 453 
rect 120 453 123 456 
rect 120 456 123 459 
rect 120 459 123 462 
rect 120 462 123 465 
rect 120 465 123 468 
rect 120 468 123 471 
rect 120 471 123 474 
rect 120 474 123 477 
rect 120 477 123 480 
rect 120 480 123 483 
rect 120 483 123 486 
rect 120 486 123 489 
rect 120 489 123 492 
rect 120 492 123 495 
rect 120 495 123 498 
rect 120 498 123 501 
rect 120 501 123 504 
rect 120 504 123 507 
rect 120 507 123 510 
rect 123 0 126 3 
rect 123 3 126 6 
rect 123 6 126 9 
rect 123 9 126 12 
rect 123 12 126 15 
rect 123 15 126 18 
rect 123 18 126 21 
rect 123 21 126 24 
rect 123 24 126 27 
rect 123 27 126 30 
rect 123 30 126 33 
rect 123 33 126 36 
rect 123 36 126 39 
rect 123 39 126 42 
rect 123 42 126 45 
rect 123 45 126 48 
rect 123 48 126 51 
rect 123 51 126 54 
rect 123 54 126 57 
rect 123 57 126 60 
rect 123 60 126 63 
rect 123 63 126 66 
rect 123 66 126 69 
rect 123 69 126 72 
rect 123 72 126 75 
rect 123 75 126 78 
rect 123 78 126 81 
rect 123 81 126 84 
rect 123 84 126 87 
rect 123 87 126 90 
rect 123 90 126 93 
rect 123 93 126 96 
rect 123 96 126 99 
rect 123 99 126 102 
rect 123 102 126 105 
rect 123 105 126 108 
rect 123 108 126 111 
rect 123 111 126 114 
rect 123 114 126 117 
rect 123 117 126 120 
rect 123 120 126 123 
rect 123 123 126 126 
rect 123 126 126 129 
rect 123 129 126 132 
rect 123 132 126 135 
rect 123 135 126 138 
rect 123 138 126 141 
rect 123 141 126 144 
rect 123 144 126 147 
rect 123 147 126 150 
rect 123 150 126 153 
rect 123 153 126 156 
rect 123 156 126 159 
rect 123 159 126 162 
rect 123 162 126 165 
rect 123 165 126 168 
rect 123 168 126 171 
rect 123 171 126 174 
rect 123 174 126 177 
rect 123 177 126 180 
rect 123 180 126 183 
rect 123 183 126 186 
rect 123 186 126 189 
rect 123 189 126 192 
rect 123 192 126 195 
rect 123 195 126 198 
rect 123 198 126 201 
rect 123 201 126 204 
rect 123 204 126 207 
rect 123 207 126 210 
rect 123 210 126 213 
rect 123 213 126 216 
rect 123 216 126 219 
rect 123 219 126 222 
rect 123 222 126 225 
rect 123 225 126 228 
rect 123 228 126 231 
rect 123 231 126 234 
rect 123 234 126 237 
rect 123 237 126 240 
rect 123 240 126 243 
rect 123 243 126 246 
rect 123 246 126 249 
rect 123 249 126 252 
rect 123 252 126 255 
rect 123 255 126 258 
rect 123 258 126 261 
rect 123 261 126 264 
rect 123 264 126 267 
rect 123 267 126 270 
rect 123 270 126 273 
rect 123 273 126 276 
rect 123 276 126 279 
rect 123 279 126 282 
rect 123 282 126 285 
rect 123 285 126 288 
rect 123 288 126 291 
rect 123 291 126 294 
rect 123 294 126 297 
rect 123 297 126 300 
rect 123 300 126 303 
rect 123 303 126 306 
rect 123 306 126 309 
rect 123 309 126 312 
rect 123 312 126 315 
rect 123 315 126 318 
rect 123 318 126 321 
rect 123 321 126 324 
rect 123 324 126 327 
rect 123 327 126 330 
rect 123 330 126 333 
rect 123 333 126 336 
rect 123 336 126 339 
rect 123 339 126 342 
rect 123 342 126 345 
rect 123 345 126 348 
rect 123 348 126 351 
rect 123 351 126 354 
rect 123 354 126 357 
rect 123 357 126 360 
rect 123 360 126 363 
rect 123 363 126 366 
rect 123 366 126 369 
rect 123 369 126 372 
rect 123 372 126 375 
rect 123 375 126 378 
rect 123 378 126 381 
rect 123 381 126 384 
rect 123 384 126 387 
rect 123 387 126 390 
rect 123 390 126 393 
rect 123 393 126 396 
rect 123 396 126 399 
rect 123 399 126 402 
rect 123 402 126 405 
rect 123 405 126 408 
rect 123 408 126 411 
rect 123 411 126 414 
rect 123 414 126 417 
rect 123 417 126 420 
rect 123 420 126 423 
rect 123 423 126 426 
rect 123 426 126 429 
rect 123 429 126 432 
rect 123 432 126 435 
rect 123 435 126 438 
rect 123 438 126 441 
rect 123 441 126 444 
rect 123 444 126 447 
rect 123 447 126 450 
rect 123 450 126 453 
rect 123 453 126 456 
rect 123 456 126 459 
rect 123 459 126 462 
rect 123 462 126 465 
rect 123 465 126 468 
rect 123 468 126 471 
rect 123 471 126 474 
rect 123 474 126 477 
rect 123 477 126 480 
rect 123 480 126 483 
rect 123 483 126 486 
rect 123 486 126 489 
rect 123 489 126 492 
rect 123 492 126 495 
rect 123 495 126 498 
rect 123 498 126 501 
rect 123 501 126 504 
rect 123 504 126 507 
rect 123 507 126 510 
rect 126 0 129 3 
rect 126 3 129 6 
rect 126 6 129 9 
rect 126 9 129 12 
rect 126 12 129 15 
rect 126 15 129 18 
rect 126 18 129 21 
rect 126 21 129 24 
rect 126 24 129 27 
rect 126 27 129 30 
rect 126 30 129 33 
rect 126 33 129 36 
rect 126 36 129 39 
rect 126 39 129 42 
rect 126 42 129 45 
rect 126 45 129 48 
rect 126 48 129 51 
rect 126 51 129 54 
rect 126 54 129 57 
rect 126 57 129 60 
rect 126 60 129 63 
rect 126 63 129 66 
rect 126 66 129 69 
rect 126 69 129 72 
rect 126 72 129 75 
rect 126 75 129 78 
rect 126 78 129 81 
rect 126 81 129 84 
rect 126 84 129 87 
rect 126 87 129 90 
rect 126 90 129 93 
rect 126 93 129 96 
rect 126 96 129 99 
rect 126 99 129 102 
rect 126 102 129 105 
rect 126 105 129 108 
rect 126 108 129 111 
rect 126 111 129 114 
rect 126 114 129 117 
rect 126 117 129 120 
rect 126 120 129 123 
rect 126 123 129 126 
rect 126 126 129 129 
rect 126 129 129 132 
rect 126 132 129 135 
rect 126 135 129 138 
rect 126 138 129 141 
rect 126 141 129 144 
rect 126 144 129 147 
rect 126 147 129 150 
rect 126 150 129 153 
rect 126 153 129 156 
rect 126 156 129 159 
rect 126 159 129 162 
rect 126 162 129 165 
rect 126 165 129 168 
rect 126 168 129 171 
rect 126 171 129 174 
rect 126 174 129 177 
rect 126 177 129 180 
rect 126 180 129 183 
rect 126 183 129 186 
rect 126 186 129 189 
rect 126 189 129 192 
rect 126 192 129 195 
rect 126 195 129 198 
rect 126 198 129 201 
rect 126 201 129 204 
rect 126 204 129 207 
rect 126 207 129 210 
rect 126 210 129 213 
rect 126 213 129 216 
rect 126 216 129 219 
rect 126 219 129 222 
rect 126 222 129 225 
rect 126 225 129 228 
rect 126 228 129 231 
rect 126 231 129 234 
rect 126 234 129 237 
rect 126 237 129 240 
rect 126 240 129 243 
rect 126 243 129 246 
rect 126 246 129 249 
rect 126 249 129 252 
rect 126 252 129 255 
rect 126 255 129 258 
rect 126 258 129 261 
rect 126 261 129 264 
rect 126 264 129 267 
rect 126 267 129 270 
rect 126 270 129 273 
rect 126 273 129 276 
rect 126 276 129 279 
rect 126 279 129 282 
rect 126 282 129 285 
rect 126 285 129 288 
rect 126 288 129 291 
rect 126 291 129 294 
rect 126 294 129 297 
rect 126 297 129 300 
rect 126 300 129 303 
rect 126 303 129 306 
rect 126 306 129 309 
rect 126 309 129 312 
rect 126 312 129 315 
rect 126 315 129 318 
rect 126 318 129 321 
rect 126 321 129 324 
rect 126 324 129 327 
rect 126 327 129 330 
rect 126 330 129 333 
rect 126 333 129 336 
rect 126 336 129 339 
rect 126 339 129 342 
rect 126 342 129 345 
rect 126 345 129 348 
rect 126 348 129 351 
rect 126 351 129 354 
rect 126 354 129 357 
rect 126 357 129 360 
rect 126 360 129 363 
rect 126 363 129 366 
rect 126 366 129 369 
rect 126 369 129 372 
rect 126 372 129 375 
rect 126 375 129 378 
rect 126 378 129 381 
rect 126 381 129 384 
rect 126 384 129 387 
rect 126 387 129 390 
rect 126 390 129 393 
rect 126 393 129 396 
rect 126 396 129 399 
rect 126 399 129 402 
rect 126 402 129 405 
rect 126 405 129 408 
rect 126 408 129 411 
rect 126 411 129 414 
rect 126 414 129 417 
rect 126 417 129 420 
rect 126 420 129 423 
rect 126 423 129 426 
rect 126 426 129 429 
rect 126 429 129 432 
rect 126 432 129 435 
rect 126 435 129 438 
rect 126 438 129 441 
rect 126 441 129 444 
rect 126 444 129 447 
rect 126 447 129 450 
rect 126 450 129 453 
rect 126 453 129 456 
rect 126 456 129 459 
rect 126 459 129 462 
rect 126 462 129 465 
rect 126 465 129 468 
rect 126 468 129 471 
rect 126 471 129 474 
rect 126 474 129 477 
rect 126 477 129 480 
rect 126 480 129 483 
rect 126 483 129 486 
rect 126 486 129 489 
rect 126 489 129 492 
rect 126 492 129 495 
rect 126 495 129 498 
rect 126 498 129 501 
rect 126 501 129 504 
rect 126 504 129 507 
rect 126 507 129 510 
rect 129 0 132 3 
rect 129 3 132 6 
rect 129 6 132 9 
rect 129 9 132 12 
rect 129 12 132 15 
rect 129 15 132 18 
rect 129 18 132 21 
rect 129 21 132 24 
rect 129 24 132 27 
rect 129 27 132 30 
rect 129 30 132 33 
rect 129 33 132 36 
rect 129 36 132 39 
rect 129 39 132 42 
rect 129 42 132 45 
rect 129 45 132 48 
rect 129 48 132 51 
rect 129 51 132 54 
rect 129 54 132 57 
rect 129 57 132 60 
rect 129 60 132 63 
rect 129 63 132 66 
rect 129 66 132 69 
rect 129 69 132 72 
rect 129 72 132 75 
rect 129 75 132 78 
rect 129 78 132 81 
rect 129 81 132 84 
rect 129 84 132 87 
rect 129 87 132 90 
rect 129 90 132 93 
rect 129 93 132 96 
rect 129 96 132 99 
rect 129 99 132 102 
rect 129 102 132 105 
rect 129 105 132 108 
rect 129 108 132 111 
rect 129 111 132 114 
rect 129 114 132 117 
rect 129 117 132 120 
rect 129 120 132 123 
rect 129 123 132 126 
rect 129 126 132 129 
rect 129 129 132 132 
rect 129 132 132 135 
rect 129 135 132 138 
rect 129 138 132 141 
rect 129 141 132 144 
rect 129 144 132 147 
rect 129 147 132 150 
rect 129 150 132 153 
rect 129 153 132 156 
rect 129 156 132 159 
rect 129 159 132 162 
rect 129 162 132 165 
rect 129 165 132 168 
rect 129 168 132 171 
rect 129 171 132 174 
rect 129 174 132 177 
rect 129 177 132 180 
rect 129 180 132 183 
rect 129 183 132 186 
rect 129 186 132 189 
rect 129 189 132 192 
rect 129 192 132 195 
rect 129 195 132 198 
rect 129 198 132 201 
rect 129 201 132 204 
rect 129 204 132 207 
rect 129 207 132 210 
rect 129 210 132 213 
rect 129 213 132 216 
rect 129 216 132 219 
rect 129 219 132 222 
rect 129 222 132 225 
rect 129 225 132 228 
rect 129 228 132 231 
rect 129 231 132 234 
rect 129 234 132 237 
rect 129 237 132 240 
rect 129 240 132 243 
rect 129 243 132 246 
rect 129 246 132 249 
rect 129 249 132 252 
rect 129 252 132 255 
rect 129 255 132 258 
rect 129 258 132 261 
rect 129 261 132 264 
rect 129 264 132 267 
rect 129 267 132 270 
rect 129 270 132 273 
rect 129 273 132 276 
rect 129 276 132 279 
rect 129 279 132 282 
rect 129 282 132 285 
rect 129 285 132 288 
rect 129 288 132 291 
rect 129 291 132 294 
rect 129 294 132 297 
rect 129 297 132 300 
rect 129 300 132 303 
rect 129 303 132 306 
rect 129 306 132 309 
rect 129 309 132 312 
rect 129 312 132 315 
rect 129 315 132 318 
rect 129 318 132 321 
rect 129 321 132 324 
rect 129 324 132 327 
rect 129 327 132 330 
rect 129 330 132 333 
rect 129 333 132 336 
rect 129 336 132 339 
rect 129 339 132 342 
rect 129 342 132 345 
rect 129 345 132 348 
rect 129 348 132 351 
rect 129 351 132 354 
rect 129 354 132 357 
rect 129 357 132 360 
rect 129 360 132 363 
rect 129 363 132 366 
rect 129 366 132 369 
rect 129 369 132 372 
rect 129 372 132 375 
rect 129 375 132 378 
rect 129 378 132 381 
rect 129 381 132 384 
rect 129 384 132 387 
rect 129 387 132 390 
rect 129 390 132 393 
rect 129 393 132 396 
rect 129 396 132 399 
rect 129 399 132 402 
rect 129 402 132 405 
rect 129 405 132 408 
rect 129 408 132 411 
rect 129 411 132 414 
rect 129 414 132 417 
rect 129 417 132 420 
rect 129 420 132 423 
rect 129 423 132 426 
rect 129 426 132 429 
rect 129 429 132 432 
rect 129 432 132 435 
rect 129 435 132 438 
rect 129 438 132 441 
rect 129 441 132 444 
rect 129 444 132 447 
rect 129 447 132 450 
rect 129 450 132 453 
rect 129 453 132 456 
rect 129 456 132 459 
rect 129 459 132 462 
rect 129 462 132 465 
rect 129 465 132 468 
rect 129 468 132 471 
rect 129 471 132 474 
rect 129 474 132 477 
rect 129 477 132 480 
rect 129 480 132 483 
rect 129 483 132 486 
rect 129 486 132 489 
rect 129 489 132 492 
rect 129 492 132 495 
rect 129 495 132 498 
rect 129 498 132 501 
rect 129 501 132 504 
rect 129 504 132 507 
rect 129 507 132 510 
rect 132 0 135 3 
rect 132 3 135 6 
rect 132 6 135 9 
rect 132 9 135 12 
rect 132 12 135 15 
rect 132 15 135 18 
rect 132 18 135 21 
rect 132 21 135 24 
rect 132 24 135 27 
rect 132 27 135 30 
rect 132 30 135 33 
rect 132 33 135 36 
rect 132 36 135 39 
rect 132 39 135 42 
rect 132 42 135 45 
rect 132 45 135 48 
rect 132 48 135 51 
rect 132 51 135 54 
rect 132 54 135 57 
rect 132 57 135 60 
rect 132 60 135 63 
rect 132 63 135 66 
rect 132 66 135 69 
rect 132 69 135 72 
rect 132 72 135 75 
rect 132 75 135 78 
rect 132 78 135 81 
rect 132 81 135 84 
rect 132 84 135 87 
rect 132 87 135 90 
rect 132 90 135 93 
rect 132 93 135 96 
rect 132 96 135 99 
rect 132 99 135 102 
rect 132 102 135 105 
rect 132 105 135 108 
rect 132 108 135 111 
rect 132 111 135 114 
rect 132 114 135 117 
rect 132 117 135 120 
rect 132 120 135 123 
rect 132 123 135 126 
rect 132 126 135 129 
rect 132 129 135 132 
rect 132 132 135 135 
rect 132 135 135 138 
rect 132 138 135 141 
rect 132 141 135 144 
rect 132 144 135 147 
rect 132 147 135 150 
rect 132 150 135 153 
rect 132 153 135 156 
rect 132 156 135 159 
rect 132 159 135 162 
rect 132 162 135 165 
rect 132 165 135 168 
rect 132 168 135 171 
rect 132 171 135 174 
rect 132 174 135 177 
rect 132 177 135 180 
rect 132 180 135 183 
rect 132 183 135 186 
rect 132 186 135 189 
rect 132 189 135 192 
rect 132 192 135 195 
rect 132 195 135 198 
rect 132 198 135 201 
rect 132 201 135 204 
rect 132 204 135 207 
rect 132 207 135 210 
rect 132 210 135 213 
rect 132 213 135 216 
rect 132 216 135 219 
rect 132 219 135 222 
rect 132 222 135 225 
rect 132 225 135 228 
rect 132 228 135 231 
rect 132 231 135 234 
rect 132 234 135 237 
rect 132 237 135 240 
rect 132 240 135 243 
rect 132 243 135 246 
rect 132 246 135 249 
rect 132 249 135 252 
rect 132 252 135 255 
rect 132 255 135 258 
rect 132 258 135 261 
rect 132 261 135 264 
rect 132 264 135 267 
rect 132 267 135 270 
rect 132 270 135 273 
rect 132 273 135 276 
rect 132 276 135 279 
rect 132 279 135 282 
rect 132 282 135 285 
rect 132 285 135 288 
rect 132 288 135 291 
rect 132 291 135 294 
rect 132 294 135 297 
rect 132 297 135 300 
rect 132 300 135 303 
rect 132 303 135 306 
rect 132 306 135 309 
rect 132 309 135 312 
rect 132 312 135 315 
rect 132 315 135 318 
rect 132 318 135 321 
rect 132 321 135 324 
rect 132 324 135 327 
rect 132 327 135 330 
rect 132 330 135 333 
rect 132 333 135 336 
rect 132 336 135 339 
rect 132 339 135 342 
rect 132 342 135 345 
rect 132 345 135 348 
rect 132 348 135 351 
rect 132 351 135 354 
rect 132 354 135 357 
rect 132 357 135 360 
rect 132 360 135 363 
rect 132 363 135 366 
rect 132 366 135 369 
rect 132 369 135 372 
rect 132 372 135 375 
rect 132 375 135 378 
rect 132 378 135 381 
rect 132 381 135 384 
rect 132 384 135 387 
rect 132 387 135 390 
rect 132 390 135 393 
rect 132 393 135 396 
rect 132 396 135 399 
rect 132 399 135 402 
rect 132 402 135 405 
rect 132 405 135 408 
rect 132 408 135 411 
rect 132 411 135 414 
rect 132 414 135 417 
rect 132 417 135 420 
rect 132 420 135 423 
rect 132 423 135 426 
rect 132 426 135 429 
rect 132 429 135 432 
rect 132 432 135 435 
rect 132 435 135 438 
rect 132 438 135 441 
rect 132 441 135 444 
rect 132 444 135 447 
rect 132 447 135 450 
rect 132 450 135 453 
rect 132 453 135 456 
rect 132 456 135 459 
rect 132 459 135 462 
rect 132 462 135 465 
rect 132 465 135 468 
rect 132 468 135 471 
rect 132 471 135 474 
rect 132 474 135 477 
rect 132 477 135 480 
rect 132 480 135 483 
rect 132 483 135 486 
rect 132 486 135 489 
rect 132 489 135 492 
rect 132 492 135 495 
rect 132 495 135 498 
rect 132 498 135 501 
rect 132 501 135 504 
rect 132 504 135 507 
rect 132 507 135 510 
rect 135 0 138 3 
rect 135 3 138 6 
rect 135 6 138 9 
rect 135 9 138 12 
rect 135 12 138 15 
rect 135 15 138 18 
rect 135 18 138 21 
rect 135 21 138 24 
rect 135 24 138 27 
rect 135 27 138 30 
rect 135 30 138 33 
rect 135 33 138 36 
rect 135 36 138 39 
rect 135 39 138 42 
rect 135 42 138 45 
rect 135 45 138 48 
rect 135 48 138 51 
rect 135 51 138 54 
rect 135 54 138 57 
rect 135 57 138 60 
rect 135 60 138 63 
rect 135 63 138 66 
rect 135 66 138 69 
rect 135 69 138 72 
rect 135 72 138 75 
rect 135 75 138 78 
rect 135 78 138 81 
rect 135 81 138 84 
rect 135 84 138 87 
rect 135 87 138 90 
rect 135 90 138 93 
rect 135 93 138 96 
rect 135 96 138 99 
rect 135 99 138 102 
rect 135 102 138 105 
rect 135 105 138 108 
rect 135 108 138 111 
rect 135 111 138 114 
rect 135 114 138 117 
rect 135 117 138 120 
rect 135 120 138 123 
rect 135 123 138 126 
rect 135 126 138 129 
rect 135 129 138 132 
rect 135 132 138 135 
rect 135 135 138 138 
rect 135 138 138 141 
rect 135 141 138 144 
rect 135 144 138 147 
rect 135 147 138 150 
rect 135 150 138 153 
rect 135 153 138 156 
rect 135 156 138 159 
rect 135 159 138 162 
rect 135 162 138 165 
rect 135 165 138 168 
rect 135 168 138 171 
rect 135 171 138 174 
rect 135 174 138 177 
rect 135 177 138 180 
rect 135 180 138 183 
rect 135 183 138 186 
rect 135 186 138 189 
rect 135 189 138 192 
rect 135 192 138 195 
rect 135 195 138 198 
rect 135 198 138 201 
rect 135 201 138 204 
rect 135 204 138 207 
rect 135 207 138 210 
rect 135 210 138 213 
rect 135 213 138 216 
rect 135 216 138 219 
rect 135 219 138 222 
rect 135 222 138 225 
rect 135 225 138 228 
rect 135 228 138 231 
rect 135 231 138 234 
rect 135 234 138 237 
rect 135 237 138 240 
rect 135 240 138 243 
rect 135 243 138 246 
rect 135 246 138 249 
rect 135 249 138 252 
rect 135 252 138 255 
rect 135 255 138 258 
rect 135 258 138 261 
rect 135 261 138 264 
rect 135 264 138 267 
rect 135 267 138 270 
rect 135 270 138 273 
rect 135 273 138 276 
rect 135 276 138 279 
rect 135 279 138 282 
rect 135 282 138 285 
rect 135 285 138 288 
rect 135 288 138 291 
rect 135 291 138 294 
rect 135 294 138 297 
rect 135 297 138 300 
rect 135 300 138 303 
rect 135 303 138 306 
rect 135 306 138 309 
rect 135 309 138 312 
rect 135 312 138 315 
rect 135 315 138 318 
rect 135 318 138 321 
rect 135 321 138 324 
rect 135 324 138 327 
rect 135 327 138 330 
rect 135 330 138 333 
rect 135 333 138 336 
rect 135 336 138 339 
rect 135 339 138 342 
rect 135 342 138 345 
rect 135 345 138 348 
rect 135 348 138 351 
rect 135 351 138 354 
rect 135 354 138 357 
rect 135 357 138 360 
rect 135 360 138 363 
rect 135 363 138 366 
rect 135 366 138 369 
rect 135 369 138 372 
rect 135 372 138 375 
rect 135 375 138 378 
rect 135 378 138 381 
rect 135 381 138 384 
rect 135 384 138 387 
rect 135 387 138 390 
rect 135 390 138 393 
rect 135 393 138 396 
rect 135 396 138 399 
rect 135 399 138 402 
rect 135 402 138 405 
rect 135 405 138 408 
rect 135 408 138 411 
rect 135 411 138 414 
rect 135 414 138 417 
rect 135 417 138 420 
rect 135 420 138 423 
rect 135 423 138 426 
rect 135 426 138 429 
rect 135 429 138 432 
rect 135 432 138 435 
rect 135 435 138 438 
rect 135 438 138 441 
rect 135 441 138 444 
rect 135 444 138 447 
rect 135 447 138 450 
rect 135 450 138 453 
rect 135 453 138 456 
rect 135 456 138 459 
rect 135 459 138 462 
rect 135 462 138 465 
rect 135 465 138 468 
rect 135 468 138 471 
rect 135 471 138 474 
rect 135 474 138 477 
rect 135 477 138 480 
rect 135 480 138 483 
rect 135 483 138 486 
rect 135 486 138 489 
rect 135 489 138 492 
rect 135 492 138 495 
rect 135 495 138 498 
rect 135 498 138 501 
rect 135 501 138 504 
rect 135 504 138 507 
rect 135 507 138 510 
rect 138 0 141 3 
rect 138 3 141 6 
rect 138 6 141 9 
rect 138 9 141 12 
rect 138 12 141 15 
rect 138 15 141 18 
rect 138 18 141 21 
rect 138 21 141 24 
rect 138 24 141 27 
rect 138 27 141 30 
rect 138 30 141 33 
rect 138 33 141 36 
rect 138 36 141 39 
rect 138 39 141 42 
rect 138 42 141 45 
rect 138 45 141 48 
rect 138 48 141 51 
rect 138 51 141 54 
rect 138 54 141 57 
rect 138 57 141 60 
rect 138 60 141 63 
rect 138 63 141 66 
rect 138 66 141 69 
rect 138 69 141 72 
rect 138 72 141 75 
rect 138 75 141 78 
rect 138 78 141 81 
rect 138 81 141 84 
rect 138 84 141 87 
rect 138 87 141 90 
rect 138 90 141 93 
rect 138 93 141 96 
rect 138 96 141 99 
rect 138 99 141 102 
rect 138 102 141 105 
rect 138 105 141 108 
rect 138 108 141 111 
rect 138 111 141 114 
rect 138 114 141 117 
rect 138 117 141 120 
rect 138 120 141 123 
rect 138 123 141 126 
rect 138 126 141 129 
rect 138 129 141 132 
rect 138 132 141 135 
rect 138 135 141 138 
rect 138 138 141 141 
rect 138 141 141 144 
rect 138 144 141 147 
rect 138 147 141 150 
rect 138 150 141 153 
rect 138 153 141 156 
rect 138 156 141 159 
rect 138 159 141 162 
rect 138 162 141 165 
rect 138 165 141 168 
rect 138 168 141 171 
rect 138 171 141 174 
rect 138 174 141 177 
rect 138 177 141 180 
rect 138 180 141 183 
rect 138 183 141 186 
rect 138 186 141 189 
rect 138 189 141 192 
rect 138 192 141 195 
rect 138 195 141 198 
rect 138 198 141 201 
rect 138 201 141 204 
rect 138 204 141 207 
rect 138 207 141 210 
rect 138 210 141 213 
rect 138 213 141 216 
rect 138 216 141 219 
rect 138 219 141 222 
rect 138 222 141 225 
rect 138 225 141 228 
rect 138 228 141 231 
rect 138 231 141 234 
rect 138 234 141 237 
rect 138 237 141 240 
rect 138 240 141 243 
rect 138 243 141 246 
rect 138 246 141 249 
rect 138 249 141 252 
rect 138 252 141 255 
rect 138 255 141 258 
rect 138 258 141 261 
rect 138 261 141 264 
rect 138 264 141 267 
rect 138 267 141 270 
rect 138 270 141 273 
rect 138 273 141 276 
rect 138 276 141 279 
rect 138 279 141 282 
rect 138 282 141 285 
rect 138 285 141 288 
rect 138 288 141 291 
rect 138 291 141 294 
rect 138 294 141 297 
rect 138 297 141 300 
rect 138 300 141 303 
rect 138 303 141 306 
rect 138 306 141 309 
rect 138 309 141 312 
rect 138 312 141 315 
rect 138 315 141 318 
rect 138 318 141 321 
rect 138 321 141 324 
rect 138 324 141 327 
rect 138 327 141 330 
rect 138 330 141 333 
rect 138 333 141 336 
rect 138 336 141 339 
rect 138 339 141 342 
rect 138 342 141 345 
rect 138 345 141 348 
rect 138 348 141 351 
rect 138 351 141 354 
rect 138 354 141 357 
rect 138 357 141 360 
rect 138 360 141 363 
rect 138 363 141 366 
rect 138 366 141 369 
rect 138 369 141 372 
rect 138 372 141 375 
rect 138 375 141 378 
rect 138 378 141 381 
rect 138 381 141 384 
rect 138 384 141 387 
rect 138 387 141 390 
rect 138 390 141 393 
rect 138 393 141 396 
rect 138 396 141 399 
rect 138 399 141 402 
rect 138 402 141 405 
rect 138 405 141 408 
rect 138 408 141 411 
rect 138 411 141 414 
rect 138 414 141 417 
rect 138 417 141 420 
rect 138 420 141 423 
rect 138 423 141 426 
rect 138 426 141 429 
rect 138 429 141 432 
rect 138 432 141 435 
rect 138 435 141 438 
rect 138 438 141 441 
rect 138 441 141 444 
rect 138 444 141 447 
rect 138 447 141 450 
rect 138 450 141 453 
rect 138 453 141 456 
rect 138 456 141 459 
rect 138 459 141 462 
rect 138 462 141 465 
rect 138 465 141 468 
rect 138 468 141 471 
rect 138 471 141 474 
rect 138 474 141 477 
rect 138 477 141 480 
rect 138 480 141 483 
rect 138 483 141 486 
rect 138 486 141 489 
rect 138 489 141 492 
rect 138 492 141 495 
rect 138 495 141 498 
rect 138 498 141 501 
rect 138 501 141 504 
rect 138 504 141 507 
rect 138 507 141 510 
rect 141 0 144 3 
rect 141 3 144 6 
rect 141 6 144 9 
rect 141 9 144 12 
rect 141 12 144 15 
rect 141 15 144 18 
rect 141 18 144 21 
rect 141 21 144 24 
rect 141 24 144 27 
rect 141 27 144 30 
rect 141 30 144 33 
rect 141 33 144 36 
rect 141 36 144 39 
rect 141 39 144 42 
rect 141 42 144 45 
rect 141 45 144 48 
rect 141 48 144 51 
rect 141 51 144 54 
rect 141 54 144 57 
rect 141 57 144 60 
rect 141 60 144 63 
rect 141 63 144 66 
rect 141 66 144 69 
rect 141 69 144 72 
rect 141 72 144 75 
rect 141 75 144 78 
rect 141 78 144 81 
rect 141 81 144 84 
rect 141 84 144 87 
rect 141 87 144 90 
rect 141 90 144 93 
rect 141 93 144 96 
rect 141 96 144 99 
rect 141 99 144 102 
rect 141 102 144 105 
rect 141 105 144 108 
rect 141 108 144 111 
rect 141 111 144 114 
rect 141 114 144 117 
rect 141 117 144 120 
rect 141 120 144 123 
rect 141 123 144 126 
rect 141 126 144 129 
rect 141 129 144 132 
rect 141 132 144 135 
rect 141 135 144 138 
rect 141 138 144 141 
rect 141 141 144 144 
rect 141 144 144 147 
rect 141 147 144 150 
rect 141 150 144 153 
rect 141 153 144 156 
rect 141 156 144 159 
rect 141 159 144 162 
rect 141 162 144 165 
rect 141 165 144 168 
rect 141 168 144 171 
rect 141 171 144 174 
rect 141 174 144 177 
rect 141 177 144 180 
rect 141 180 144 183 
rect 141 183 144 186 
rect 141 186 144 189 
rect 141 189 144 192 
rect 141 192 144 195 
rect 141 195 144 198 
rect 141 198 144 201 
rect 141 201 144 204 
rect 141 204 144 207 
rect 141 207 144 210 
rect 141 210 144 213 
rect 141 213 144 216 
rect 141 216 144 219 
rect 141 219 144 222 
rect 141 222 144 225 
rect 141 225 144 228 
rect 141 228 144 231 
rect 141 231 144 234 
rect 141 234 144 237 
rect 141 237 144 240 
rect 141 240 144 243 
rect 141 243 144 246 
rect 141 246 144 249 
rect 141 249 144 252 
rect 141 252 144 255 
rect 141 255 144 258 
rect 141 258 144 261 
rect 141 261 144 264 
rect 141 264 144 267 
rect 141 267 144 270 
rect 141 270 144 273 
rect 141 273 144 276 
rect 141 276 144 279 
rect 141 279 144 282 
rect 141 282 144 285 
rect 141 285 144 288 
rect 141 288 144 291 
rect 141 291 144 294 
rect 141 294 144 297 
rect 141 297 144 300 
rect 141 300 144 303 
rect 141 303 144 306 
rect 141 306 144 309 
rect 141 309 144 312 
rect 141 312 144 315 
rect 141 315 144 318 
rect 141 318 144 321 
rect 141 321 144 324 
rect 141 324 144 327 
rect 141 327 144 330 
rect 141 330 144 333 
rect 141 333 144 336 
rect 141 336 144 339 
rect 141 339 144 342 
rect 141 342 144 345 
rect 141 345 144 348 
rect 141 348 144 351 
rect 141 351 144 354 
rect 141 354 144 357 
rect 141 357 144 360 
rect 141 360 144 363 
rect 141 363 144 366 
rect 141 366 144 369 
rect 141 369 144 372 
rect 141 372 144 375 
rect 141 375 144 378 
rect 141 378 144 381 
rect 141 381 144 384 
rect 141 384 144 387 
rect 141 387 144 390 
rect 141 390 144 393 
rect 141 393 144 396 
rect 141 396 144 399 
rect 141 399 144 402 
rect 141 402 144 405 
rect 141 405 144 408 
rect 141 408 144 411 
rect 141 411 144 414 
rect 141 414 144 417 
rect 141 417 144 420 
rect 141 420 144 423 
rect 141 423 144 426 
rect 141 426 144 429 
rect 141 429 144 432 
rect 141 432 144 435 
rect 141 435 144 438 
rect 141 438 144 441 
rect 141 441 144 444 
rect 141 444 144 447 
rect 141 447 144 450 
rect 141 450 144 453 
rect 141 453 144 456 
rect 141 456 144 459 
rect 141 459 144 462 
rect 141 462 144 465 
rect 141 465 144 468 
rect 141 468 144 471 
rect 141 471 144 474 
rect 141 474 144 477 
rect 141 477 144 480 
rect 141 480 144 483 
rect 141 483 144 486 
rect 141 486 144 489 
rect 141 489 144 492 
rect 141 492 144 495 
rect 141 495 144 498 
rect 141 498 144 501 
rect 141 501 144 504 
rect 141 504 144 507 
rect 141 507 144 510 
rect 144 0 147 3 
rect 144 3 147 6 
rect 144 6 147 9 
rect 144 9 147 12 
rect 144 12 147 15 
rect 144 15 147 18 
rect 144 18 147 21 
rect 144 21 147 24 
rect 144 24 147 27 
rect 144 27 147 30 
rect 144 30 147 33 
rect 144 33 147 36 
rect 144 36 147 39 
rect 144 39 147 42 
rect 144 42 147 45 
rect 144 45 147 48 
rect 144 48 147 51 
rect 144 51 147 54 
rect 144 54 147 57 
rect 144 57 147 60 
rect 144 60 147 63 
rect 144 63 147 66 
rect 144 66 147 69 
rect 144 69 147 72 
rect 144 72 147 75 
rect 144 75 147 78 
rect 144 78 147 81 
rect 144 81 147 84 
rect 144 84 147 87 
rect 144 87 147 90 
rect 144 90 147 93 
rect 144 93 147 96 
rect 144 96 147 99 
rect 144 99 147 102 
rect 144 102 147 105 
rect 144 105 147 108 
rect 144 108 147 111 
rect 144 111 147 114 
rect 144 114 147 117 
rect 144 117 147 120 
rect 144 120 147 123 
rect 144 123 147 126 
rect 144 126 147 129 
rect 144 129 147 132 
rect 144 132 147 135 
rect 144 135 147 138 
rect 144 138 147 141 
rect 144 141 147 144 
rect 144 144 147 147 
rect 144 147 147 150 
rect 144 150 147 153 
rect 144 153 147 156 
rect 144 156 147 159 
rect 144 159 147 162 
rect 144 162 147 165 
rect 144 165 147 168 
rect 144 168 147 171 
rect 144 171 147 174 
rect 144 174 147 177 
rect 144 177 147 180 
rect 144 180 147 183 
rect 144 183 147 186 
rect 144 186 147 189 
rect 144 189 147 192 
rect 144 192 147 195 
rect 144 195 147 198 
rect 144 198 147 201 
rect 144 201 147 204 
rect 144 204 147 207 
rect 144 207 147 210 
rect 144 210 147 213 
rect 144 213 147 216 
rect 144 216 147 219 
rect 144 219 147 222 
rect 144 222 147 225 
rect 144 225 147 228 
rect 144 228 147 231 
rect 144 231 147 234 
rect 144 234 147 237 
rect 144 237 147 240 
rect 144 240 147 243 
rect 144 243 147 246 
rect 144 246 147 249 
rect 144 249 147 252 
rect 144 252 147 255 
rect 144 255 147 258 
rect 144 258 147 261 
rect 144 261 147 264 
rect 144 264 147 267 
rect 144 267 147 270 
rect 144 270 147 273 
rect 144 273 147 276 
rect 144 276 147 279 
rect 144 279 147 282 
rect 144 282 147 285 
rect 144 285 147 288 
rect 144 288 147 291 
rect 144 291 147 294 
rect 144 294 147 297 
rect 144 297 147 300 
rect 144 300 147 303 
rect 144 303 147 306 
rect 144 306 147 309 
rect 144 309 147 312 
rect 144 312 147 315 
rect 144 315 147 318 
rect 144 318 147 321 
rect 144 321 147 324 
rect 144 324 147 327 
rect 144 327 147 330 
rect 144 330 147 333 
rect 144 333 147 336 
rect 144 336 147 339 
rect 144 339 147 342 
rect 144 342 147 345 
rect 144 345 147 348 
rect 144 348 147 351 
rect 144 351 147 354 
rect 144 354 147 357 
rect 144 357 147 360 
rect 144 360 147 363 
rect 144 363 147 366 
rect 144 366 147 369 
rect 144 369 147 372 
rect 144 372 147 375 
rect 144 375 147 378 
rect 144 378 147 381 
rect 144 381 147 384 
rect 144 384 147 387 
rect 144 387 147 390 
rect 144 390 147 393 
rect 144 393 147 396 
rect 144 396 147 399 
rect 144 399 147 402 
rect 144 402 147 405 
rect 144 405 147 408 
rect 144 408 147 411 
rect 144 411 147 414 
rect 144 414 147 417 
rect 144 417 147 420 
rect 144 420 147 423 
rect 144 423 147 426 
rect 144 426 147 429 
rect 144 429 147 432 
rect 144 432 147 435 
rect 144 435 147 438 
rect 144 438 147 441 
rect 144 441 147 444 
rect 144 444 147 447 
rect 144 447 147 450 
rect 144 450 147 453 
rect 144 453 147 456 
rect 144 456 147 459 
rect 144 459 147 462 
rect 144 462 147 465 
rect 144 465 147 468 
rect 144 468 147 471 
rect 144 471 147 474 
rect 144 474 147 477 
rect 144 477 147 480 
rect 144 480 147 483 
rect 144 483 147 486 
rect 144 486 147 489 
rect 144 489 147 492 
rect 144 492 147 495 
rect 144 495 147 498 
rect 144 498 147 501 
rect 144 501 147 504 
rect 144 504 147 507 
rect 144 507 147 510 
rect 147 0 150 3 
rect 147 3 150 6 
rect 147 6 150 9 
rect 147 9 150 12 
rect 147 12 150 15 
rect 147 15 150 18 
rect 147 18 150 21 
rect 147 21 150 24 
rect 147 24 150 27 
rect 147 27 150 30 
rect 147 30 150 33 
rect 147 33 150 36 
rect 147 36 150 39 
rect 147 39 150 42 
rect 147 42 150 45 
rect 147 45 150 48 
rect 147 48 150 51 
rect 147 51 150 54 
rect 147 54 150 57 
rect 147 57 150 60 
rect 147 60 150 63 
rect 147 63 150 66 
rect 147 66 150 69 
rect 147 69 150 72 
rect 147 72 150 75 
rect 147 75 150 78 
rect 147 78 150 81 
rect 147 81 150 84 
rect 147 84 150 87 
rect 147 87 150 90 
rect 147 90 150 93 
rect 147 93 150 96 
rect 147 96 150 99 
rect 147 99 150 102 
rect 147 102 150 105 
rect 147 105 150 108 
rect 147 108 150 111 
rect 147 111 150 114 
rect 147 114 150 117 
rect 147 117 150 120 
rect 147 120 150 123 
rect 147 123 150 126 
rect 147 126 150 129 
rect 147 129 150 132 
rect 147 132 150 135 
rect 147 135 150 138 
rect 147 138 150 141 
rect 147 141 150 144 
rect 147 144 150 147 
rect 147 147 150 150 
rect 147 150 150 153 
rect 147 153 150 156 
rect 147 156 150 159 
rect 147 159 150 162 
rect 147 162 150 165 
rect 147 165 150 168 
rect 147 168 150 171 
rect 147 171 150 174 
rect 147 174 150 177 
rect 147 177 150 180 
rect 147 180 150 183 
rect 147 183 150 186 
rect 147 186 150 189 
rect 147 189 150 192 
rect 147 192 150 195 
rect 147 195 150 198 
rect 147 198 150 201 
rect 147 201 150 204 
rect 147 204 150 207 
rect 147 207 150 210 
rect 147 210 150 213 
rect 147 213 150 216 
rect 147 216 150 219 
rect 147 219 150 222 
rect 147 222 150 225 
rect 147 225 150 228 
rect 147 228 150 231 
rect 147 231 150 234 
rect 147 234 150 237 
rect 147 237 150 240 
rect 147 240 150 243 
rect 147 243 150 246 
rect 147 246 150 249 
rect 147 249 150 252 
rect 147 252 150 255 
rect 147 255 150 258 
rect 147 258 150 261 
rect 147 261 150 264 
rect 147 264 150 267 
rect 147 267 150 270 
rect 147 270 150 273 
rect 147 273 150 276 
rect 147 276 150 279 
rect 147 279 150 282 
rect 147 282 150 285 
rect 147 285 150 288 
rect 147 288 150 291 
rect 147 291 150 294 
rect 147 294 150 297 
rect 147 297 150 300 
rect 147 300 150 303 
rect 147 303 150 306 
rect 147 306 150 309 
rect 147 309 150 312 
rect 147 312 150 315 
rect 147 315 150 318 
rect 147 318 150 321 
rect 147 321 150 324 
rect 147 324 150 327 
rect 147 327 150 330 
rect 147 330 150 333 
rect 147 333 150 336 
rect 147 336 150 339 
rect 147 339 150 342 
rect 147 342 150 345 
rect 147 345 150 348 
rect 147 348 150 351 
rect 147 351 150 354 
rect 147 354 150 357 
rect 147 357 150 360 
rect 147 360 150 363 
rect 147 363 150 366 
rect 147 366 150 369 
rect 147 369 150 372 
rect 147 372 150 375 
rect 147 375 150 378 
rect 147 378 150 381 
rect 147 381 150 384 
rect 147 384 150 387 
rect 147 387 150 390 
rect 147 390 150 393 
rect 147 393 150 396 
rect 147 396 150 399 
rect 147 399 150 402 
rect 147 402 150 405 
rect 147 405 150 408 
rect 147 408 150 411 
rect 147 411 150 414 
rect 147 414 150 417 
rect 147 417 150 420 
rect 147 420 150 423 
rect 147 423 150 426 
rect 147 426 150 429 
rect 147 429 150 432 
rect 147 432 150 435 
rect 147 435 150 438 
rect 147 438 150 441 
rect 147 441 150 444 
rect 147 444 150 447 
rect 147 447 150 450 
rect 147 450 150 453 
rect 147 453 150 456 
rect 147 456 150 459 
rect 147 459 150 462 
rect 147 462 150 465 
rect 147 465 150 468 
rect 147 468 150 471 
rect 147 471 150 474 
rect 147 474 150 477 
rect 147 477 150 480 
rect 147 480 150 483 
rect 147 483 150 486 
rect 147 486 150 489 
rect 147 489 150 492 
rect 147 492 150 495 
rect 147 495 150 498 
rect 147 498 150 501 
rect 147 501 150 504 
rect 147 504 150 507 
rect 147 507 150 510 
rect 150 0 153 3 
rect 150 3 153 6 
rect 150 6 153 9 
rect 150 9 153 12 
rect 150 12 153 15 
rect 150 15 153 18 
rect 150 18 153 21 
rect 150 21 153 24 
rect 150 24 153 27 
rect 150 27 153 30 
rect 150 30 153 33 
rect 150 33 153 36 
rect 150 36 153 39 
rect 150 39 153 42 
rect 150 42 153 45 
rect 150 45 153 48 
rect 150 48 153 51 
rect 150 51 153 54 
rect 150 54 153 57 
rect 150 57 153 60 
rect 150 60 153 63 
rect 150 63 153 66 
rect 150 66 153 69 
rect 150 69 153 72 
rect 150 72 153 75 
rect 150 75 153 78 
rect 150 78 153 81 
rect 150 81 153 84 
rect 150 84 153 87 
rect 150 87 153 90 
rect 150 90 153 93 
rect 150 93 153 96 
rect 150 96 153 99 
rect 150 99 153 102 
rect 150 102 153 105 
rect 150 105 153 108 
rect 150 108 153 111 
rect 150 111 153 114 
rect 150 114 153 117 
rect 150 117 153 120 
rect 150 120 153 123 
rect 150 123 153 126 
rect 150 126 153 129 
rect 150 129 153 132 
rect 150 132 153 135 
rect 150 135 153 138 
rect 150 138 153 141 
rect 150 141 153 144 
rect 150 144 153 147 
rect 150 147 153 150 
rect 150 150 153 153 
rect 150 153 153 156 
rect 150 156 153 159 
rect 150 159 153 162 
rect 150 162 153 165 
rect 150 165 153 168 
rect 150 168 153 171 
rect 150 171 153 174 
rect 150 174 153 177 
rect 150 177 153 180 
rect 150 180 153 183 
rect 150 183 153 186 
rect 150 186 153 189 
rect 150 189 153 192 
rect 150 192 153 195 
rect 150 195 153 198 
rect 150 198 153 201 
rect 150 201 153 204 
rect 150 204 153 207 
rect 150 207 153 210 
rect 150 210 153 213 
rect 150 213 153 216 
rect 150 216 153 219 
rect 150 219 153 222 
rect 150 222 153 225 
rect 150 225 153 228 
rect 150 228 153 231 
rect 150 231 153 234 
rect 150 234 153 237 
rect 150 237 153 240 
rect 150 240 153 243 
rect 150 243 153 246 
rect 150 246 153 249 
rect 150 249 153 252 
rect 150 252 153 255 
rect 150 255 153 258 
rect 150 258 153 261 
rect 150 261 153 264 
rect 150 264 153 267 
rect 150 267 153 270 
rect 150 270 153 273 
rect 150 273 153 276 
rect 150 276 153 279 
rect 150 279 153 282 
rect 150 282 153 285 
rect 150 285 153 288 
rect 150 288 153 291 
rect 150 291 153 294 
rect 150 294 153 297 
rect 150 297 153 300 
rect 150 300 153 303 
rect 150 303 153 306 
rect 150 306 153 309 
rect 150 309 153 312 
rect 150 312 153 315 
rect 150 315 153 318 
rect 150 318 153 321 
rect 150 321 153 324 
rect 150 324 153 327 
rect 150 327 153 330 
rect 150 330 153 333 
rect 150 333 153 336 
rect 150 336 153 339 
rect 150 339 153 342 
rect 150 342 153 345 
rect 150 345 153 348 
rect 150 348 153 351 
rect 150 351 153 354 
rect 150 354 153 357 
rect 150 357 153 360 
rect 150 360 153 363 
rect 150 363 153 366 
rect 150 366 153 369 
rect 150 369 153 372 
rect 150 372 153 375 
rect 150 375 153 378 
rect 150 378 153 381 
rect 150 381 153 384 
rect 150 384 153 387 
rect 150 387 153 390 
rect 150 390 153 393 
rect 150 393 153 396 
rect 150 396 153 399 
rect 150 399 153 402 
rect 150 402 153 405 
rect 150 405 153 408 
rect 150 408 153 411 
rect 150 411 153 414 
rect 150 414 153 417 
rect 150 417 153 420 
rect 150 420 153 423 
rect 150 423 153 426 
rect 150 426 153 429 
rect 150 429 153 432 
rect 150 432 153 435 
rect 150 435 153 438 
rect 150 438 153 441 
rect 150 441 153 444 
rect 150 444 153 447 
rect 150 447 153 450 
rect 150 450 153 453 
rect 150 453 153 456 
rect 150 456 153 459 
rect 150 459 153 462 
rect 150 462 153 465 
rect 150 465 153 468 
rect 150 468 153 471 
rect 150 471 153 474 
rect 150 474 153 477 
rect 150 477 153 480 
rect 150 480 153 483 
rect 150 483 153 486 
rect 150 486 153 489 
rect 150 489 153 492 
rect 150 492 153 495 
rect 150 495 153 498 
rect 150 498 153 501 
rect 150 501 153 504 
rect 150 504 153 507 
rect 150 507 153 510 
rect 153 0 156 3 
rect 153 3 156 6 
rect 153 6 156 9 
rect 153 9 156 12 
rect 153 12 156 15 
rect 153 15 156 18 
rect 153 18 156 21 
rect 153 21 156 24 
rect 153 24 156 27 
rect 153 27 156 30 
rect 153 30 156 33 
rect 153 33 156 36 
rect 153 36 156 39 
rect 153 39 156 42 
rect 153 42 156 45 
rect 153 45 156 48 
rect 153 48 156 51 
rect 153 51 156 54 
rect 153 54 156 57 
rect 153 57 156 60 
rect 153 60 156 63 
rect 153 63 156 66 
rect 153 66 156 69 
rect 153 69 156 72 
rect 153 72 156 75 
rect 153 75 156 78 
rect 153 78 156 81 
rect 153 81 156 84 
rect 153 84 156 87 
rect 153 87 156 90 
rect 153 90 156 93 
rect 153 93 156 96 
rect 153 96 156 99 
rect 153 99 156 102 
rect 153 102 156 105 
rect 153 105 156 108 
rect 153 108 156 111 
rect 153 111 156 114 
rect 153 114 156 117 
rect 153 117 156 120 
rect 153 120 156 123 
rect 153 123 156 126 
rect 153 126 156 129 
rect 153 129 156 132 
rect 153 132 156 135 
rect 153 135 156 138 
rect 153 138 156 141 
rect 153 141 156 144 
rect 153 144 156 147 
rect 153 147 156 150 
rect 153 150 156 153 
rect 153 153 156 156 
rect 153 156 156 159 
rect 153 159 156 162 
rect 153 162 156 165 
rect 153 165 156 168 
rect 153 168 156 171 
rect 153 171 156 174 
rect 153 174 156 177 
rect 153 177 156 180 
rect 153 180 156 183 
rect 153 183 156 186 
rect 153 186 156 189 
rect 153 189 156 192 
rect 153 192 156 195 
rect 153 195 156 198 
rect 153 198 156 201 
rect 153 201 156 204 
rect 153 204 156 207 
rect 153 207 156 210 
rect 153 210 156 213 
rect 153 213 156 216 
rect 153 216 156 219 
rect 153 219 156 222 
rect 153 222 156 225 
rect 153 225 156 228 
rect 153 228 156 231 
rect 153 231 156 234 
rect 153 234 156 237 
rect 153 237 156 240 
rect 153 240 156 243 
rect 153 243 156 246 
rect 153 246 156 249 
rect 153 249 156 252 
rect 153 252 156 255 
rect 153 255 156 258 
rect 153 258 156 261 
rect 153 261 156 264 
rect 153 264 156 267 
rect 153 267 156 270 
rect 153 270 156 273 
rect 153 273 156 276 
rect 153 276 156 279 
rect 153 279 156 282 
rect 153 282 156 285 
rect 153 285 156 288 
rect 153 288 156 291 
rect 153 291 156 294 
rect 153 294 156 297 
rect 153 297 156 300 
rect 153 300 156 303 
rect 153 303 156 306 
rect 153 306 156 309 
rect 153 309 156 312 
rect 153 312 156 315 
rect 153 315 156 318 
rect 153 318 156 321 
rect 153 321 156 324 
rect 153 324 156 327 
rect 153 327 156 330 
rect 153 330 156 333 
rect 153 333 156 336 
rect 153 336 156 339 
rect 153 339 156 342 
rect 153 342 156 345 
rect 153 345 156 348 
rect 153 348 156 351 
rect 153 351 156 354 
rect 153 354 156 357 
rect 153 357 156 360 
rect 153 360 156 363 
rect 153 363 156 366 
rect 153 366 156 369 
rect 153 369 156 372 
rect 153 372 156 375 
rect 153 375 156 378 
rect 153 378 156 381 
rect 153 381 156 384 
rect 153 384 156 387 
rect 153 387 156 390 
rect 153 390 156 393 
rect 153 393 156 396 
rect 153 396 156 399 
rect 153 399 156 402 
rect 153 402 156 405 
rect 153 405 156 408 
rect 153 408 156 411 
rect 153 411 156 414 
rect 153 414 156 417 
rect 153 417 156 420 
rect 153 420 156 423 
rect 153 423 156 426 
rect 153 426 156 429 
rect 153 429 156 432 
rect 153 432 156 435 
rect 153 435 156 438 
rect 153 438 156 441 
rect 153 441 156 444 
rect 153 444 156 447 
rect 153 447 156 450 
rect 153 450 156 453 
rect 153 453 156 456 
rect 153 456 156 459 
rect 153 459 156 462 
rect 153 462 156 465 
rect 153 465 156 468 
rect 153 468 156 471 
rect 153 471 156 474 
rect 153 474 156 477 
rect 153 477 156 480 
rect 153 480 156 483 
rect 153 483 156 486 
rect 153 486 156 489 
rect 153 489 156 492 
rect 153 492 156 495 
rect 153 495 156 498 
rect 153 498 156 501 
rect 153 501 156 504 
rect 153 504 156 507 
rect 153 507 156 510 
rect 156 0 159 3 
rect 156 3 159 6 
rect 156 6 159 9 
rect 156 9 159 12 
rect 156 12 159 15 
rect 156 15 159 18 
rect 156 18 159 21 
rect 156 21 159 24 
rect 156 24 159 27 
rect 156 27 159 30 
rect 156 30 159 33 
rect 156 33 159 36 
rect 156 36 159 39 
rect 156 39 159 42 
rect 156 42 159 45 
rect 156 45 159 48 
rect 156 48 159 51 
rect 156 51 159 54 
rect 156 54 159 57 
rect 156 57 159 60 
rect 156 60 159 63 
rect 156 63 159 66 
rect 156 66 159 69 
rect 156 69 159 72 
rect 156 72 159 75 
rect 156 75 159 78 
rect 156 78 159 81 
rect 156 81 159 84 
rect 156 84 159 87 
rect 156 87 159 90 
rect 156 90 159 93 
rect 156 93 159 96 
rect 156 96 159 99 
rect 156 99 159 102 
rect 156 102 159 105 
rect 156 105 159 108 
rect 156 108 159 111 
rect 156 111 159 114 
rect 156 114 159 117 
rect 156 117 159 120 
rect 156 120 159 123 
rect 156 123 159 126 
rect 156 126 159 129 
rect 156 129 159 132 
rect 156 132 159 135 
rect 156 135 159 138 
rect 156 138 159 141 
rect 156 141 159 144 
rect 156 144 159 147 
rect 156 147 159 150 
rect 156 150 159 153 
rect 156 153 159 156 
rect 156 156 159 159 
rect 156 159 159 162 
rect 156 162 159 165 
rect 156 165 159 168 
rect 156 168 159 171 
rect 156 171 159 174 
rect 156 174 159 177 
rect 156 177 159 180 
rect 156 180 159 183 
rect 156 183 159 186 
rect 156 186 159 189 
rect 156 189 159 192 
rect 156 192 159 195 
rect 156 195 159 198 
rect 156 198 159 201 
rect 156 201 159 204 
rect 156 204 159 207 
rect 156 207 159 210 
rect 156 210 159 213 
rect 156 213 159 216 
rect 156 216 159 219 
rect 156 219 159 222 
rect 156 222 159 225 
rect 156 225 159 228 
rect 156 228 159 231 
rect 156 231 159 234 
rect 156 234 159 237 
rect 156 237 159 240 
rect 156 240 159 243 
rect 156 243 159 246 
rect 156 246 159 249 
rect 156 249 159 252 
rect 156 252 159 255 
rect 156 255 159 258 
rect 156 258 159 261 
rect 156 261 159 264 
rect 156 264 159 267 
rect 156 267 159 270 
rect 156 270 159 273 
rect 156 273 159 276 
rect 156 276 159 279 
rect 156 279 159 282 
rect 156 282 159 285 
rect 156 285 159 288 
rect 156 288 159 291 
rect 156 291 159 294 
rect 156 294 159 297 
rect 156 297 159 300 
rect 156 300 159 303 
rect 156 303 159 306 
rect 156 306 159 309 
rect 156 309 159 312 
rect 156 312 159 315 
rect 156 315 159 318 
rect 156 318 159 321 
rect 156 321 159 324 
rect 156 324 159 327 
rect 156 327 159 330 
rect 156 330 159 333 
rect 156 333 159 336 
rect 156 336 159 339 
rect 156 339 159 342 
rect 156 342 159 345 
rect 156 345 159 348 
rect 156 348 159 351 
rect 156 351 159 354 
rect 156 354 159 357 
rect 156 357 159 360 
rect 156 360 159 363 
rect 156 363 159 366 
rect 156 366 159 369 
rect 156 369 159 372 
rect 156 372 159 375 
rect 156 375 159 378 
rect 156 378 159 381 
rect 156 381 159 384 
rect 156 384 159 387 
rect 156 387 159 390 
rect 156 390 159 393 
rect 156 393 159 396 
rect 156 396 159 399 
rect 156 399 159 402 
rect 156 402 159 405 
rect 156 405 159 408 
rect 156 408 159 411 
rect 156 411 159 414 
rect 156 414 159 417 
rect 156 417 159 420 
rect 156 420 159 423 
rect 156 423 159 426 
rect 156 426 159 429 
rect 156 429 159 432 
rect 156 432 159 435 
rect 156 435 159 438 
rect 156 438 159 441 
rect 156 441 159 444 
rect 156 444 159 447 
rect 156 447 159 450 
rect 156 450 159 453 
rect 156 453 159 456 
rect 156 456 159 459 
rect 156 459 159 462 
rect 156 462 159 465 
rect 156 465 159 468 
rect 156 468 159 471 
rect 156 471 159 474 
rect 156 474 159 477 
rect 156 477 159 480 
rect 156 480 159 483 
rect 156 483 159 486 
rect 156 486 159 489 
rect 156 489 159 492 
rect 156 492 159 495 
rect 156 495 159 498 
rect 156 498 159 501 
rect 156 501 159 504 
rect 156 504 159 507 
rect 156 507 159 510 
rect 159 0 162 3 
rect 159 3 162 6 
rect 159 6 162 9 
rect 159 9 162 12 
rect 159 12 162 15 
rect 159 15 162 18 
rect 159 18 162 21 
rect 159 21 162 24 
rect 159 24 162 27 
rect 159 27 162 30 
rect 159 30 162 33 
rect 159 33 162 36 
rect 159 36 162 39 
rect 159 39 162 42 
rect 159 42 162 45 
rect 159 45 162 48 
rect 159 48 162 51 
rect 159 51 162 54 
rect 159 54 162 57 
rect 159 57 162 60 
rect 159 60 162 63 
rect 159 63 162 66 
rect 159 66 162 69 
rect 159 69 162 72 
rect 159 72 162 75 
rect 159 75 162 78 
rect 159 78 162 81 
rect 159 81 162 84 
rect 159 84 162 87 
rect 159 87 162 90 
rect 159 90 162 93 
rect 159 93 162 96 
rect 159 96 162 99 
rect 159 99 162 102 
rect 159 102 162 105 
rect 159 105 162 108 
rect 159 108 162 111 
rect 159 111 162 114 
rect 159 114 162 117 
rect 159 117 162 120 
rect 159 120 162 123 
rect 159 123 162 126 
rect 159 126 162 129 
rect 159 129 162 132 
rect 159 132 162 135 
rect 159 135 162 138 
rect 159 138 162 141 
rect 159 141 162 144 
rect 159 144 162 147 
rect 159 147 162 150 
rect 159 150 162 153 
rect 159 153 162 156 
rect 159 156 162 159 
rect 159 159 162 162 
rect 159 162 162 165 
rect 159 165 162 168 
rect 159 168 162 171 
rect 159 171 162 174 
rect 159 174 162 177 
rect 159 177 162 180 
rect 159 180 162 183 
rect 159 183 162 186 
rect 159 186 162 189 
rect 159 189 162 192 
rect 159 192 162 195 
rect 159 195 162 198 
rect 159 198 162 201 
rect 159 201 162 204 
rect 159 204 162 207 
rect 159 207 162 210 
rect 159 210 162 213 
rect 159 213 162 216 
rect 159 216 162 219 
rect 159 219 162 222 
rect 159 222 162 225 
rect 159 225 162 228 
rect 159 228 162 231 
rect 159 231 162 234 
rect 159 234 162 237 
rect 159 237 162 240 
rect 159 240 162 243 
rect 159 243 162 246 
rect 159 246 162 249 
rect 159 249 162 252 
rect 159 252 162 255 
rect 159 255 162 258 
rect 159 258 162 261 
rect 159 261 162 264 
rect 159 264 162 267 
rect 159 267 162 270 
rect 159 270 162 273 
rect 159 273 162 276 
rect 159 276 162 279 
rect 159 279 162 282 
rect 159 282 162 285 
rect 159 285 162 288 
rect 159 288 162 291 
rect 159 291 162 294 
rect 159 294 162 297 
rect 159 297 162 300 
rect 159 300 162 303 
rect 159 303 162 306 
rect 159 306 162 309 
rect 159 309 162 312 
rect 159 312 162 315 
rect 159 315 162 318 
rect 159 318 162 321 
rect 159 321 162 324 
rect 159 324 162 327 
rect 159 327 162 330 
rect 159 330 162 333 
rect 159 333 162 336 
rect 159 336 162 339 
rect 159 339 162 342 
rect 159 342 162 345 
rect 159 345 162 348 
rect 159 348 162 351 
rect 159 351 162 354 
rect 159 354 162 357 
rect 159 357 162 360 
rect 159 360 162 363 
rect 159 363 162 366 
rect 159 366 162 369 
rect 159 369 162 372 
rect 159 372 162 375 
rect 159 375 162 378 
rect 159 378 162 381 
rect 159 381 162 384 
rect 159 384 162 387 
rect 159 387 162 390 
rect 159 390 162 393 
rect 159 393 162 396 
rect 159 396 162 399 
rect 159 399 162 402 
rect 159 402 162 405 
rect 159 405 162 408 
rect 159 408 162 411 
rect 159 411 162 414 
rect 159 414 162 417 
rect 159 417 162 420 
rect 159 420 162 423 
rect 159 423 162 426 
rect 159 426 162 429 
rect 159 429 162 432 
rect 159 432 162 435 
rect 159 435 162 438 
rect 159 438 162 441 
rect 159 441 162 444 
rect 159 444 162 447 
rect 159 447 162 450 
rect 159 450 162 453 
rect 159 453 162 456 
rect 159 456 162 459 
rect 159 459 162 462 
rect 159 462 162 465 
rect 159 465 162 468 
rect 159 468 162 471 
rect 159 471 162 474 
rect 159 474 162 477 
rect 159 477 162 480 
rect 159 480 162 483 
rect 159 483 162 486 
rect 159 486 162 489 
rect 159 489 162 492 
rect 159 492 162 495 
rect 159 495 162 498 
rect 159 498 162 501 
rect 159 501 162 504 
rect 159 504 162 507 
rect 159 507 162 510 
rect 162 0 165 3 
rect 162 3 165 6 
rect 162 6 165 9 
rect 162 9 165 12 
rect 162 12 165 15 
rect 162 15 165 18 
rect 162 18 165 21 
rect 162 21 165 24 
rect 162 24 165 27 
rect 162 27 165 30 
rect 162 30 165 33 
rect 162 33 165 36 
rect 162 36 165 39 
rect 162 39 165 42 
rect 162 42 165 45 
rect 162 45 165 48 
rect 162 48 165 51 
rect 162 51 165 54 
rect 162 54 165 57 
rect 162 57 165 60 
rect 162 60 165 63 
rect 162 63 165 66 
rect 162 66 165 69 
rect 162 69 165 72 
rect 162 72 165 75 
rect 162 75 165 78 
rect 162 78 165 81 
rect 162 81 165 84 
rect 162 84 165 87 
rect 162 87 165 90 
rect 162 90 165 93 
rect 162 93 165 96 
rect 162 96 165 99 
rect 162 99 165 102 
rect 162 102 165 105 
rect 162 105 165 108 
rect 162 108 165 111 
rect 162 111 165 114 
rect 162 114 165 117 
rect 162 117 165 120 
rect 162 120 165 123 
rect 162 123 165 126 
rect 162 126 165 129 
rect 162 129 165 132 
rect 162 132 165 135 
rect 162 135 165 138 
rect 162 138 165 141 
rect 162 141 165 144 
rect 162 144 165 147 
rect 162 147 165 150 
rect 162 150 165 153 
rect 162 153 165 156 
rect 162 156 165 159 
rect 162 159 165 162 
rect 162 162 165 165 
rect 162 165 165 168 
rect 162 168 165 171 
rect 162 171 165 174 
rect 162 174 165 177 
rect 162 177 165 180 
rect 162 180 165 183 
rect 162 183 165 186 
rect 162 186 165 189 
rect 162 189 165 192 
rect 162 192 165 195 
rect 162 195 165 198 
rect 162 198 165 201 
rect 162 201 165 204 
rect 162 204 165 207 
rect 162 207 165 210 
rect 162 210 165 213 
rect 162 213 165 216 
rect 162 216 165 219 
rect 162 219 165 222 
rect 162 222 165 225 
rect 162 225 165 228 
rect 162 228 165 231 
rect 162 231 165 234 
rect 162 234 165 237 
rect 162 237 165 240 
rect 162 240 165 243 
rect 162 243 165 246 
rect 162 246 165 249 
rect 162 249 165 252 
rect 162 252 165 255 
rect 162 255 165 258 
rect 162 258 165 261 
rect 162 261 165 264 
rect 162 264 165 267 
rect 162 267 165 270 
rect 162 270 165 273 
rect 162 273 165 276 
rect 162 276 165 279 
rect 162 279 165 282 
rect 162 282 165 285 
rect 162 285 165 288 
rect 162 288 165 291 
rect 162 291 165 294 
rect 162 294 165 297 
rect 162 297 165 300 
rect 162 300 165 303 
rect 162 303 165 306 
rect 162 306 165 309 
rect 162 309 165 312 
rect 162 312 165 315 
rect 162 315 165 318 
rect 162 318 165 321 
rect 162 321 165 324 
rect 162 324 165 327 
rect 162 327 165 330 
rect 162 330 165 333 
rect 162 333 165 336 
rect 162 336 165 339 
rect 162 339 165 342 
rect 162 342 165 345 
rect 162 345 165 348 
rect 162 348 165 351 
rect 162 351 165 354 
rect 162 354 165 357 
rect 162 357 165 360 
rect 162 360 165 363 
rect 162 363 165 366 
rect 162 366 165 369 
rect 162 369 165 372 
rect 162 372 165 375 
rect 162 375 165 378 
rect 162 378 165 381 
rect 162 381 165 384 
rect 162 384 165 387 
rect 162 387 165 390 
rect 162 390 165 393 
rect 162 393 165 396 
rect 162 396 165 399 
rect 162 399 165 402 
rect 162 402 165 405 
rect 162 405 165 408 
rect 162 408 165 411 
rect 162 411 165 414 
rect 162 414 165 417 
rect 162 417 165 420 
rect 162 420 165 423 
rect 162 423 165 426 
rect 162 426 165 429 
rect 162 429 165 432 
rect 162 432 165 435 
rect 162 435 165 438 
rect 162 438 165 441 
rect 162 441 165 444 
rect 162 444 165 447 
rect 162 447 165 450 
rect 162 450 165 453 
rect 162 453 165 456 
rect 162 456 165 459 
rect 162 459 165 462 
rect 162 462 165 465 
rect 162 465 165 468 
rect 162 468 165 471 
rect 162 471 165 474 
rect 162 474 165 477 
rect 162 477 165 480 
rect 162 480 165 483 
rect 162 483 165 486 
rect 162 486 165 489 
rect 162 489 165 492 
rect 162 492 165 495 
rect 162 495 165 498 
rect 162 498 165 501 
rect 162 501 165 504 
rect 162 504 165 507 
rect 162 507 165 510 
rect 165 0 168 3 
rect 165 3 168 6 
rect 165 6 168 9 
rect 165 9 168 12 
rect 165 12 168 15 
rect 165 15 168 18 
rect 165 18 168 21 
rect 165 21 168 24 
rect 165 24 168 27 
rect 165 27 168 30 
rect 165 30 168 33 
rect 165 33 168 36 
rect 165 36 168 39 
rect 165 39 168 42 
rect 165 42 168 45 
rect 165 45 168 48 
rect 165 48 168 51 
rect 165 51 168 54 
rect 165 54 168 57 
rect 165 57 168 60 
rect 165 60 168 63 
rect 165 63 168 66 
rect 165 66 168 69 
rect 165 69 168 72 
rect 165 72 168 75 
rect 165 75 168 78 
rect 165 78 168 81 
rect 165 81 168 84 
rect 165 84 168 87 
rect 165 87 168 90 
rect 165 90 168 93 
rect 165 93 168 96 
rect 165 96 168 99 
rect 165 99 168 102 
rect 165 102 168 105 
rect 165 105 168 108 
rect 165 108 168 111 
rect 165 111 168 114 
rect 165 114 168 117 
rect 165 117 168 120 
rect 165 120 168 123 
rect 165 123 168 126 
rect 165 126 168 129 
rect 165 129 168 132 
rect 165 132 168 135 
rect 165 135 168 138 
rect 165 138 168 141 
rect 165 141 168 144 
rect 165 144 168 147 
rect 165 147 168 150 
rect 165 150 168 153 
rect 165 153 168 156 
rect 165 156 168 159 
rect 165 159 168 162 
rect 165 162 168 165 
rect 165 165 168 168 
rect 165 168 168 171 
rect 165 171 168 174 
rect 165 174 168 177 
rect 165 177 168 180 
rect 165 180 168 183 
rect 165 183 168 186 
rect 165 186 168 189 
rect 165 189 168 192 
rect 165 192 168 195 
rect 165 195 168 198 
rect 165 198 168 201 
rect 165 201 168 204 
rect 165 204 168 207 
rect 165 207 168 210 
rect 165 210 168 213 
rect 165 213 168 216 
rect 165 216 168 219 
rect 165 219 168 222 
rect 165 222 168 225 
rect 165 225 168 228 
rect 165 228 168 231 
rect 165 231 168 234 
rect 165 234 168 237 
rect 165 237 168 240 
rect 165 240 168 243 
rect 165 243 168 246 
rect 165 246 168 249 
rect 165 249 168 252 
rect 165 252 168 255 
rect 165 255 168 258 
rect 165 258 168 261 
rect 165 261 168 264 
rect 165 264 168 267 
rect 165 267 168 270 
rect 165 270 168 273 
rect 165 273 168 276 
rect 165 276 168 279 
rect 165 279 168 282 
rect 165 282 168 285 
rect 165 285 168 288 
rect 165 288 168 291 
rect 165 291 168 294 
rect 165 294 168 297 
rect 165 297 168 300 
rect 165 300 168 303 
rect 165 303 168 306 
rect 165 306 168 309 
rect 165 309 168 312 
rect 165 312 168 315 
rect 165 315 168 318 
rect 165 318 168 321 
rect 165 321 168 324 
rect 165 324 168 327 
rect 165 327 168 330 
rect 165 330 168 333 
rect 165 333 168 336 
rect 165 336 168 339 
rect 165 339 168 342 
rect 165 342 168 345 
rect 165 345 168 348 
rect 165 348 168 351 
rect 165 351 168 354 
rect 165 354 168 357 
rect 165 357 168 360 
rect 165 360 168 363 
rect 165 363 168 366 
rect 165 366 168 369 
rect 165 369 168 372 
rect 165 372 168 375 
rect 165 375 168 378 
rect 165 378 168 381 
rect 165 381 168 384 
rect 165 384 168 387 
rect 165 387 168 390 
rect 165 390 168 393 
rect 165 393 168 396 
rect 165 396 168 399 
rect 165 399 168 402 
rect 165 402 168 405 
rect 165 405 168 408 
rect 165 408 168 411 
rect 165 411 168 414 
rect 165 414 168 417 
rect 165 417 168 420 
rect 165 420 168 423 
rect 165 423 168 426 
rect 165 426 168 429 
rect 165 429 168 432 
rect 165 432 168 435 
rect 165 435 168 438 
rect 165 438 168 441 
rect 165 441 168 444 
rect 165 444 168 447 
rect 165 447 168 450 
rect 165 450 168 453 
rect 165 453 168 456 
rect 165 456 168 459 
rect 165 459 168 462 
rect 165 462 168 465 
rect 165 465 168 468 
rect 165 468 168 471 
rect 165 471 168 474 
rect 165 474 168 477 
rect 165 477 168 480 
rect 165 480 168 483 
rect 165 483 168 486 
rect 165 486 168 489 
rect 165 489 168 492 
rect 165 492 168 495 
rect 165 495 168 498 
rect 165 498 168 501 
rect 165 501 168 504 
rect 165 504 168 507 
rect 165 507 168 510 
rect 168 0 171 3 
rect 168 3 171 6 
rect 168 6 171 9 
rect 168 9 171 12 
rect 168 12 171 15 
rect 168 15 171 18 
rect 168 18 171 21 
rect 168 21 171 24 
rect 168 24 171 27 
rect 168 27 171 30 
rect 168 30 171 33 
rect 168 33 171 36 
rect 168 36 171 39 
rect 168 39 171 42 
rect 168 42 171 45 
rect 168 45 171 48 
rect 168 48 171 51 
rect 168 51 171 54 
rect 168 54 171 57 
rect 168 57 171 60 
rect 168 60 171 63 
rect 168 63 171 66 
rect 168 66 171 69 
rect 168 69 171 72 
rect 168 72 171 75 
rect 168 75 171 78 
rect 168 78 171 81 
rect 168 81 171 84 
rect 168 84 171 87 
rect 168 87 171 90 
rect 168 90 171 93 
rect 168 93 171 96 
rect 168 96 171 99 
rect 168 99 171 102 
rect 168 102 171 105 
rect 168 105 171 108 
rect 168 108 171 111 
rect 168 111 171 114 
rect 168 114 171 117 
rect 168 117 171 120 
rect 168 120 171 123 
rect 168 123 171 126 
rect 168 126 171 129 
rect 168 129 171 132 
rect 168 132 171 135 
rect 168 135 171 138 
rect 168 138 171 141 
rect 168 141 171 144 
rect 168 144 171 147 
rect 168 147 171 150 
rect 168 150 171 153 
rect 168 153 171 156 
rect 168 156 171 159 
rect 168 159 171 162 
rect 168 162 171 165 
rect 168 165 171 168 
rect 168 168 171 171 
rect 168 171 171 174 
rect 168 174 171 177 
rect 168 177 171 180 
rect 168 180 171 183 
rect 168 183 171 186 
rect 168 186 171 189 
rect 168 189 171 192 
rect 168 192 171 195 
rect 168 195 171 198 
rect 168 198 171 201 
rect 168 201 171 204 
rect 168 204 171 207 
rect 168 207 171 210 
rect 168 210 171 213 
rect 168 213 171 216 
rect 168 216 171 219 
rect 168 219 171 222 
rect 168 222 171 225 
rect 168 225 171 228 
rect 168 228 171 231 
rect 168 231 171 234 
rect 168 234 171 237 
rect 168 237 171 240 
rect 168 240 171 243 
rect 168 243 171 246 
rect 168 246 171 249 
rect 168 249 171 252 
rect 168 252 171 255 
rect 168 255 171 258 
rect 168 258 171 261 
rect 168 261 171 264 
rect 168 264 171 267 
rect 168 267 171 270 
rect 168 270 171 273 
rect 168 273 171 276 
rect 168 276 171 279 
rect 168 279 171 282 
rect 168 282 171 285 
rect 168 285 171 288 
rect 168 288 171 291 
rect 168 291 171 294 
rect 168 294 171 297 
rect 168 297 171 300 
rect 168 300 171 303 
rect 168 303 171 306 
rect 168 306 171 309 
rect 168 309 171 312 
rect 168 312 171 315 
rect 168 315 171 318 
rect 168 318 171 321 
rect 168 321 171 324 
rect 168 324 171 327 
rect 168 327 171 330 
rect 168 330 171 333 
rect 168 333 171 336 
rect 168 336 171 339 
rect 168 339 171 342 
rect 168 342 171 345 
rect 168 345 171 348 
rect 168 348 171 351 
rect 168 351 171 354 
rect 168 354 171 357 
rect 168 357 171 360 
rect 168 360 171 363 
rect 168 363 171 366 
rect 168 366 171 369 
rect 168 369 171 372 
rect 168 372 171 375 
rect 168 375 171 378 
rect 168 378 171 381 
rect 168 381 171 384 
rect 168 384 171 387 
rect 168 387 171 390 
rect 168 390 171 393 
rect 168 393 171 396 
rect 168 396 171 399 
rect 168 399 171 402 
rect 168 402 171 405 
rect 168 405 171 408 
rect 168 408 171 411 
rect 168 411 171 414 
rect 168 414 171 417 
rect 168 417 171 420 
rect 168 420 171 423 
rect 168 423 171 426 
rect 168 426 171 429 
rect 168 429 171 432 
rect 168 432 171 435 
rect 168 435 171 438 
rect 168 438 171 441 
rect 168 441 171 444 
rect 168 444 171 447 
rect 168 447 171 450 
rect 168 450 171 453 
rect 168 453 171 456 
rect 168 456 171 459 
rect 168 459 171 462 
rect 168 462 171 465 
rect 168 465 171 468 
rect 168 468 171 471 
rect 168 471 171 474 
rect 168 474 171 477 
rect 168 477 171 480 
rect 168 480 171 483 
rect 168 483 171 486 
rect 168 486 171 489 
rect 168 489 171 492 
rect 168 492 171 495 
rect 168 495 171 498 
rect 168 498 171 501 
rect 168 501 171 504 
rect 168 504 171 507 
rect 168 507 171 510 
rect 171 0 174 3 
rect 171 3 174 6 
rect 171 6 174 9 
rect 171 9 174 12 
rect 171 12 174 15 
rect 171 15 174 18 
rect 171 18 174 21 
rect 171 21 174 24 
rect 171 24 174 27 
rect 171 27 174 30 
rect 171 30 174 33 
rect 171 33 174 36 
rect 171 36 174 39 
rect 171 39 174 42 
rect 171 42 174 45 
rect 171 45 174 48 
rect 171 48 174 51 
rect 171 51 174 54 
rect 171 54 174 57 
rect 171 57 174 60 
rect 171 60 174 63 
rect 171 63 174 66 
rect 171 66 174 69 
rect 171 69 174 72 
rect 171 72 174 75 
rect 171 75 174 78 
rect 171 78 174 81 
rect 171 81 174 84 
rect 171 84 174 87 
rect 171 87 174 90 
rect 171 90 174 93 
rect 171 93 174 96 
rect 171 96 174 99 
rect 171 99 174 102 
rect 171 102 174 105 
rect 171 105 174 108 
rect 171 108 174 111 
rect 171 111 174 114 
rect 171 114 174 117 
rect 171 117 174 120 
rect 171 120 174 123 
rect 171 123 174 126 
rect 171 126 174 129 
rect 171 129 174 132 
rect 171 132 174 135 
rect 171 135 174 138 
rect 171 138 174 141 
rect 171 141 174 144 
rect 171 144 174 147 
rect 171 147 174 150 
rect 171 150 174 153 
rect 171 153 174 156 
rect 171 156 174 159 
rect 171 159 174 162 
rect 171 162 174 165 
rect 171 165 174 168 
rect 171 168 174 171 
rect 171 171 174 174 
rect 171 174 174 177 
rect 171 177 174 180 
rect 171 180 174 183 
rect 171 183 174 186 
rect 171 186 174 189 
rect 171 189 174 192 
rect 171 192 174 195 
rect 171 195 174 198 
rect 171 198 174 201 
rect 171 201 174 204 
rect 171 204 174 207 
rect 171 207 174 210 
rect 171 210 174 213 
rect 171 213 174 216 
rect 171 216 174 219 
rect 171 219 174 222 
rect 171 222 174 225 
rect 171 225 174 228 
rect 171 228 174 231 
rect 171 231 174 234 
rect 171 234 174 237 
rect 171 237 174 240 
rect 171 240 174 243 
rect 171 243 174 246 
rect 171 246 174 249 
rect 171 249 174 252 
rect 171 252 174 255 
rect 171 255 174 258 
rect 171 258 174 261 
rect 171 261 174 264 
rect 171 264 174 267 
rect 171 267 174 270 
rect 171 270 174 273 
rect 171 273 174 276 
rect 171 276 174 279 
rect 171 279 174 282 
rect 171 282 174 285 
rect 171 285 174 288 
rect 171 288 174 291 
rect 171 291 174 294 
rect 171 294 174 297 
rect 171 297 174 300 
rect 171 300 174 303 
rect 171 303 174 306 
rect 171 306 174 309 
rect 171 309 174 312 
rect 171 312 174 315 
rect 171 315 174 318 
rect 171 318 174 321 
rect 171 321 174 324 
rect 171 324 174 327 
rect 171 327 174 330 
rect 171 330 174 333 
rect 171 333 174 336 
rect 171 336 174 339 
rect 171 339 174 342 
rect 171 342 174 345 
rect 171 345 174 348 
rect 171 348 174 351 
rect 171 351 174 354 
rect 171 354 174 357 
rect 171 357 174 360 
rect 171 360 174 363 
rect 171 363 174 366 
rect 171 366 174 369 
rect 171 369 174 372 
rect 171 372 174 375 
rect 171 375 174 378 
rect 171 378 174 381 
rect 171 381 174 384 
rect 171 384 174 387 
rect 171 387 174 390 
rect 171 390 174 393 
rect 171 393 174 396 
rect 171 396 174 399 
rect 171 399 174 402 
rect 171 402 174 405 
rect 171 405 174 408 
rect 171 408 174 411 
rect 171 411 174 414 
rect 171 414 174 417 
rect 171 417 174 420 
rect 171 420 174 423 
rect 171 423 174 426 
rect 171 426 174 429 
rect 171 429 174 432 
rect 171 432 174 435 
rect 171 435 174 438 
rect 171 438 174 441 
rect 171 441 174 444 
rect 171 444 174 447 
rect 171 447 174 450 
rect 171 450 174 453 
rect 171 453 174 456 
rect 171 456 174 459 
rect 171 459 174 462 
rect 171 462 174 465 
rect 171 465 174 468 
rect 171 468 174 471 
rect 171 471 174 474 
rect 171 474 174 477 
rect 171 477 174 480 
rect 171 480 174 483 
rect 171 483 174 486 
rect 171 486 174 489 
rect 171 489 174 492 
rect 171 492 174 495 
rect 171 495 174 498 
rect 171 498 174 501 
rect 171 501 174 504 
rect 171 504 174 507 
rect 171 507 174 510 
rect 174 0 177 3 
rect 174 3 177 6 
rect 174 6 177 9 
rect 174 9 177 12 
rect 174 12 177 15 
rect 174 15 177 18 
rect 174 18 177 21 
rect 174 21 177 24 
rect 174 24 177 27 
rect 174 27 177 30 
rect 174 30 177 33 
rect 174 33 177 36 
rect 174 36 177 39 
rect 174 39 177 42 
rect 174 42 177 45 
rect 174 45 177 48 
rect 174 48 177 51 
rect 174 51 177 54 
rect 174 54 177 57 
rect 174 57 177 60 
rect 174 60 177 63 
rect 174 63 177 66 
rect 174 66 177 69 
rect 174 69 177 72 
rect 174 72 177 75 
rect 174 75 177 78 
rect 174 78 177 81 
rect 174 81 177 84 
rect 174 84 177 87 
rect 174 87 177 90 
rect 174 90 177 93 
rect 174 93 177 96 
rect 174 96 177 99 
rect 174 99 177 102 
rect 174 102 177 105 
rect 174 105 177 108 
rect 174 108 177 111 
rect 174 111 177 114 
rect 174 114 177 117 
rect 174 117 177 120 
rect 174 120 177 123 
rect 174 123 177 126 
rect 174 126 177 129 
rect 174 129 177 132 
rect 174 132 177 135 
rect 174 135 177 138 
rect 174 138 177 141 
rect 174 141 177 144 
rect 174 144 177 147 
rect 174 147 177 150 
rect 174 150 177 153 
rect 174 153 177 156 
rect 174 156 177 159 
rect 174 159 177 162 
rect 174 162 177 165 
rect 174 165 177 168 
rect 174 168 177 171 
rect 174 171 177 174 
rect 174 174 177 177 
rect 174 177 177 180 
rect 174 180 177 183 
rect 174 183 177 186 
rect 174 186 177 189 
rect 174 189 177 192 
rect 174 192 177 195 
rect 174 195 177 198 
rect 174 198 177 201 
rect 174 201 177 204 
rect 174 204 177 207 
rect 174 207 177 210 
rect 174 210 177 213 
rect 174 213 177 216 
rect 174 216 177 219 
rect 174 219 177 222 
rect 174 222 177 225 
rect 174 225 177 228 
rect 174 228 177 231 
rect 174 231 177 234 
rect 174 234 177 237 
rect 174 237 177 240 
rect 174 240 177 243 
rect 174 243 177 246 
rect 174 246 177 249 
rect 174 249 177 252 
rect 174 252 177 255 
rect 174 255 177 258 
rect 174 258 177 261 
rect 174 261 177 264 
rect 174 264 177 267 
rect 174 267 177 270 
rect 174 270 177 273 
rect 174 273 177 276 
rect 174 276 177 279 
rect 174 279 177 282 
rect 174 282 177 285 
rect 174 285 177 288 
rect 174 288 177 291 
rect 174 291 177 294 
rect 174 294 177 297 
rect 174 297 177 300 
rect 174 300 177 303 
rect 174 303 177 306 
rect 174 306 177 309 
rect 174 309 177 312 
rect 174 312 177 315 
rect 174 315 177 318 
rect 174 318 177 321 
rect 174 321 177 324 
rect 174 324 177 327 
rect 174 327 177 330 
rect 174 330 177 333 
rect 174 333 177 336 
rect 174 336 177 339 
rect 174 339 177 342 
rect 174 342 177 345 
rect 174 345 177 348 
rect 174 348 177 351 
rect 174 351 177 354 
rect 174 354 177 357 
rect 174 357 177 360 
rect 174 360 177 363 
rect 174 363 177 366 
rect 174 366 177 369 
rect 174 369 177 372 
rect 174 372 177 375 
rect 174 375 177 378 
rect 174 378 177 381 
rect 174 381 177 384 
rect 174 384 177 387 
rect 174 387 177 390 
rect 174 390 177 393 
rect 174 393 177 396 
rect 174 396 177 399 
rect 174 399 177 402 
rect 174 402 177 405 
rect 174 405 177 408 
rect 174 408 177 411 
rect 174 411 177 414 
rect 174 414 177 417 
rect 174 417 177 420 
rect 174 420 177 423 
rect 174 423 177 426 
rect 174 426 177 429 
rect 174 429 177 432 
rect 174 432 177 435 
rect 174 435 177 438 
rect 174 438 177 441 
rect 174 441 177 444 
rect 174 444 177 447 
rect 174 447 177 450 
rect 174 450 177 453 
rect 174 453 177 456 
rect 174 456 177 459 
rect 174 459 177 462 
rect 174 462 177 465 
rect 174 465 177 468 
rect 174 468 177 471 
rect 174 471 177 474 
rect 174 474 177 477 
rect 174 477 177 480 
rect 174 480 177 483 
rect 174 483 177 486 
rect 174 486 177 489 
rect 174 489 177 492 
rect 174 492 177 495 
rect 174 495 177 498 
rect 174 498 177 501 
rect 174 501 177 504 
rect 174 504 177 507 
rect 174 507 177 510 
rect 177 0 180 3 
rect 177 3 180 6 
rect 177 6 180 9 
rect 177 9 180 12 
rect 177 12 180 15 
rect 177 15 180 18 
rect 177 18 180 21 
rect 177 21 180 24 
rect 177 24 180 27 
rect 177 27 180 30 
rect 177 30 180 33 
rect 177 33 180 36 
rect 177 36 180 39 
rect 177 39 180 42 
rect 177 42 180 45 
rect 177 45 180 48 
rect 177 48 180 51 
rect 177 51 180 54 
rect 177 54 180 57 
rect 177 57 180 60 
rect 177 60 180 63 
rect 177 63 180 66 
rect 177 66 180 69 
rect 177 69 180 72 
rect 177 72 180 75 
rect 177 75 180 78 
rect 177 78 180 81 
rect 177 81 180 84 
rect 177 84 180 87 
rect 177 87 180 90 
rect 177 90 180 93 
rect 177 93 180 96 
rect 177 96 180 99 
rect 177 99 180 102 
rect 177 102 180 105 
rect 177 105 180 108 
rect 177 108 180 111 
rect 177 111 180 114 
rect 177 114 180 117 
rect 177 117 180 120 
rect 177 120 180 123 
rect 177 123 180 126 
rect 177 126 180 129 
rect 177 129 180 132 
rect 177 132 180 135 
rect 177 135 180 138 
rect 177 138 180 141 
rect 177 141 180 144 
rect 177 144 180 147 
rect 177 147 180 150 
rect 177 150 180 153 
rect 177 153 180 156 
rect 177 156 180 159 
rect 177 159 180 162 
rect 177 162 180 165 
rect 177 165 180 168 
rect 177 168 180 171 
rect 177 171 180 174 
rect 177 174 180 177 
rect 177 177 180 180 
rect 177 180 180 183 
rect 177 183 180 186 
rect 177 186 180 189 
rect 177 189 180 192 
rect 177 192 180 195 
rect 177 195 180 198 
rect 177 198 180 201 
rect 177 201 180 204 
rect 177 204 180 207 
rect 177 207 180 210 
rect 177 210 180 213 
rect 177 213 180 216 
rect 177 216 180 219 
rect 177 219 180 222 
rect 177 222 180 225 
rect 177 225 180 228 
rect 177 228 180 231 
rect 177 231 180 234 
rect 177 234 180 237 
rect 177 237 180 240 
rect 177 240 180 243 
rect 177 243 180 246 
rect 177 246 180 249 
rect 177 249 180 252 
rect 177 252 180 255 
rect 177 255 180 258 
rect 177 258 180 261 
rect 177 261 180 264 
rect 177 264 180 267 
rect 177 267 180 270 
rect 177 270 180 273 
rect 177 273 180 276 
rect 177 276 180 279 
rect 177 279 180 282 
rect 177 282 180 285 
rect 177 285 180 288 
rect 177 288 180 291 
rect 177 291 180 294 
rect 177 294 180 297 
rect 177 297 180 300 
rect 177 300 180 303 
rect 177 303 180 306 
rect 177 306 180 309 
rect 177 309 180 312 
rect 177 312 180 315 
rect 177 315 180 318 
rect 177 318 180 321 
rect 177 321 180 324 
rect 177 324 180 327 
rect 177 327 180 330 
rect 177 330 180 333 
rect 177 333 180 336 
rect 177 336 180 339 
rect 177 339 180 342 
rect 177 342 180 345 
rect 177 345 180 348 
rect 177 348 180 351 
rect 177 351 180 354 
rect 177 354 180 357 
rect 177 357 180 360 
rect 177 360 180 363 
rect 177 363 180 366 
rect 177 366 180 369 
rect 177 369 180 372 
rect 177 372 180 375 
rect 177 375 180 378 
rect 177 378 180 381 
rect 177 381 180 384 
rect 177 384 180 387 
rect 177 387 180 390 
rect 177 390 180 393 
rect 177 393 180 396 
rect 177 396 180 399 
rect 177 399 180 402 
rect 177 402 180 405 
rect 177 405 180 408 
rect 177 408 180 411 
rect 177 411 180 414 
rect 177 414 180 417 
rect 177 417 180 420 
rect 177 420 180 423 
rect 177 423 180 426 
rect 177 426 180 429 
rect 177 429 180 432 
rect 177 432 180 435 
rect 177 435 180 438 
rect 177 438 180 441 
rect 177 441 180 444 
rect 177 444 180 447 
rect 177 447 180 450 
rect 177 450 180 453 
rect 177 453 180 456 
rect 177 456 180 459 
rect 177 459 180 462 
rect 177 462 180 465 
rect 177 465 180 468 
rect 177 468 180 471 
rect 177 471 180 474 
rect 177 474 180 477 
rect 177 477 180 480 
rect 177 480 180 483 
rect 177 483 180 486 
rect 177 486 180 489 
rect 177 489 180 492 
rect 177 492 180 495 
rect 177 495 180 498 
rect 177 498 180 501 
rect 177 501 180 504 
rect 177 504 180 507 
rect 177 507 180 510 
rect 180 0 183 3 
rect 180 3 183 6 
rect 180 6 183 9 
rect 180 9 183 12 
rect 180 12 183 15 
rect 180 15 183 18 
rect 180 18 183 21 
rect 180 21 183 24 
rect 180 24 183 27 
rect 180 27 183 30 
rect 180 30 183 33 
rect 180 33 183 36 
rect 180 36 183 39 
rect 180 39 183 42 
rect 180 42 183 45 
rect 180 45 183 48 
rect 180 48 183 51 
rect 180 51 183 54 
rect 180 54 183 57 
rect 180 57 183 60 
rect 180 60 183 63 
rect 180 63 183 66 
rect 180 66 183 69 
rect 180 69 183 72 
rect 180 72 183 75 
rect 180 75 183 78 
rect 180 78 183 81 
rect 180 81 183 84 
rect 180 84 183 87 
rect 180 87 183 90 
rect 180 90 183 93 
rect 180 93 183 96 
rect 180 96 183 99 
rect 180 99 183 102 
rect 180 102 183 105 
rect 180 105 183 108 
rect 180 108 183 111 
rect 180 111 183 114 
rect 180 114 183 117 
rect 180 117 183 120 
rect 180 120 183 123 
rect 180 123 183 126 
rect 180 126 183 129 
rect 180 129 183 132 
rect 180 132 183 135 
rect 180 135 183 138 
rect 180 138 183 141 
rect 180 141 183 144 
rect 180 144 183 147 
rect 180 147 183 150 
rect 180 150 183 153 
rect 180 153 183 156 
rect 180 156 183 159 
rect 180 159 183 162 
rect 180 162 183 165 
rect 180 165 183 168 
rect 180 168 183 171 
rect 180 171 183 174 
rect 180 174 183 177 
rect 180 177 183 180 
rect 180 180 183 183 
rect 180 183 183 186 
rect 180 186 183 189 
rect 180 189 183 192 
rect 180 192 183 195 
rect 180 195 183 198 
rect 180 198 183 201 
rect 180 201 183 204 
rect 180 204 183 207 
rect 180 207 183 210 
rect 180 210 183 213 
rect 180 213 183 216 
rect 180 216 183 219 
rect 180 219 183 222 
rect 180 222 183 225 
rect 180 225 183 228 
rect 180 228 183 231 
rect 180 231 183 234 
rect 180 234 183 237 
rect 180 237 183 240 
rect 180 240 183 243 
rect 180 243 183 246 
rect 180 246 183 249 
rect 180 249 183 252 
rect 180 252 183 255 
rect 180 255 183 258 
rect 180 258 183 261 
rect 180 261 183 264 
rect 180 264 183 267 
rect 180 267 183 270 
rect 180 270 183 273 
rect 180 273 183 276 
rect 180 276 183 279 
rect 180 279 183 282 
rect 180 282 183 285 
rect 180 285 183 288 
rect 180 288 183 291 
rect 180 291 183 294 
rect 180 294 183 297 
rect 180 297 183 300 
rect 180 300 183 303 
rect 180 303 183 306 
rect 180 306 183 309 
rect 180 309 183 312 
rect 180 312 183 315 
rect 180 315 183 318 
rect 180 318 183 321 
rect 180 321 183 324 
rect 180 324 183 327 
rect 180 327 183 330 
rect 180 330 183 333 
rect 180 333 183 336 
rect 180 336 183 339 
rect 180 339 183 342 
rect 180 342 183 345 
rect 180 345 183 348 
rect 180 348 183 351 
rect 180 351 183 354 
rect 180 354 183 357 
rect 180 357 183 360 
rect 180 360 183 363 
rect 180 363 183 366 
rect 180 366 183 369 
rect 180 369 183 372 
rect 180 372 183 375 
rect 180 375 183 378 
rect 180 378 183 381 
rect 180 381 183 384 
rect 180 384 183 387 
rect 180 387 183 390 
rect 180 390 183 393 
rect 180 393 183 396 
rect 180 396 183 399 
rect 180 399 183 402 
rect 180 402 183 405 
rect 180 405 183 408 
rect 180 408 183 411 
rect 180 411 183 414 
rect 180 414 183 417 
rect 180 417 183 420 
rect 180 420 183 423 
rect 180 423 183 426 
rect 180 426 183 429 
rect 180 429 183 432 
rect 180 432 183 435 
rect 180 435 183 438 
rect 180 438 183 441 
rect 180 441 183 444 
rect 180 444 183 447 
rect 180 447 183 450 
rect 180 450 183 453 
rect 180 453 183 456 
rect 180 456 183 459 
rect 180 459 183 462 
rect 180 462 183 465 
rect 180 465 183 468 
rect 180 468 183 471 
rect 180 471 183 474 
rect 180 474 183 477 
rect 180 477 183 480 
rect 180 480 183 483 
rect 180 483 183 486 
rect 180 486 183 489 
rect 180 489 183 492 
rect 180 492 183 495 
rect 180 495 183 498 
rect 180 498 183 501 
rect 180 501 183 504 
rect 180 504 183 507 
rect 180 507 183 510 
rect 183 0 186 3 
rect 183 3 186 6 
rect 183 6 186 9 
rect 183 9 186 12 
rect 183 12 186 15 
rect 183 15 186 18 
rect 183 18 186 21 
rect 183 21 186 24 
rect 183 24 186 27 
rect 183 27 186 30 
rect 183 30 186 33 
rect 183 33 186 36 
rect 183 36 186 39 
rect 183 39 186 42 
rect 183 42 186 45 
rect 183 45 186 48 
rect 183 48 186 51 
rect 183 51 186 54 
rect 183 54 186 57 
rect 183 57 186 60 
rect 183 60 186 63 
rect 183 63 186 66 
rect 183 66 186 69 
rect 183 69 186 72 
rect 183 72 186 75 
rect 183 75 186 78 
rect 183 78 186 81 
rect 183 81 186 84 
rect 183 84 186 87 
rect 183 87 186 90 
rect 183 90 186 93 
rect 183 93 186 96 
rect 183 96 186 99 
rect 183 99 186 102 
rect 183 102 186 105 
rect 183 105 186 108 
rect 183 108 186 111 
rect 183 111 186 114 
rect 183 114 186 117 
rect 183 117 186 120 
rect 183 120 186 123 
rect 183 123 186 126 
rect 183 126 186 129 
rect 183 129 186 132 
rect 183 132 186 135 
rect 183 135 186 138 
rect 183 138 186 141 
rect 183 141 186 144 
rect 183 144 186 147 
rect 183 147 186 150 
rect 183 150 186 153 
rect 183 153 186 156 
rect 183 156 186 159 
rect 183 159 186 162 
rect 183 162 186 165 
rect 183 165 186 168 
rect 183 168 186 171 
rect 183 171 186 174 
rect 183 174 186 177 
rect 183 177 186 180 
rect 183 180 186 183 
rect 183 183 186 186 
rect 183 186 186 189 
rect 183 189 186 192 
rect 183 192 186 195 
rect 183 195 186 198 
rect 183 198 186 201 
rect 183 201 186 204 
rect 183 204 186 207 
rect 183 207 186 210 
rect 183 210 186 213 
rect 183 213 186 216 
rect 183 216 186 219 
rect 183 219 186 222 
rect 183 222 186 225 
rect 183 225 186 228 
rect 183 228 186 231 
rect 183 231 186 234 
rect 183 234 186 237 
rect 183 237 186 240 
rect 183 240 186 243 
rect 183 243 186 246 
rect 183 246 186 249 
rect 183 249 186 252 
rect 183 252 186 255 
rect 183 255 186 258 
rect 183 258 186 261 
rect 183 261 186 264 
rect 183 264 186 267 
rect 183 267 186 270 
rect 183 270 186 273 
rect 183 273 186 276 
rect 183 276 186 279 
rect 183 279 186 282 
rect 183 282 186 285 
rect 183 285 186 288 
rect 183 288 186 291 
rect 183 291 186 294 
rect 183 294 186 297 
rect 183 297 186 300 
rect 183 300 186 303 
rect 183 303 186 306 
rect 183 306 186 309 
rect 183 309 186 312 
rect 183 312 186 315 
rect 183 315 186 318 
rect 183 318 186 321 
rect 183 321 186 324 
rect 183 324 186 327 
rect 183 327 186 330 
rect 183 330 186 333 
rect 183 333 186 336 
rect 183 336 186 339 
rect 183 339 186 342 
rect 183 342 186 345 
rect 183 345 186 348 
rect 183 348 186 351 
rect 183 351 186 354 
rect 183 354 186 357 
rect 183 357 186 360 
rect 183 360 186 363 
rect 183 363 186 366 
rect 183 366 186 369 
rect 183 369 186 372 
rect 183 372 186 375 
rect 183 375 186 378 
rect 183 378 186 381 
rect 183 381 186 384 
rect 183 384 186 387 
rect 183 387 186 390 
rect 183 390 186 393 
rect 183 393 186 396 
rect 183 396 186 399 
rect 183 399 186 402 
rect 183 402 186 405 
rect 183 405 186 408 
rect 183 408 186 411 
rect 183 411 186 414 
rect 183 414 186 417 
rect 183 417 186 420 
rect 183 420 186 423 
rect 183 423 186 426 
rect 183 426 186 429 
rect 183 429 186 432 
rect 183 432 186 435 
rect 183 435 186 438 
rect 183 438 186 441 
rect 183 441 186 444 
rect 183 444 186 447 
rect 183 447 186 450 
rect 183 450 186 453 
rect 183 453 186 456 
rect 183 456 186 459 
rect 183 459 186 462 
rect 183 462 186 465 
rect 183 465 186 468 
rect 183 468 186 471 
rect 183 471 186 474 
rect 183 474 186 477 
rect 183 477 186 480 
rect 183 480 186 483 
rect 183 483 186 486 
rect 183 486 186 489 
rect 183 489 186 492 
rect 183 492 186 495 
rect 183 495 186 498 
rect 183 498 186 501 
rect 183 501 186 504 
rect 183 504 186 507 
rect 183 507 186 510 
rect 186 0 189 3 
rect 186 3 189 6 
rect 186 6 189 9 
rect 186 9 189 12 
rect 186 12 189 15 
rect 186 15 189 18 
rect 186 18 189 21 
rect 186 21 189 24 
rect 186 24 189 27 
rect 186 27 189 30 
rect 186 30 189 33 
rect 186 33 189 36 
rect 186 36 189 39 
rect 186 39 189 42 
rect 186 42 189 45 
rect 186 45 189 48 
rect 186 48 189 51 
rect 186 51 189 54 
rect 186 54 189 57 
rect 186 57 189 60 
rect 186 60 189 63 
rect 186 63 189 66 
rect 186 66 189 69 
rect 186 69 189 72 
rect 186 72 189 75 
rect 186 75 189 78 
rect 186 78 189 81 
rect 186 81 189 84 
rect 186 84 189 87 
rect 186 87 189 90 
rect 186 90 189 93 
rect 186 93 189 96 
rect 186 96 189 99 
rect 186 99 189 102 
rect 186 102 189 105 
rect 186 105 189 108 
rect 186 108 189 111 
rect 186 111 189 114 
rect 186 114 189 117 
rect 186 117 189 120 
rect 186 120 189 123 
rect 186 123 189 126 
rect 186 126 189 129 
rect 186 129 189 132 
rect 186 132 189 135 
rect 186 135 189 138 
rect 186 138 189 141 
rect 186 141 189 144 
rect 186 144 189 147 
rect 186 147 189 150 
rect 186 150 189 153 
rect 186 153 189 156 
rect 186 156 189 159 
rect 186 159 189 162 
rect 186 162 189 165 
rect 186 165 189 168 
rect 186 168 189 171 
rect 186 171 189 174 
rect 186 174 189 177 
rect 186 177 189 180 
rect 186 180 189 183 
rect 186 183 189 186 
rect 186 186 189 189 
rect 186 189 189 192 
rect 186 192 189 195 
rect 186 195 189 198 
rect 186 198 189 201 
rect 186 201 189 204 
rect 186 204 189 207 
rect 186 207 189 210 
rect 186 210 189 213 
rect 186 213 189 216 
rect 186 216 189 219 
rect 186 219 189 222 
rect 186 222 189 225 
rect 186 225 189 228 
rect 186 228 189 231 
rect 186 231 189 234 
rect 186 234 189 237 
rect 186 237 189 240 
rect 186 240 189 243 
rect 186 243 189 246 
rect 186 246 189 249 
rect 186 249 189 252 
rect 186 252 189 255 
rect 186 255 189 258 
rect 186 258 189 261 
rect 186 261 189 264 
rect 186 264 189 267 
rect 186 267 189 270 
rect 186 270 189 273 
rect 186 273 189 276 
rect 186 276 189 279 
rect 186 279 189 282 
rect 186 282 189 285 
rect 186 285 189 288 
rect 186 288 189 291 
rect 186 291 189 294 
rect 186 294 189 297 
rect 186 297 189 300 
rect 186 300 189 303 
rect 186 303 189 306 
rect 186 306 189 309 
rect 186 309 189 312 
rect 186 312 189 315 
rect 186 315 189 318 
rect 186 318 189 321 
rect 186 321 189 324 
rect 186 324 189 327 
rect 186 327 189 330 
rect 186 330 189 333 
rect 186 333 189 336 
rect 186 336 189 339 
rect 186 339 189 342 
rect 186 342 189 345 
rect 186 345 189 348 
rect 186 348 189 351 
rect 186 351 189 354 
rect 186 354 189 357 
rect 186 357 189 360 
rect 186 360 189 363 
rect 186 363 189 366 
rect 186 366 189 369 
rect 186 369 189 372 
rect 186 372 189 375 
rect 186 375 189 378 
rect 186 378 189 381 
rect 186 381 189 384 
rect 186 384 189 387 
rect 186 387 189 390 
rect 186 390 189 393 
rect 186 393 189 396 
rect 186 396 189 399 
rect 186 399 189 402 
rect 186 402 189 405 
rect 186 405 189 408 
rect 186 408 189 411 
rect 186 411 189 414 
rect 186 414 189 417 
rect 186 417 189 420 
rect 186 420 189 423 
rect 186 423 189 426 
rect 186 426 189 429 
rect 186 429 189 432 
rect 186 432 189 435 
rect 186 435 189 438 
rect 186 438 189 441 
rect 186 441 189 444 
rect 186 444 189 447 
rect 186 447 189 450 
rect 186 450 189 453 
rect 186 453 189 456 
rect 186 456 189 459 
rect 186 459 189 462 
rect 186 462 189 465 
rect 186 465 189 468 
rect 186 468 189 471 
rect 186 471 189 474 
rect 186 474 189 477 
rect 186 477 189 480 
rect 186 480 189 483 
rect 186 483 189 486 
rect 186 486 189 489 
rect 186 489 189 492 
rect 186 492 189 495 
rect 186 495 189 498 
rect 186 498 189 501 
rect 186 501 189 504 
rect 186 504 189 507 
rect 186 507 189 510 
rect 189 0 192 3 
rect 189 3 192 6 
rect 189 6 192 9 
rect 189 9 192 12 
rect 189 12 192 15 
rect 189 15 192 18 
rect 189 18 192 21 
rect 189 21 192 24 
rect 189 24 192 27 
rect 189 27 192 30 
rect 189 30 192 33 
rect 189 33 192 36 
rect 189 36 192 39 
rect 189 39 192 42 
rect 189 42 192 45 
rect 189 45 192 48 
rect 189 48 192 51 
rect 189 51 192 54 
rect 189 54 192 57 
rect 189 57 192 60 
rect 189 60 192 63 
rect 189 63 192 66 
rect 189 66 192 69 
rect 189 69 192 72 
rect 189 72 192 75 
rect 189 75 192 78 
rect 189 78 192 81 
rect 189 81 192 84 
rect 189 84 192 87 
rect 189 87 192 90 
rect 189 90 192 93 
rect 189 93 192 96 
rect 189 96 192 99 
rect 189 99 192 102 
rect 189 102 192 105 
rect 189 105 192 108 
rect 189 108 192 111 
rect 189 111 192 114 
rect 189 114 192 117 
rect 189 117 192 120 
rect 189 120 192 123 
rect 189 123 192 126 
rect 189 126 192 129 
rect 189 129 192 132 
rect 189 132 192 135 
rect 189 135 192 138 
rect 189 138 192 141 
rect 189 141 192 144 
rect 189 144 192 147 
rect 189 147 192 150 
rect 189 150 192 153 
rect 189 153 192 156 
rect 189 156 192 159 
rect 189 159 192 162 
rect 189 162 192 165 
rect 189 165 192 168 
rect 189 168 192 171 
rect 189 171 192 174 
rect 189 174 192 177 
rect 189 177 192 180 
rect 189 180 192 183 
rect 189 183 192 186 
rect 189 186 192 189 
rect 189 189 192 192 
rect 189 192 192 195 
rect 189 195 192 198 
rect 189 198 192 201 
rect 189 201 192 204 
rect 189 204 192 207 
rect 189 207 192 210 
rect 189 210 192 213 
rect 189 213 192 216 
rect 189 216 192 219 
rect 189 219 192 222 
rect 189 222 192 225 
rect 189 225 192 228 
rect 189 228 192 231 
rect 189 231 192 234 
rect 189 234 192 237 
rect 189 237 192 240 
rect 189 240 192 243 
rect 189 243 192 246 
rect 189 246 192 249 
rect 189 249 192 252 
rect 189 252 192 255 
rect 189 255 192 258 
rect 189 258 192 261 
rect 189 261 192 264 
rect 189 264 192 267 
rect 189 267 192 270 
rect 189 270 192 273 
rect 189 273 192 276 
rect 189 276 192 279 
rect 189 279 192 282 
rect 189 282 192 285 
rect 189 285 192 288 
rect 189 288 192 291 
rect 189 291 192 294 
rect 189 294 192 297 
rect 189 297 192 300 
rect 189 300 192 303 
rect 189 303 192 306 
rect 189 306 192 309 
rect 189 309 192 312 
rect 189 312 192 315 
rect 189 315 192 318 
rect 189 318 192 321 
rect 189 321 192 324 
rect 189 324 192 327 
rect 189 327 192 330 
rect 189 330 192 333 
rect 189 333 192 336 
rect 189 336 192 339 
rect 189 339 192 342 
rect 189 342 192 345 
rect 189 345 192 348 
rect 189 348 192 351 
rect 189 351 192 354 
rect 189 354 192 357 
rect 189 357 192 360 
rect 189 360 192 363 
rect 189 363 192 366 
rect 189 366 192 369 
rect 189 369 192 372 
rect 189 372 192 375 
rect 189 375 192 378 
rect 189 378 192 381 
rect 189 381 192 384 
rect 189 384 192 387 
rect 189 387 192 390 
rect 189 390 192 393 
rect 189 393 192 396 
rect 189 396 192 399 
rect 189 399 192 402 
rect 189 402 192 405 
rect 189 405 192 408 
rect 189 408 192 411 
rect 189 411 192 414 
rect 189 414 192 417 
rect 189 417 192 420 
rect 189 420 192 423 
rect 189 423 192 426 
rect 189 426 192 429 
rect 189 429 192 432 
rect 189 432 192 435 
rect 189 435 192 438 
rect 189 438 192 441 
rect 189 441 192 444 
rect 189 444 192 447 
rect 189 447 192 450 
rect 189 450 192 453 
rect 189 453 192 456 
rect 189 456 192 459 
rect 189 459 192 462 
rect 189 462 192 465 
rect 189 465 192 468 
rect 189 468 192 471 
rect 189 471 192 474 
rect 189 474 192 477 
rect 189 477 192 480 
rect 189 480 192 483 
rect 189 483 192 486 
rect 189 486 192 489 
rect 189 489 192 492 
rect 189 492 192 495 
rect 189 495 192 498 
rect 189 498 192 501 
rect 189 501 192 504 
rect 189 504 192 507 
rect 189 507 192 510 
rect 192 0 195 3 
rect 192 3 195 6 
rect 192 6 195 9 
rect 192 9 195 12 
rect 192 12 195 15 
rect 192 15 195 18 
rect 192 18 195 21 
rect 192 21 195 24 
rect 192 24 195 27 
rect 192 27 195 30 
rect 192 30 195 33 
rect 192 33 195 36 
rect 192 36 195 39 
rect 192 39 195 42 
rect 192 42 195 45 
rect 192 45 195 48 
rect 192 48 195 51 
rect 192 51 195 54 
rect 192 54 195 57 
rect 192 57 195 60 
rect 192 60 195 63 
rect 192 63 195 66 
rect 192 66 195 69 
rect 192 69 195 72 
rect 192 72 195 75 
rect 192 75 195 78 
rect 192 78 195 81 
rect 192 81 195 84 
rect 192 84 195 87 
rect 192 87 195 90 
rect 192 90 195 93 
rect 192 93 195 96 
rect 192 96 195 99 
rect 192 99 195 102 
rect 192 102 195 105 
rect 192 105 195 108 
rect 192 108 195 111 
rect 192 111 195 114 
rect 192 114 195 117 
rect 192 117 195 120 
rect 192 120 195 123 
rect 192 123 195 126 
rect 192 126 195 129 
rect 192 129 195 132 
rect 192 132 195 135 
rect 192 135 195 138 
rect 192 138 195 141 
rect 192 141 195 144 
rect 192 144 195 147 
rect 192 147 195 150 
rect 192 150 195 153 
rect 192 153 195 156 
rect 192 156 195 159 
rect 192 159 195 162 
rect 192 162 195 165 
rect 192 165 195 168 
rect 192 168 195 171 
rect 192 171 195 174 
rect 192 174 195 177 
rect 192 177 195 180 
rect 192 180 195 183 
rect 192 183 195 186 
rect 192 186 195 189 
rect 192 189 195 192 
rect 192 192 195 195 
rect 192 195 195 198 
rect 192 198 195 201 
rect 192 201 195 204 
rect 192 204 195 207 
rect 192 207 195 210 
rect 192 210 195 213 
rect 192 213 195 216 
rect 192 216 195 219 
rect 192 219 195 222 
rect 192 222 195 225 
rect 192 225 195 228 
rect 192 228 195 231 
rect 192 231 195 234 
rect 192 234 195 237 
rect 192 237 195 240 
rect 192 240 195 243 
rect 192 243 195 246 
rect 192 246 195 249 
rect 192 249 195 252 
rect 192 252 195 255 
rect 192 255 195 258 
rect 192 258 195 261 
rect 192 261 195 264 
rect 192 264 195 267 
rect 192 267 195 270 
rect 192 270 195 273 
rect 192 273 195 276 
rect 192 276 195 279 
rect 192 279 195 282 
rect 192 282 195 285 
rect 192 285 195 288 
rect 192 288 195 291 
rect 192 291 195 294 
rect 192 294 195 297 
rect 192 297 195 300 
rect 192 300 195 303 
rect 192 303 195 306 
rect 192 306 195 309 
rect 192 309 195 312 
rect 192 312 195 315 
rect 192 315 195 318 
rect 192 318 195 321 
rect 192 321 195 324 
rect 192 324 195 327 
rect 192 327 195 330 
rect 192 330 195 333 
rect 192 333 195 336 
rect 192 336 195 339 
rect 192 339 195 342 
rect 192 342 195 345 
rect 192 345 195 348 
rect 192 348 195 351 
rect 192 351 195 354 
rect 192 354 195 357 
rect 192 357 195 360 
rect 192 360 195 363 
rect 192 363 195 366 
rect 192 366 195 369 
rect 192 369 195 372 
rect 192 372 195 375 
rect 192 375 195 378 
rect 192 378 195 381 
rect 192 381 195 384 
rect 192 384 195 387 
rect 192 387 195 390 
rect 192 390 195 393 
rect 192 393 195 396 
rect 192 396 195 399 
rect 192 399 195 402 
rect 192 402 195 405 
rect 192 405 195 408 
rect 192 408 195 411 
rect 192 411 195 414 
rect 192 414 195 417 
rect 192 417 195 420 
rect 192 420 195 423 
rect 192 423 195 426 
rect 192 426 195 429 
rect 192 429 195 432 
rect 192 432 195 435 
rect 192 435 195 438 
rect 192 438 195 441 
rect 192 441 195 444 
rect 192 444 195 447 
rect 192 447 195 450 
rect 192 450 195 453 
rect 192 453 195 456 
rect 192 456 195 459 
rect 192 459 195 462 
rect 192 462 195 465 
rect 192 465 195 468 
rect 192 468 195 471 
rect 192 471 195 474 
rect 192 474 195 477 
rect 192 477 195 480 
rect 192 480 195 483 
rect 192 483 195 486 
rect 192 486 195 489 
rect 192 489 195 492 
rect 192 492 195 495 
rect 192 495 195 498 
rect 192 498 195 501 
rect 192 501 195 504 
rect 192 504 195 507 
rect 192 507 195 510 
rect 195 0 198 3 
rect 195 3 198 6 
rect 195 6 198 9 
rect 195 9 198 12 
rect 195 12 198 15 
rect 195 15 198 18 
rect 195 18 198 21 
rect 195 21 198 24 
rect 195 24 198 27 
rect 195 27 198 30 
rect 195 30 198 33 
rect 195 33 198 36 
rect 195 36 198 39 
rect 195 39 198 42 
rect 195 42 198 45 
rect 195 45 198 48 
rect 195 48 198 51 
rect 195 51 198 54 
rect 195 54 198 57 
rect 195 57 198 60 
rect 195 60 198 63 
rect 195 63 198 66 
rect 195 66 198 69 
rect 195 69 198 72 
rect 195 72 198 75 
rect 195 75 198 78 
rect 195 78 198 81 
rect 195 81 198 84 
rect 195 84 198 87 
rect 195 87 198 90 
rect 195 90 198 93 
rect 195 93 198 96 
rect 195 96 198 99 
rect 195 99 198 102 
rect 195 102 198 105 
rect 195 105 198 108 
rect 195 108 198 111 
rect 195 111 198 114 
rect 195 114 198 117 
rect 195 117 198 120 
rect 195 120 198 123 
rect 195 123 198 126 
rect 195 126 198 129 
rect 195 129 198 132 
rect 195 132 198 135 
rect 195 135 198 138 
rect 195 138 198 141 
rect 195 141 198 144 
rect 195 144 198 147 
rect 195 147 198 150 
rect 195 150 198 153 
rect 195 153 198 156 
rect 195 156 198 159 
rect 195 159 198 162 
rect 195 162 198 165 
rect 195 165 198 168 
rect 195 168 198 171 
rect 195 171 198 174 
rect 195 174 198 177 
rect 195 177 198 180 
rect 195 180 198 183 
rect 195 183 198 186 
rect 195 186 198 189 
rect 195 189 198 192 
rect 195 192 198 195 
rect 195 195 198 198 
rect 195 198 198 201 
rect 195 201 198 204 
rect 195 204 198 207 
rect 195 207 198 210 
rect 195 210 198 213 
rect 195 213 198 216 
rect 195 216 198 219 
rect 195 219 198 222 
rect 195 222 198 225 
rect 195 225 198 228 
rect 195 228 198 231 
rect 195 231 198 234 
rect 195 234 198 237 
rect 195 237 198 240 
rect 195 240 198 243 
rect 195 243 198 246 
rect 195 246 198 249 
rect 195 249 198 252 
rect 195 252 198 255 
rect 195 255 198 258 
rect 195 258 198 261 
rect 195 261 198 264 
rect 195 264 198 267 
rect 195 267 198 270 
rect 195 270 198 273 
rect 195 273 198 276 
rect 195 276 198 279 
rect 195 279 198 282 
rect 195 282 198 285 
rect 195 285 198 288 
rect 195 288 198 291 
rect 195 291 198 294 
rect 195 294 198 297 
rect 195 297 198 300 
rect 195 300 198 303 
rect 195 303 198 306 
rect 195 306 198 309 
rect 195 309 198 312 
rect 195 312 198 315 
rect 195 315 198 318 
rect 195 318 198 321 
rect 195 321 198 324 
rect 195 324 198 327 
rect 195 327 198 330 
rect 195 330 198 333 
rect 195 333 198 336 
rect 195 336 198 339 
rect 195 339 198 342 
rect 195 342 198 345 
rect 195 345 198 348 
rect 195 348 198 351 
rect 195 351 198 354 
rect 195 354 198 357 
rect 195 357 198 360 
rect 195 360 198 363 
rect 195 363 198 366 
rect 195 366 198 369 
rect 195 369 198 372 
rect 195 372 198 375 
rect 195 375 198 378 
rect 195 378 198 381 
rect 195 381 198 384 
rect 195 384 198 387 
rect 195 387 198 390 
rect 195 390 198 393 
rect 195 393 198 396 
rect 195 396 198 399 
rect 195 399 198 402 
rect 195 402 198 405 
rect 195 405 198 408 
rect 195 408 198 411 
rect 195 411 198 414 
rect 195 414 198 417 
rect 195 417 198 420 
rect 195 420 198 423 
rect 195 423 198 426 
rect 195 426 198 429 
rect 195 429 198 432 
rect 195 432 198 435 
rect 195 435 198 438 
rect 195 438 198 441 
rect 195 441 198 444 
rect 195 444 198 447 
rect 195 447 198 450 
rect 195 450 198 453 
rect 195 453 198 456 
rect 195 456 198 459 
rect 195 459 198 462 
rect 195 462 198 465 
rect 195 465 198 468 
rect 195 468 198 471 
rect 195 471 198 474 
rect 195 474 198 477 
rect 195 477 198 480 
rect 195 480 198 483 
rect 195 483 198 486 
rect 195 486 198 489 
rect 195 489 198 492 
rect 195 492 198 495 
rect 195 495 198 498 
rect 195 498 198 501 
rect 195 501 198 504 
rect 195 504 198 507 
rect 195 507 198 510 
rect 198 0 201 3 
rect 198 3 201 6 
rect 198 6 201 9 
rect 198 9 201 12 
rect 198 12 201 15 
rect 198 15 201 18 
rect 198 18 201 21 
rect 198 21 201 24 
rect 198 24 201 27 
rect 198 27 201 30 
rect 198 30 201 33 
rect 198 33 201 36 
rect 198 36 201 39 
rect 198 39 201 42 
rect 198 42 201 45 
rect 198 45 201 48 
rect 198 48 201 51 
rect 198 51 201 54 
rect 198 54 201 57 
rect 198 57 201 60 
rect 198 60 201 63 
rect 198 63 201 66 
rect 198 66 201 69 
rect 198 69 201 72 
rect 198 72 201 75 
rect 198 75 201 78 
rect 198 78 201 81 
rect 198 81 201 84 
rect 198 84 201 87 
rect 198 87 201 90 
rect 198 90 201 93 
rect 198 93 201 96 
rect 198 96 201 99 
rect 198 99 201 102 
rect 198 102 201 105 
rect 198 105 201 108 
rect 198 108 201 111 
rect 198 111 201 114 
rect 198 114 201 117 
rect 198 117 201 120 
rect 198 120 201 123 
rect 198 123 201 126 
rect 198 126 201 129 
rect 198 129 201 132 
rect 198 132 201 135 
rect 198 135 201 138 
rect 198 138 201 141 
rect 198 141 201 144 
rect 198 144 201 147 
rect 198 147 201 150 
rect 198 150 201 153 
rect 198 153 201 156 
rect 198 156 201 159 
rect 198 159 201 162 
rect 198 162 201 165 
rect 198 165 201 168 
rect 198 168 201 171 
rect 198 171 201 174 
rect 198 174 201 177 
rect 198 177 201 180 
rect 198 180 201 183 
rect 198 183 201 186 
rect 198 186 201 189 
rect 198 189 201 192 
rect 198 192 201 195 
rect 198 195 201 198 
rect 198 198 201 201 
rect 198 201 201 204 
rect 198 204 201 207 
rect 198 207 201 210 
rect 198 210 201 213 
rect 198 213 201 216 
rect 198 216 201 219 
rect 198 219 201 222 
rect 198 222 201 225 
rect 198 225 201 228 
rect 198 228 201 231 
rect 198 231 201 234 
rect 198 234 201 237 
rect 198 237 201 240 
rect 198 240 201 243 
rect 198 243 201 246 
rect 198 246 201 249 
rect 198 249 201 252 
rect 198 252 201 255 
rect 198 255 201 258 
rect 198 258 201 261 
rect 198 261 201 264 
rect 198 264 201 267 
rect 198 267 201 270 
rect 198 270 201 273 
rect 198 273 201 276 
rect 198 276 201 279 
rect 198 279 201 282 
rect 198 282 201 285 
rect 198 285 201 288 
rect 198 288 201 291 
rect 198 291 201 294 
rect 198 294 201 297 
rect 198 297 201 300 
rect 198 300 201 303 
rect 198 303 201 306 
rect 198 306 201 309 
rect 198 309 201 312 
rect 198 312 201 315 
rect 198 315 201 318 
rect 198 318 201 321 
rect 198 321 201 324 
rect 198 324 201 327 
rect 198 327 201 330 
rect 198 330 201 333 
rect 198 333 201 336 
rect 198 336 201 339 
rect 198 339 201 342 
rect 198 342 201 345 
rect 198 345 201 348 
rect 198 348 201 351 
rect 198 351 201 354 
rect 198 354 201 357 
rect 198 357 201 360 
rect 198 360 201 363 
rect 198 363 201 366 
rect 198 366 201 369 
rect 198 369 201 372 
rect 198 372 201 375 
rect 198 375 201 378 
rect 198 378 201 381 
rect 198 381 201 384 
rect 198 384 201 387 
rect 198 387 201 390 
rect 198 390 201 393 
rect 198 393 201 396 
rect 198 396 201 399 
rect 198 399 201 402 
rect 198 402 201 405 
rect 198 405 201 408 
rect 198 408 201 411 
rect 198 411 201 414 
rect 198 414 201 417 
rect 198 417 201 420 
rect 198 420 201 423 
rect 198 423 201 426 
rect 198 426 201 429 
rect 198 429 201 432 
rect 198 432 201 435 
rect 198 435 201 438 
rect 198 438 201 441 
rect 198 441 201 444 
rect 198 444 201 447 
rect 198 447 201 450 
rect 198 450 201 453 
rect 198 453 201 456 
rect 198 456 201 459 
rect 198 459 201 462 
rect 198 462 201 465 
rect 198 465 201 468 
rect 198 468 201 471 
rect 198 471 201 474 
rect 198 474 201 477 
rect 198 477 201 480 
rect 198 480 201 483 
rect 198 483 201 486 
rect 198 486 201 489 
rect 198 489 201 492 
rect 198 492 201 495 
rect 198 495 201 498 
rect 198 498 201 501 
rect 198 501 201 504 
rect 198 504 201 507 
rect 198 507 201 510 
rect 201 0 204 3 
rect 201 3 204 6 
rect 201 6 204 9 
rect 201 9 204 12 
rect 201 12 204 15 
rect 201 15 204 18 
rect 201 18 204 21 
rect 201 21 204 24 
rect 201 24 204 27 
rect 201 27 204 30 
rect 201 30 204 33 
rect 201 33 204 36 
rect 201 36 204 39 
rect 201 39 204 42 
rect 201 42 204 45 
rect 201 45 204 48 
rect 201 48 204 51 
rect 201 51 204 54 
rect 201 54 204 57 
rect 201 57 204 60 
rect 201 60 204 63 
rect 201 63 204 66 
rect 201 66 204 69 
rect 201 69 204 72 
rect 201 72 204 75 
rect 201 75 204 78 
rect 201 78 204 81 
rect 201 81 204 84 
rect 201 84 204 87 
rect 201 87 204 90 
rect 201 90 204 93 
rect 201 93 204 96 
rect 201 96 204 99 
rect 201 99 204 102 
rect 201 102 204 105 
rect 201 105 204 108 
rect 201 108 204 111 
rect 201 111 204 114 
rect 201 114 204 117 
rect 201 117 204 120 
rect 201 120 204 123 
rect 201 123 204 126 
rect 201 126 204 129 
rect 201 129 204 132 
rect 201 132 204 135 
rect 201 135 204 138 
rect 201 138 204 141 
rect 201 141 204 144 
rect 201 144 204 147 
rect 201 147 204 150 
rect 201 150 204 153 
rect 201 153 204 156 
rect 201 156 204 159 
rect 201 159 204 162 
rect 201 162 204 165 
rect 201 165 204 168 
rect 201 168 204 171 
rect 201 171 204 174 
rect 201 174 204 177 
rect 201 177 204 180 
rect 201 180 204 183 
rect 201 183 204 186 
rect 201 186 204 189 
rect 201 189 204 192 
rect 201 192 204 195 
rect 201 195 204 198 
rect 201 198 204 201 
rect 201 201 204 204 
rect 201 204 204 207 
rect 201 207 204 210 
rect 201 210 204 213 
rect 201 213 204 216 
rect 201 216 204 219 
rect 201 219 204 222 
rect 201 222 204 225 
rect 201 225 204 228 
rect 201 228 204 231 
rect 201 231 204 234 
rect 201 234 204 237 
rect 201 237 204 240 
rect 201 240 204 243 
rect 201 243 204 246 
rect 201 246 204 249 
rect 201 249 204 252 
rect 201 252 204 255 
rect 201 255 204 258 
rect 201 258 204 261 
rect 201 261 204 264 
rect 201 264 204 267 
rect 201 267 204 270 
rect 201 270 204 273 
rect 201 273 204 276 
rect 201 276 204 279 
rect 201 279 204 282 
rect 201 282 204 285 
rect 201 285 204 288 
rect 201 288 204 291 
rect 201 291 204 294 
rect 201 294 204 297 
rect 201 297 204 300 
rect 201 300 204 303 
rect 201 303 204 306 
rect 201 306 204 309 
rect 201 309 204 312 
rect 201 312 204 315 
rect 201 315 204 318 
rect 201 318 204 321 
rect 201 321 204 324 
rect 201 324 204 327 
rect 201 327 204 330 
rect 201 330 204 333 
rect 201 333 204 336 
rect 201 336 204 339 
rect 201 339 204 342 
rect 201 342 204 345 
rect 201 345 204 348 
rect 201 348 204 351 
rect 201 351 204 354 
rect 201 354 204 357 
rect 201 357 204 360 
rect 201 360 204 363 
rect 201 363 204 366 
rect 201 366 204 369 
rect 201 369 204 372 
rect 201 372 204 375 
rect 201 375 204 378 
rect 201 378 204 381 
rect 201 381 204 384 
rect 201 384 204 387 
rect 201 387 204 390 
rect 201 390 204 393 
rect 201 393 204 396 
rect 201 396 204 399 
rect 201 399 204 402 
rect 201 402 204 405 
rect 201 405 204 408 
rect 201 408 204 411 
rect 201 411 204 414 
rect 201 414 204 417 
rect 201 417 204 420 
rect 201 420 204 423 
rect 201 423 204 426 
rect 201 426 204 429 
rect 201 429 204 432 
rect 201 432 204 435 
rect 201 435 204 438 
rect 201 438 204 441 
rect 201 441 204 444 
rect 201 444 204 447 
rect 201 447 204 450 
rect 201 450 204 453 
rect 201 453 204 456 
rect 201 456 204 459 
rect 201 459 204 462 
rect 201 462 204 465 
rect 201 465 204 468 
rect 201 468 204 471 
rect 201 471 204 474 
rect 201 474 204 477 
rect 201 477 204 480 
rect 201 480 204 483 
rect 201 483 204 486 
rect 201 486 204 489 
rect 201 489 204 492 
rect 201 492 204 495 
rect 201 495 204 498 
rect 201 498 204 501 
rect 201 501 204 504 
rect 201 504 204 507 
rect 201 507 204 510 
rect 204 0 207 3 
rect 204 3 207 6 
rect 204 6 207 9 
rect 204 9 207 12 
rect 204 12 207 15 
rect 204 15 207 18 
rect 204 18 207 21 
rect 204 21 207 24 
rect 204 24 207 27 
rect 204 27 207 30 
rect 204 30 207 33 
rect 204 33 207 36 
rect 204 36 207 39 
rect 204 39 207 42 
rect 204 42 207 45 
rect 204 45 207 48 
rect 204 48 207 51 
rect 204 51 207 54 
rect 204 54 207 57 
rect 204 57 207 60 
rect 204 60 207 63 
rect 204 63 207 66 
rect 204 66 207 69 
rect 204 69 207 72 
rect 204 72 207 75 
rect 204 75 207 78 
rect 204 78 207 81 
rect 204 81 207 84 
rect 204 84 207 87 
rect 204 87 207 90 
rect 204 90 207 93 
rect 204 93 207 96 
rect 204 96 207 99 
rect 204 99 207 102 
rect 204 102 207 105 
rect 204 105 207 108 
rect 204 108 207 111 
rect 204 111 207 114 
rect 204 114 207 117 
rect 204 117 207 120 
rect 204 120 207 123 
rect 204 123 207 126 
rect 204 126 207 129 
rect 204 129 207 132 
rect 204 132 207 135 
rect 204 135 207 138 
rect 204 138 207 141 
rect 204 141 207 144 
rect 204 144 207 147 
rect 204 147 207 150 
rect 204 150 207 153 
rect 204 153 207 156 
rect 204 156 207 159 
rect 204 159 207 162 
rect 204 162 207 165 
rect 204 165 207 168 
rect 204 168 207 171 
rect 204 171 207 174 
rect 204 174 207 177 
rect 204 177 207 180 
rect 204 180 207 183 
rect 204 183 207 186 
rect 204 186 207 189 
rect 204 189 207 192 
rect 204 192 207 195 
rect 204 195 207 198 
rect 204 198 207 201 
rect 204 201 207 204 
rect 204 204 207 207 
rect 204 207 207 210 
rect 204 210 207 213 
rect 204 213 207 216 
rect 204 216 207 219 
rect 204 219 207 222 
rect 204 222 207 225 
rect 204 225 207 228 
rect 204 228 207 231 
rect 204 231 207 234 
rect 204 234 207 237 
rect 204 237 207 240 
rect 204 240 207 243 
rect 204 243 207 246 
rect 204 246 207 249 
rect 204 249 207 252 
rect 204 252 207 255 
rect 204 255 207 258 
rect 204 258 207 261 
rect 204 261 207 264 
rect 204 264 207 267 
rect 204 267 207 270 
rect 204 270 207 273 
rect 204 273 207 276 
rect 204 276 207 279 
rect 204 279 207 282 
rect 204 282 207 285 
rect 204 285 207 288 
rect 204 288 207 291 
rect 204 291 207 294 
rect 204 294 207 297 
rect 204 297 207 300 
rect 204 300 207 303 
rect 204 303 207 306 
rect 204 306 207 309 
rect 204 309 207 312 
rect 204 312 207 315 
rect 204 315 207 318 
rect 204 318 207 321 
rect 204 321 207 324 
rect 204 324 207 327 
rect 204 327 207 330 
rect 204 330 207 333 
rect 204 333 207 336 
rect 204 336 207 339 
rect 204 339 207 342 
rect 204 342 207 345 
rect 204 345 207 348 
rect 204 348 207 351 
rect 204 351 207 354 
rect 204 354 207 357 
rect 204 357 207 360 
rect 204 360 207 363 
rect 204 363 207 366 
rect 204 366 207 369 
rect 204 369 207 372 
rect 204 372 207 375 
rect 204 375 207 378 
rect 204 378 207 381 
rect 204 381 207 384 
rect 204 384 207 387 
rect 204 387 207 390 
rect 204 390 207 393 
rect 204 393 207 396 
rect 204 396 207 399 
rect 204 399 207 402 
rect 204 402 207 405 
rect 204 405 207 408 
rect 204 408 207 411 
rect 204 411 207 414 
rect 204 414 207 417 
rect 204 417 207 420 
rect 204 420 207 423 
rect 204 423 207 426 
rect 204 426 207 429 
rect 204 429 207 432 
rect 204 432 207 435 
rect 204 435 207 438 
rect 204 438 207 441 
rect 204 441 207 444 
rect 204 444 207 447 
rect 204 447 207 450 
rect 204 450 207 453 
rect 204 453 207 456 
rect 204 456 207 459 
rect 204 459 207 462 
rect 204 462 207 465 
rect 204 465 207 468 
rect 204 468 207 471 
rect 204 471 207 474 
rect 204 474 207 477 
rect 204 477 207 480 
rect 204 480 207 483 
rect 204 483 207 486 
rect 204 486 207 489 
rect 204 489 207 492 
rect 204 492 207 495 
rect 204 495 207 498 
rect 204 498 207 501 
rect 204 501 207 504 
rect 204 504 207 507 
rect 204 507 207 510 
rect 207 0 210 3 
rect 207 3 210 6 
rect 207 6 210 9 
rect 207 9 210 12 
rect 207 12 210 15 
rect 207 15 210 18 
rect 207 18 210 21 
rect 207 21 210 24 
rect 207 24 210 27 
rect 207 27 210 30 
rect 207 30 210 33 
rect 207 33 210 36 
rect 207 36 210 39 
rect 207 39 210 42 
rect 207 42 210 45 
rect 207 45 210 48 
rect 207 48 210 51 
rect 207 51 210 54 
rect 207 54 210 57 
rect 207 57 210 60 
rect 207 60 210 63 
rect 207 63 210 66 
rect 207 66 210 69 
rect 207 69 210 72 
rect 207 72 210 75 
rect 207 75 210 78 
rect 207 78 210 81 
rect 207 81 210 84 
rect 207 84 210 87 
rect 207 87 210 90 
rect 207 90 210 93 
rect 207 93 210 96 
rect 207 96 210 99 
rect 207 99 210 102 
rect 207 102 210 105 
rect 207 105 210 108 
rect 207 108 210 111 
rect 207 111 210 114 
rect 207 114 210 117 
rect 207 117 210 120 
rect 207 120 210 123 
rect 207 123 210 126 
rect 207 126 210 129 
rect 207 129 210 132 
rect 207 132 210 135 
rect 207 135 210 138 
rect 207 138 210 141 
rect 207 141 210 144 
rect 207 144 210 147 
rect 207 147 210 150 
rect 207 150 210 153 
rect 207 153 210 156 
rect 207 156 210 159 
rect 207 159 210 162 
rect 207 162 210 165 
rect 207 165 210 168 
rect 207 168 210 171 
rect 207 171 210 174 
rect 207 174 210 177 
rect 207 177 210 180 
rect 207 180 210 183 
rect 207 183 210 186 
rect 207 186 210 189 
rect 207 189 210 192 
rect 207 192 210 195 
rect 207 195 210 198 
rect 207 198 210 201 
rect 207 201 210 204 
rect 207 204 210 207 
rect 207 207 210 210 
rect 207 210 210 213 
rect 207 213 210 216 
rect 207 216 210 219 
rect 207 219 210 222 
rect 207 222 210 225 
rect 207 225 210 228 
rect 207 228 210 231 
rect 207 231 210 234 
rect 207 234 210 237 
rect 207 237 210 240 
rect 207 240 210 243 
rect 207 243 210 246 
rect 207 246 210 249 
rect 207 249 210 252 
rect 207 252 210 255 
rect 207 255 210 258 
rect 207 258 210 261 
rect 207 261 210 264 
rect 207 264 210 267 
rect 207 267 210 270 
rect 207 270 210 273 
rect 207 273 210 276 
rect 207 276 210 279 
rect 207 279 210 282 
rect 207 282 210 285 
rect 207 285 210 288 
rect 207 288 210 291 
rect 207 291 210 294 
rect 207 294 210 297 
rect 207 297 210 300 
rect 207 300 210 303 
rect 207 303 210 306 
rect 207 306 210 309 
rect 207 309 210 312 
rect 207 312 210 315 
rect 207 315 210 318 
rect 207 318 210 321 
rect 207 321 210 324 
rect 207 324 210 327 
rect 207 327 210 330 
rect 207 330 210 333 
rect 207 333 210 336 
rect 207 336 210 339 
rect 207 339 210 342 
rect 207 342 210 345 
rect 207 345 210 348 
rect 207 348 210 351 
rect 207 351 210 354 
rect 207 354 210 357 
rect 207 357 210 360 
rect 207 360 210 363 
rect 207 363 210 366 
rect 207 366 210 369 
rect 207 369 210 372 
rect 207 372 210 375 
rect 207 375 210 378 
rect 207 378 210 381 
rect 207 381 210 384 
rect 207 384 210 387 
rect 207 387 210 390 
rect 207 390 210 393 
rect 207 393 210 396 
rect 207 396 210 399 
rect 207 399 210 402 
rect 207 402 210 405 
rect 207 405 210 408 
rect 207 408 210 411 
rect 207 411 210 414 
rect 207 414 210 417 
rect 207 417 210 420 
rect 207 420 210 423 
rect 207 423 210 426 
rect 207 426 210 429 
rect 207 429 210 432 
rect 207 432 210 435 
rect 207 435 210 438 
rect 207 438 210 441 
rect 207 441 210 444 
rect 207 444 210 447 
rect 207 447 210 450 
rect 207 450 210 453 
rect 207 453 210 456 
rect 207 456 210 459 
rect 207 459 210 462 
rect 207 462 210 465 
rect 207 465 210 468 
rect 207 468 210 471 
rect 207 471 210 474 
rect 207 474 210 477 
rect 207 477 210 480 
rect 207 480 210 483 
rect 207 483 210 486 
rect 207 486 210 489 
rect 207 489 210 492 
rect 207 492 210 495 
rect 207 495 210 498 
rect 207 498 210 501 
rect 207 501 210 504 
rect 207 504 210 507 
rect 207 507 210 510 
rect 210 0 213 3 
rect 210 3 213 6 
rect 210 6 213 9 
rect 210 9 213 12 
rect 210 12 213 15 
rect 210 15 213 18 
rect 210 18 213 21 
rect 210 21 213 24 
rect 210 24 213 27 
rect 210 27 213 30 
rect 210 30 213 33 
rect 210 33 213 36 
rect 210 36 213 39 
rect 210 39 213 42 
rect 210 42 213 45 
rect 210 45 213 48 
rect 210 48 213 51 
rect 210 51 213 54 
rect 210 54 213 57 
rect 210 57 213 60 
rect 210 60 213 63 
rect 210 63 213 66 
rect 210 66 213 69 
rect 210 69 213 72 
rect 210 72 213 75 
rect 210 75 213 78 
rect 210 78 213 81 
rect 210 81 213 84 
rect 210 84 213 87 
rect 210 87 213 90 
rect 210 90 213 93 
rect 210 93 213 96 
rect 210 96 213 99 
rect 210 99 213 102 
rect 210 102 213 105 
rect 210 105 213 108 
rect 210 108 213 111 
rect 210 111 213 114 
rect 210 114 213 117 
rect 210 117 213 120 
rect 210 120 213 123 
rect 210 123 213 126 
rect 210 126 213 129 
rect 210 129 213 132 
rect 210 132 213 135 
rect 210 135 213 138 
rect 210 138 213 141 
rect 210 141 213 144 
rect 210 144 213 147 
rect 210 147 213 150 
rect 210 150 213 153 
rect 210 153 213 156 
rect 210 156 213 159 
rect 210 159 213 162 
rect 210 162 213 165 
rect 210 165 213 168 
rect 210 168 213 171 
rect 210 171 213 174 
rect 210 174 213 177 
rect 210 177 213 180 
rect 210 180 213 183 
rect 210 183 213 186 
rect 210 186 213 189 
rect 210 189 213 192 
rect 210 192 213 195 
rect 210 195 213 198 
rect 210 198 213 201 
rect 210 201 213 204 
rect 210 204 213 207 
rect 210 207 213 210 
rect 210 210 213 213 
rect 210 213 213 216 
rect 210 216 213 219 
rect 210 219 213 222 
rect 210 222 213 225 
rect 210 225 213 228 
rect 210 228 213 231 
rect 210 231 213 234 
rect 210 234 213 237 
rect 210 237 213 240 
rect 210 240 213 243 
rect 210 243 213 246 
rect 210 246 213 249 
rect 210 249 213 252 
rect 210 252 213 255 
rect 210 255 213 258 
rect 210 258 213 261 
rect 210 261 213 264 
rect 210 264 213 267 
rect 210 267 213 270 
rect 210 270 213 273 
rect 210 273 213 276 
rect 210 276 213 279 
rect 210 279 213 282 
rect 210 282 213 285 
rect 210 285 213 288 
rect 210 288 213 291 
rect 210 291 213 294 
rect 210 294 213 297 
rect 210 297 213 300 
rect 210 300 213 303 
rect 210 303 213 306 
rect 210 306 213 309 
rect 210 309 213 312 
rect 210 312 213 315 
rect 210 315 213 318 
rect 210 318 213 321 
rect 210 321 213 324 
rect 210 324 213 327 
rect 210 327 213 330 
rect 210 330 213 333 
rect 210 333 213 336 
rect 210 336 213 339 
rect 210 339 213 342 
rect 210 342 213 345 
rect 210 345 213 348 
rect 210 348 213 351 
rect 210 351 213 354 
rect 210 354 213 357 
rect 210 357 213 360 
rect 210 360 213 363 
rect 210 363 213 366 
rect 210 366 213 369 
rect 210 369 213 372 
rect 210 372 213 375 
rect 210 375 213 378 
rect 210 378 213 381 
rect 210 381 213 384 
rect 210 384 213 387 
rect 210 387 213 390 
rect 210 390 213 393 
rect 210 393 213 396 
rect 210 396 213 399 
rect 210 399 213 402 
rect 210 402 213 405 
rect 210 405 213 408 
rect 210 408 213 411 
rect 210 411 213 414 
rect 210 414 213 417 
rect 210 417 213 420 
rect 210 420 213 423 
rect 210 423 213 426 
rect 210 426 213 429 
rect 210 429 213 432 
rect 210 432 213 435 
rect 210 435 213 438 
rect 210 438 213 441 
rect 210 441 213 444 
rect 210 444 213 447 
rect 210 447 213 450 
rect 210 450 213 453 
rect 210 453 213 456 
rect 210 456 213 459 
rect 210 459 213 462 
rect 210 462 213 465 
rect 210 465 213 468 
rect 210 468 213 471 
rect 210 471 213 474 
rect 210 474 213 477 
rect 210 477 213 480 
rect 210 480 213 483 
rect 210 483 213 486 
rect 210 486 213 489 
rect 210 489 213 492 
rect 210 492 213 495 
rect 210 495 213 498 
rect 210 498 213 501 
rect 210 501 213 504 
rect 210 504 213 507 
rect 210 507 213 510 
rect 213 0 216 3 
rect 213 3 216 6 
rect 213 6 216 9 
rect 213 9 216 12 
rect 213 12 216 15 
rect 213 15 216 18 
rect 213 18 216 21 
rect 213 21 216 24 
rect 213 24 216 27 
rect 213 27 216 30 
rect 213 30 216 33 
rect 213 33 216 36 
rect 213 36 216 39 
rect 213 39 216 42 
rect 213 42 216 45 
rect 213 45 216 48 
rect 213 48 216 51 
rect 213 51 216 54 
rect 213 54 216 57 
rect 213 57 216 60 
rect 213 60 216 63 
rect 213 63 216 66 
rect 213 66 216 69 
rect 213 69 216 72 
rect 213 72 216 75 
rect 213 75 216 78 
rect 213 78 216 81 
rect 213 81 216 84 
rect 213 84 216 87 
rect 213 87 216 90 
rect 213 90 216 93 
rect 213 93 216 96 
rect 213 96 216 99 
rect 213 99 216 102 
rect 213 102 216 105 
rect 213 105 216 108 
rect 213 108 216 111 
rect 213 111 216 114 
rect 213 114 216 117 
rect 213 117 216 120 
rect 213 120 216 123 
rect 213 123 216 126 
rect 213 126 216 129 
rect 213 129 216 132 
rect 213 132 216 135 
rect 213 135 216 138 
rect 213 138 216 141 
rect 213 141 216 144 
rect 213 144 216 147 
rect 213 147 216 150 
rect 213 150 216 153 
rect 213 153 216 156 
rect 213 156 216 159 
rect 213 159 216 162 
rect 213 162 216 165 
rect 213 165 216 168 
rect 213 168 216 171 
rect 213 171 216 174 
rect 213 174 216 177 
rect 213 177 216 180 
rect 213 180 216 183 
rect 213 183 216 186 
rect 213 186 216 189 
rect 213 189 216 192 
rect 213 192 216 195 
rect 213 195 216 198 
rect 213 198 216 201 
rect 213 201 216 204 
rect 213 204 216 207 
rect 213 207 216 210 
rect 213 210 216 213 
rect 213 213 216 216 
rect 213 216 216 219 
rect 213 219 216 222 
rect 213 222 216 225 
rect 213 225 216 228 
rect 213 228 216 231 
rect 213 231 216 234 
rect 213 234 216 237 
rect 213 237 216 240 
rect 213 240 216 243 
rect 213 243 216 246 
rect 213 246 216 249 
rect 213 249 216 252 
rect 213 252 216 255 
rect 213 255 216 258 
rect 213 258 216 261 
rect 213 261 216 264 
rect 213 264 216 267 
rect 213 267 216 270 
rect 213 270 216 273 
rect 213 273 216 276 
rect 213 276 216 279 
rect 213 279 216 282 
rect 213 282 216 285 
rect 213 285 216 288 
rect 213 288 216 291 
rect 213 291 216 294 
rect 213 294 216 297 
rect 213 297 216 300 
rect 213 300 216 303 
rect 213 303 216 306 
rect 213 306 216 309 
rect 213 309 216 312 
rect 213 312 216 315 
rect 213 315 216 318 
rect 213 318 216 321 
rect 213 321 216 324 
rect 213 324 216 327 
rect 213 327 216 330 
rect 213 330 216 333 
rect 213 333 216 336 
rect 213 336 216 339 
rect 213 339 216 342 
rect 213 342 216 345 
rect 213 345 216 348 
rect 213 348 216 351 
rect 213 351 216 354 
rect 213 354 216 357 
rect 213 357 216 360 
rect 213 360 216 363 
rect 213 363 216 366 
rect 213 366 216 369 
rect 213 369 216 372 
rect 213 372 216 375 
rect 213 375 216 378 
rect 213 378 216 381 
rect 213 381 216 384 
rect 213 384 216 387 
rect 213 387 216 390 
rect 213 390 216 393 
rect 213 393 216 396 
rect 213 396 216 399 
rect 213 399 216 402 
rect 213 402 216 405 
rect 213 405 216 408 
rect 213 408 216 411 
rect 213 411 216 414 
rect 213 414 216 417 
rect 213 417 216 420 
rect 213 420 216 423 
rect 213 423 216 426 
rect 213 426 216 429 
rect 213 429 216 432 
rect 213 432 216 435 
rect 213 435 216 438 
rect 213 438 216 441 
rect 213 441 216 444 
rect 213 444 216 447 
rect 213 447 216 450 
rect 213 450 216 453 
rect 213 453 216 456 
rect 213 456 216 459 
rect 213 459 216 462 
rect 213 462 216 465 
rect 213 465 216 468 
rect 213 468 216 471 
rect 213 471 216 474 
rect 213 474 216 477 
rect 213 477 216 480 
rect 213 480 216 483 
rect 213 483 216 486 
rect 213 486 216 489 
rect 213 489 216 492 
rect 213 492 216 495 
rect 213 495 216 498 
rect 213 498 216 501 
rect 213 501 216 504 
rect 213 504 216 507 
rect 213 507 216 510 
rect 216 0 219 3 
rect 216 3 219 6 
rect 216 6 219 9 
rect 216 9 219 12 
rect 216 12 219 15 
rect 216 15 219 18 
rect 216 18 219 21 
rect 216 21 219 24 
rect 216 24 219 27 
rect 216 27 219 30 
rect 216 30 219 33 
rect 216 33 219 36 
rect 216 36 219 39 
rect 216 39 219 42 
rect 216 42 219 45 
rect 216 45 219 48 
rect 216 48 219 51 
rect 216 51 219 54 
rect 216 54 219 57 
rect 216 57 219 60 
rect 216 60 219 63 
rect 216 63 219 66 
rect 216 66 219 69 
rect 216 69 219 72 
rect 216 72 219 75 
rect 216 75 219 78 
rect 216 78 219 81 
rect 216 81 219 84 
rect 216 84 219 87 
rect 216 87 219 90 
rect 216 90 219 93 
rect 216 93 219 96 
rect 216 96 219 99 
rect 216 99 219 102 
rect 216 102 219 105 
rect 216 105 219 108 
rect 216 108 219 111 
rect 216 111 219 114 
rect 216 114 219 117 
rect 216 117 219 120 
rect 216 120 219 123 
rect 216 123 219 126 
rect 216 126 219 129 
rect 216 129 219 132 
rect 216 132 219 135 
rect 216 135 219 138 
rect 216 138 219 141 
rect 216 141 219 144 
rect 216 144 219 147 
rect 216 147 219 150 
rect 216 150 219 153 
rect 216 153 219 156 
rect 216 156 219 159 
rect 216 159 219 162 
rect 216 162 219 165 
rect 216 165 219 168 
rect 216 168 219 171 
rect 216 171 219 174 
rect 216 174 219 177 
rect 216 177 219 180 
rect 216 180 219 183 
rect 216 183 219 186 
rect 216 186 219 189 
rect 216 189 219 192 
rect 216 192 219 195 
rect 216 195 219 198 
rect 216 198 219 201 
rect 216 201 219 204 
rect 216 204 219 207 
rect 216 207 219 210 
rect 216 210 219 213 
rect 216 213 219 216 
rect 216 216 219 219 
rect 216 219 219 222 
rect 216 222 219 225 
rect 216 225 219 228 
rect 216 228 219 231 
rect 216 231 219 234 
rect 216 234 219 237 
rect 216 237 219 240 
rect 216 240 219 243 
rect 216 243 219 246 
rect 216 246 219 249 
rect 216 249 219 252 
rect 216 252 219 255 
rect 216 255 219 258 
rect 216 258 219 261 
rect 216 261 219 264 
rect 216 264 219 267 
rect 216 267 219 270 
rect 216 270 219 273 
rect 216 273 219 276 
rect 216 276 219 279 
rect 216 279 219 282 
rect 216 282 219 285 
rect 216 285 219 288 
rect 216 288 219 291 
rect 216 291 219 294 
rect 216 294 219 297 
rect 216 297 219 300 
rect 216 300 219 303 
rect 216 303 219 306 
rect 216 306 219 309 
rect 216 309 219 312 
rect 216 312 219 315 
rect 216 315 219 318 
rect 216 318 219 321 
rect 216 321 219 324 
rect 216 324 219 327 
rect 216 327 219 330 
rect 216 330 219 333 
rect 216 333 219 336 
rect 216 336 219 339 
rect 216 339 219 342 
rect 216 342 219 345 
rect 216 345 219 348 
rect 216 348 219 351 
rect 216 351 219 354 
rect 216 354 219 357 
rect 216 357 219 360 
rect 216 360 219 363 
rect 216 363 219 366 
rect 216 366 219 369 
rect 216 369 219 372 
rect 216 372 219 375 
rect 216 375 219 378 
rect 216 378 219 381 
rect 216 381 219 384 
rect 216 384 219 387 
rect 216 387 219 390 
rect 216 390 219 393 
rect 216 393 219 396 
rect 216 396 219 399 
rect 216 399 219 402 
rect 216 402 219 405 
rect 216 405 219 408 
rect 216 408 219 411 
rect 216 411 219 414 
rect 216 414 219 417 
rect 216 417 219 420 
rect 216 420 219 423 
rect 216 423 219 426 
rect 216 426 219 429 
rect 216 429 219 432 
rect 216 432 219 435 
rect 216 435 219 438 
rect 216 438 219 441 
rect 216 441 219 444 
rect 216 444 219 447 
rect 216 447 219 450 
rect 216 450 219 453 
rect 216 453 219 456 
rect 216 456 219 459 
rect 216 459 219 462 
rect 216 462 219 465 
rect 216 465 219 468 
rect 216 468 219 471 
rect 216 471 219 474 
rect 216 474 219 477 
rect 216 477 219 480 
rect 216 480 219 483 
rect 216 483 219 486 
rect 216 486 219 489 
rect 216 489 219 492 
rect 216 492 219 495 
rect 216 495 219 498 
rect 216 498 219 501 
rect 216 501 219 504 
rect 216 504 219 507 
rect 216 507 219 510 
rect 219 0 222 3 
rect 219 3 222 6 
rect 219 6 222 9 
rect 219 9 222 12 
rect 219 12 222 15 
rect 219 15 222 18 
rect 219 18 222 21 
rect 219 21 222 24 
rect 219 24 222 27 
rect 219 27 222 30 
rect 219 30 222 33 
rect 219 33 222 36 
rect 219 36 222 39 
rect 219 39 222 42 
rect 219 42 222 45 
rect 219 45 222 48 
rect 219 48 222 51 
rect 219 51 222 54 
rect 219 54 222 57 
rect 219 57 222 60 
rect 219 60 222 63 
rect 219 63 222 66 
rect 219 66 222 69 
rect 219 69 222 72 
rect 219 72 222 75 
rect 219 75 222 78 
rect 219 78 222 81 
rect 219 81 222 84 
rect 219 84 222 87 
rect 219 87 222 90 
rect 219 90 222 93 
rect 219 93 222 96 
rect 219 96 222 99 
rect 219 99 222 102 
rect 219 102 222 105 
rect 219 105 222 108 
rect 219 108 222 111 
rect 219 111 222 114 
rect 219 114 222 117 
rect 219 117 222 120 
rect 219 120 222 123 
rect 219 123 222 126 
rect 219 126 222 129 
rect 219 129 222 132 
rect 219 132 222 135 
rect 219 135 222 138 
rect 219 138 222 141 
rect 219 141 222 144 
rect 219 144 222 147 
rect 219 147 222 150 
rect 219 150 222 153 
rect 219 153 222 156 
rect 219 156 222 159 
rect 219 159 222 162 
rect 219 162 222 165 
rect 219 165 222 168 
rect 219 168 222 171 
rect 219 171 222 174 
rect 219 174 222 177 
rect 219 177 222 180 
rect 219 180 222 183 
rect 219 183 222 186 
rect 219 186 222 189 
rect 219 189 222 192 
rect 219 192 222 195 
rect 219 195 222 198 
rect 219 198 222 201 
rect 219 201 222 204 
rect 219 204 222 207 
rect 219 207 222 210 
rect 219 210 222 213 
rect 219 213 222 216 
rect 219 216 222 219 
rect 219 219 222 222 
rect 219 222 222 225 
rect 219 225 222 228 
rect 219 228 222 231 
rect 219 231 222 234 
rect 219 234 222 237 
rect 219 237 222 240 
rect 219 240 222 243 
rect 219 243 222 246 
rect 219 246 222 249 
rect 219 249 222 252 
rect 219 252 222 255 
rect 219 255 222 258 
rect 219 258 222 261 
rect 219 261 222 264 
rect 219 264 222 267 
rect 219 267 222 270 
rect 219 270 222 273 
rect 219 273 222 276 
rect 219 276 222 279 
rect 219 279 222 282 
rect 219 282 222 285 
rect 219 285 222 288 
rect 219 288 222 291 
rect 219 291 222 294 
rect 219 294 222 297 
rect 219 297 222 300 
rect 219 300 222 303 
rect 219 303 222 306 
rect 219 306 222 309 
rect 219 309 222 312 
rect 219 312 222 315 
rect 219 315 222 318 
rect 219 318 222 321 
rect 219 321 222 324 
rect 219 324 222 327 
rect 219 327 222 330 
rect 219 330 222 333 
rect 219 333 222 336 
rect 219 336 222 339 
rect 219 339 222 342 
rect 219 342 222 345 
rect 219 345 222 348 
rect 219 348 222 351 
rect 219 351 222 354 
rect 219 354 222 357 
rect 219 357 222 360 
rect 219 360 222 363 
rect 219 363 222 366 
rect 219 366 222 369 
rect 219 369 222 372 
rect 219 372 222 375 
rect 219 375 222 378 
rect 219 378 222 381 
rect 219 381 222 384 
rect 219 384 222 387 
rect 219 387 222 390 
rect 219 390 222 393 
rect 219 393 222 396 
rect 219 396 222 399 
rect 219 399 222 402 
rect 219 402 222 405 
rect 219 405 222 408 
rect 219 408 222 411 
rect 219 411 222 414 
rect 219 414 222 417 
rect 219 417 222 420 
rect 219 420 222 423 
rect 219 423 222 426 
rect 219 426 222 429 
rect 219 429 222 432 
rect 219 432 222 435 
rect 219 435 222 438 
rect 219 438 222 441 
rect 219 441 222 444 
rect 219 444 222 447 
rect 219 447 222 450 
rect 219 450 222 453 
rect 219 453 222 456 
rect 219 456 222 459 
rect 219 459 222 462 
rect 219 462 222 465 
rect 219 465 222 468 
rect 219 468 222 471 
rect 219 471 222 474 
rect 219 474 222 477 
rect 219 477 222 480 
rect 219 480 222 483 
rect 219 483 222 486 
rect 219 486 222 489 
rect 219 489 222 492 
rect 219 492 222 495 
rect 219 495 222 498 
rect 219 498 222 501 
rect 219 501 222 504 
rect 219 504 222 507 
rect 219 507 222 510 
rect 222 0 225 3 
rect 222 3 225 6 
rect 222 6 225 9 
rect 222 9 225 12 
rect 222 12 225 15 
rect 222 15 225 18 
rect 222 18 225 21 
rect 222 21 225 24 
rect 222 24 225 27 
rect 222 27 225 30 
rect 222 30 225 33 
rect 222 33 225 36 
rect 222 36 225 39 
rect 222 39 225 42 
rect 222 42 225 45 
rect 222 45 225 48 
rect 222 48 225 51 
rect 222 51 225 54 
rect 222 54 225 57 
rect 222 57 225 60 
rect 222 60 225 63 
rect 222 63 225 66 
rect 222 66 225 69 
rect 222 69 225 72 
rect 222 72 225 75 
rect 222 75 225 78 
rect 222 78 225 81 
rect 222 81 225 84 
rect 222 84 225 87 
rect 222 87 225 90 
rect 222 90 225 93 
rect 222 93 225 96 
rect 222 96 225 99 
rect 222 99 225 102 
rect 222 102 225 105 
rect 222 105 225 108 
rect 222 108 225 111 
rect 222 111 225 114 
rect 222 114 225 117 
rect 222 117 225 120 
rect 222 120 225 123 
rect 222 123 225 126 
rect 222 126 225 129 
rect 222 129 225 132 
rect 222 132 225 135 
rect 222 135 225 138 
rect 222 138 225 141 
rect 222 141 225 144 
rect 222 144 225 147 
rect 222 147 225 150 
rect 222 150 225 153 
rect 222 153 225 156 
rect 222 156 225 159 
rect 222 159 225 162 
rect 222 162 225 165 
rect 222 165 225 168 
rect 222 168 225 171 
rect 222 171 225 174 
rect 222 174 225 177 
rect 222 177 225 180 
rect 222 180 225 183 
rect 222 183 225 186 
rect 222 186 225 189 
rect 222 189 225 192 
rect 222 192 225 195 
rect 222 195 225 198 
rect 222 198 225 201 
rect 222 201 225 204 
rect 222 204 225 207 
rect 222 207 225 210 
rect 222 210 225 213 
rect 222 213 225 216 
rect 222 216 225 219 
rect 222 219 225 222 
rect 222 222 225 225 
rect 222 225 225 228 
rect 222 228 225 231 
rect 222 231 225 234 
rect 222 234 225 237 
rect 222 237 225 240 
rect 222 240 225 243 
rect 222 243 225 246 
rect 222 246 225 249 
rect 222 249 225 252 
rect 222 252 225 255 
rect 222 255 225 258 
rect 222 258 225 261 
rect 222 261 225 264 
rect 222 264 225 267 
rect 222 267 225 270 
rect 222 270 225 273 
rect 222 273 225 276 
rect 222 276 225 279 
rect 222 279 225 282 
rect 222 282 225 285 
rect 222 285 225 288 
rect 222 288 225 291 
rect 222 291 225 294 
rect 222 294 225 297 
rect 222 297 225 300 
rect 222 300 225 303 
rect 222 303 225 306 
rect 222 306 225 309 
rect 222 309 225 312 
rect 222 312 225 315 
rect 222 315 225 318 
rect 222 318 225 321 
rect 222 321 225 324 
rect 222 324 225 327 
rect 222 327 225 330 
rect 222 330 225 333 
rect 222 333 225 336 
rect 222 336 225 339 
rect 222 339 225 342 
rect 222 342 225 345 
rect 222 345 225 348 
rect 222 348 225 351 
rect 222 351 225 354 
rect 222 354 225 357 
rect 222 357 225 360 
rect 222 360 225 363 
rect 222 363 225 366 
rect 222 366 225 369 
rect 222 369 225 372 
rect 222 372 225 375 
rect 222 375 225 378 
rect 222 378 225 381 
rect 222 381 225 384 
rect 222 384 225 387 
rect 222 387 225 390 
rect 222 390 225 393 
rect 222 393 225 396 
rect 222 396 225 399 
rect 222 399 225 402 
rect 222 402 225 405 
rect 222 405 225 408 
rect 222 408 225 411 
rect 222 411 225 414 
rect 222 414 225 417 
rect 222 417 225 420 
rect 222 420 225 423 
rect 222 423 225 426 
rect 222 426 225 429 
rect 222 429 225 432 
rect 222 432 225 435 
rect 222 435 225 438 
rect 222 438 225 441 
rect 222 441 225 444 
rect 222 444 225 447 
rect 222 447 225 450 
rect 222 450 225 453 
rect 222 453 225 456 
rect 222 456 225 459 
rect 222 459 225 462 
rect 222 462 225 465 
rect 222 465 225 468 
rect 222 468 225 471 
rect 222 471 225 474 
rect 222 474 225 477 
rect 222 477 225 480 
rect 222 480 225 483 
rect 222 483 225 486 
rect 222 486 225 489 
rect 222 489 225 492 
rect 222 492 225 495 
rect 222 495 225 498 
rect 222 498 225 501 
rect 222 501 225 504 
rect 222 504 225 507 
rect 222 507 225 510 
rect 225 0 228 3 
rect 225 3 228 6 
rect 225 6 228 9 
rect 225 9 228 12 
rect 225 12 228 15 
rect 225 15 228 18 
rect 225 18 228 21 
rect 225 21 228 24 
rect 225 24 228 27 
rect 225 27 228 30 
rect 225 30 228 33 
rect 225 33 228 36 
rect 225 36 228 39 
rect 225 39 228 42 
rect 225 42 228 45 
rect 225 45 228 48 
rect 225 48 228 51 
rect 225 51 228 54 
rect 225 54 228 57 
rect 225 57 228 60 
rect 225 60 228 63 
rect 225 63 228 66 
rect 225 66 228 69 
rect 225 69 228 72 
rect 225 72 228 75 
rect 225 75 228 78 
rect 225 78 228 81 
rect 225 81 228 84 
rect 225 84 228 87 
rect 225 87 228 90 
rect 225 90 228 93 
rect 225 93 228 96 
rect 225 96 228 99 
rect 225 99 228 102 
rect 225 102 228 105 
rect 225 105 228 108 
rect 225 108 228 111 
rect 225 111 228 114 
rect 225 114 228 117 
rect 225 117 228 120 
rect 225 120 228 123 
rect 225 123 228 126 
rect 225 126 228 129 
rect 225 129 228 132 
rect 225 132 228 135 
rect 225 135 228 138 
rect 225 138 228 141 
rect 225 141 228 144 
rect 225 144 228 147 
rect 225 147 228 150 
rect 225 150 228 153 
rect 225 153 228 156 
rect 225 156 228 159 
rect 225 159 228 162 
rect 225 162 228 165 
rect 225 165 228 168 
rect 225 168 228 171 
rect 225 171 228 174 
rect 225 174 228 177 
rect 225 177 228 180 
rect 225 180 228 183 
rect 225 183 228 186 
rect 225 186 228 189 
rect 225 189 228 192 
rect 225 192 228 195 
rect 225 195 228 198 
rect 225 198 228 201 
rect 225 201 228 204 
rect 225 204 228 207 
rect 225 207 228 210 
rect 225 210 228 213 
rect 225 213 228 216 
rect 225 216 228 219 
rect 225 219 228 222 
rect 225 222 228 225 
rect 225 225 228 228 
rect 225 228 228 231 
rect 225 231 228 234 
rect 225 234 228 237 
rect 225 237 228 240 
rect 225 240 228 243 
rect 225 243 228 246 
rect 225 246 228 249 
rect 225 249 228 252 
rect 225 252 228 255 
rect 225 255 228 258 
rect 225 258 228 261 
rect 225 261 228 264 
rect 225 264 228 267 
rect 225 267 228 270 
rect 225 270 228 273 
rect 225 273 228 276 
rect 225 276 228 279 
rect 225 279 228 282 
rect 225 282 228 285 
rect 225 285 228 288 
rect 225 288 228 291 
rect 225 291 228 294 
rect 225 294 228 297 
rect 225 297 228 300 
rect 225 300 228 303 
rect 225 303 228 306 
rect 225 306 228 309 
rect 225 309 228 312 
rect 225 312 228 315 
rect 225 315 228 318 
rect 225 318 228 321 
rect 225 321 228 324 
rect 225 324 228 327 
rect 225 327 228 330 
rect 225 330 228 333 
rect 225 333 228 336 
rect 225 336 228 339 
rect 225 339 228 342 
rect 225 342 228 345 
rect 225 345 228 348 
rect 225 348 228 351 
rect 225 351 228 354 
rect 225 354 228 357 
rect 225 357 228 360 
rect 225 360 228 363 
rect 225 363 228 366 
rect 225 366 228 369 
rect 225 369 228 372 
rect 225 372 228 375 
rect 225 375 228 378 
rect 225 378 228 381 
rect 225 381 228 384 
rect 225 384 228 387 
rect 225 387 228 390 
rect 225 390 228 393 
rect 225 393 228 396 
rect 225 396 228 399 
rect 225 399 228 402 
rect 225 402 228 405 
rect 225 405 228 408 
rect 225 408 228 411 
rect 225 411 228 414 
rect 225 414 228 417 
rect 225 417 228 420 
rect 225 420 228 423 
rect 225 423 228 426 
rect 225 426 228 429 
rect 225 429 228 432 
rect 225 432 228 435 
rect 225 435 228 438 
rect 225 438 228 441 
rect 225 441 228 444 
rect 225 444 228 447 
rect 225 447 228 450 
rect 225 450 228 453 
rect 225 453 228 456 
rect 225 456 228 459 
rect 225 459 228 462 
rect 225 462 228 465 
rect 225 465 228 468 
rect 225 468 228 471 
rect 225 471 228 474 
rect 225 474 228 477 
rect 225 477 228 480 
rect 225 480 228 483 
rect 225 483 228 486 
rect 225 486 228 489 
rect 225 489 228 492 
rect 225 492 228 495 
rect 225 495 228 498 
rect 225 498 228 501 
rect 225 501 228 504 
rect 225 504 228 507 
rect 225 507 228 510 
rect 228 0 231 3 
rect 228 3 231 6 
rect 228 6 231 9 
rect 228 9 231 12 
rect 228 12 231 15 
rect 228 15 231 18 
rect 228 18 231 21 
rect 228 21 231 24 
rect 228 24 231 27 
rect 228 27 231 30 
rect 228 30 231 33 
rect 228 33 231 36 
rect 228 36 231 39 
rect 228 39 231 42 
rect 228 42 231 45 
rect 228 45 231 48 
rect 228 48 231 51 
rect 228 51 231 54 
rect 228 54 231 57 
rect 228 57 231 60 
rect 228 60 231 63 
rect 228 63 231 66 
rect 228 66 231 69 
rect 228 69 231 72 
rect 228 72 231 75 
rect 228 75 231 78 
rect 228 78 231 81 
rect 228 81 231 84 
rect 228 84 231 87 
rect 228 87 231 90 
rect 228 90 231 93 
rect 228 93 231 96 
rect 228 96 231 99 
rect 228 99 231 102 
rect 228 102 231 105 
rect 228 105 231 108 
rect 228 108 231 111 
rect 228 111 231 114 
rect 228 114 231 117 
rect 228 117 231 120 
rect 228 120 231 123 
rect 228 123 231 126 
rect 228 126 231 129 
rect 228 129 231 132 
rect 228 132 231 135 
rect 228 135 231 138 
rect 228 138 231 141 
rect 228 141 231 144 
rect 228 144 231 147 
rect 228 147 231 150 
rect 228 150 231 153 
rect 228 153 231 156 
rect 228 156 231 159 
rect 228 159 231 162 
rect 228 162 231 165 
rect 228 165 231 168 
rect 228 168 231 171 
rect 228 171 231 174 
rect 228 174 231 177 
rect 228 177 231 180 
rect 228 180 231 183 
rect 228 183 231 186 
rect 228 186 231 189 
rect 228 189 231 192 
rect 228 192 231 195 
rect 228 195 231 198 
rect 228 198 231 201 
rect 228 201 231 204 
rect 228 204 231 207 
rect 228 207 231 210 
rect 228 210 231 213 
rect 228 213 231 216 
rect 228 216 231 219 
rect 228 219 231 222 
rect 228 222 231 225 
rect 228 225 231 228 
rect 228 228 231 231 
rect 228 231 231 234 
rect 228 234 231 237 
rect 228 237 231 240 
rect 228 240 231 243 
rect 228 243 231 246 
rect 228 246 231 249 
rect 228 249 231 252 
rect 228 252 231 255 
rect 228 255 231 258 
rect 228 258 231 261 
rect 228 261 231 264 
rect 228 264 231 267 
rect 228 267 231 270 
rect 228 270 231 273 
rect 228 273 231 276 
rect 228 276 231 279 
rect 228 279 231 282 
rect 228 282 231 285 
rect 228 285 231 288 
rect 228 288 231 291 
rect 228 291 231 294 
rect 228 294 231 297 
rect 228 297 231 300 
rect 228 300 231 303 
rect 228 303 231 306 
rect 228 306 231 309 
rect 228 309 231 312 
rect 228 312 231 315 
rect 228 315 231 318 
rect 228 318 231 321 
rect 228 321 231 324 
rect 228 324 231 327 
rect 228 327 231 330 
rect 228 330 231 333 
rect 228 333 231 336 
rect 228 336 231 339 
rect 228 339 231 342 
rect 228 342 231 345 
rect 228 345 231 348 
rect 228 348 231 351 
rect 228 351 231 354 
rect 228 354 231 357 
rect 228 357 231 360 
rect 228 360 231 363 
rect 228 363 231 366 
rect 228 366 231 369 
rect 228 369 231 372 
rect 228 372 231 375 
rect 228 375 231 378 
rect 228 378 231 381 
rect 228 381 231 384 
rect 228 384 231 387 
rect 228 387 231 390 
rect 228 390 231 393 
rect 228 393 231 396 
rect 228 396 231 399 
rect 228 399 231 402 
rect 228 402 231 405 
rect 228 405 231 408 
rect 228 408 231 411 
rect 228 411 231 414 
rect 228 414 231 417 
rect 228 417 231 420 
rect 228 420 231 423 
rect 228 423 231 426 
rect 228 426 231 429 
rect 228 429 231 432 
rect 228 432 231 435 
rect 228 435 231 438 
rect 228 438 231 441 
rect 228 441 231 444 
rect 228 444 231 447 
rect 228 447 231 450 
rect 228 450 231 453 
rect 228 453 231 456 
rect 228 456 231 459 
rect 228 459 231 462 
rect 228 462 231 465 
rect 228 465 231 468 
rect 228 468 231 471 
rect 228 471 231 474 
rect 228 474 231 477 
rect 228 477 231 480 
rect 228 480 231 483 
rect 228 483 231 486 
rect 228 486 231 489 
rect 228 489 231 492 
rect 228 492 231 495 
rect 228 495 231 498 
rect 228 498 231 501 
rect 228 501 231 504 
rect 228 504 231 507 
rect 228 507 231 510 
rect 231 0 234 3 
rect 231 3 234 6 
rect 231 6 234 9 
rect 231 9 234 12 
rect 231 12 234 15 
rect 231 15 234 18 
rect 231 18 234 21 
rect 231 21 234 24 
rect 231 24 234 27 
rect 231 27 234 30 
rect 231 30 234 33 
rect 231 33 234 36 
rect 231 36 234 39 
rect 231 39 234 42 
rect 231 42 234 45 
rect 231 45 234 48 
rect 231 48 234 51 
rect 231 51 234 54 
rect 231 54 234 57 
rect 231 57 234 60 
rect 231 60 234 63 
rect 231 63 234 66 
rect 231 66 234 69 
rect 231 69 234 72 
rect 231 72 234 75 
rect 231 75 234 78 
rect 231 78 234 81 
rect 231 81 234 84 
rect 231 84 234 87 
rect 231 87 234 90 
rect 231 90 234 93 
rect 231 93 234 96 
rect 231 96 234 99 
rect 231 99 234 102 
rect 231 102 234 105 
rect 231 105 234 108 
rect 231 108 234 111 
rect 231 111 234 114 
rect 231 114 234 117 
rect 231 117 234 120 
rect 231 120 234 123 
rect 231 123 234 126 
rect 231 126 234 129 
rect 231 129 234 132 
rect 231 132 234 135 
rect 231 135 234 138 
rect 231 138 234 141 
rect 231 141 234 144 
rect 231 144 234 147 
rect 231 147 234 150 
rect 231 150 234 153 
rect 231 153 234 156 
rect 231 156 234 159 
rect 231 159 234 162 
rect 231 162 234 165 
rect 231 165 234 168 
rect 231 168 234 171 
rect 231 171 234 174 
rect 231 174 234 177 
rect 231 177 234 180 
rect 231 180 234 183 
rect 231 183 234 186 
rect 231 186 234 189 
rect 231 189 234 192 
rect 231 192 234 195 
rect 231 195 234 198 
rect 231 198 234 201 
rect 231 201 234 204 
rect 231 204 234 207 
rect 231 207 234 210 
rect 231 210 234 213 
rect 231 213 234 216 
rect 231 216 234 219 
rect 231 219 234 222 
rect 231 222 234 225 
rect 231 225 234 228 
rect 231 228 234 231 
rect 231 231 234 234 
rect 231 234 234 237 
rect 231 237 234 240 
rect 231 240 234 243 
rect 231 243 234 246 
rect 231 246 234 249 
rect 231 249 234 252 
rect 231 252 234 255 
rect 231 255 234 258 
rect 231 258 234 261 
rect 231 261 234 264 
rect 231 264 234 267 
rect 231 267 234 270 
rect 231 270 234 273 
rect 231 273 234 276 
rect 231 276 234 279 
rect 231 279 234 282 
rect 231 282 234 285 
rect 231 285 234 288 
rect 231 288 234 291 
rect 231 291 234 294 
rect 231 294 234 297 
rect 231 297 234 300 
rect 231 300 234 303 
rect 231 303 234 306 
rect 231 306 234 309 
rect 231 309 234 312 
rect 231 312 234 315 
rect 231 315 234 318 
rect 231 318 234 321 
rect 231 321 234 324 
rect 231 324 234 327 
rect 231 327 234 330 
rect 231 330 234 333 
rect 231 333 234 336 
rect 231 336 234 339 
rect 231 339 234 342 
rect 231 342 234 345 
rect 231 345 234 348 
rect 231 348 234 351 
rect 231 351 234 354 
rect 231 354 234 357 
rect 231 357 234 360 
rect 231 360 234 363 
rect 231 363 234 366 
rect 231 366 234 369 
rect 231 369 234 372 
rect 231 372 234 375 
rect 231 375 234 378 
rect 231 378 234 381 
rect 231 381 234 384 
rect 231 384 234 387 
rect 231 387 234 390 
rect 231 390 234 393 
rect 231 393 234 396 
rect 231 396 234 399 
rect 231 399 234 402 
rect 231 402 234 405 
rect 231 405 234 408 
rect 231 408 234 411 
rect 231 411 234 414 
rect 231 414 234 417 
rect 231 417 234 420 
rect 231 420 234 423 
rect 231 423 234 426 
rect 231 426 234 429 
rect 231 429 234 432 
rect 231 432 234 435 
rect 231 435 234 438 
rect 231 438 234 441 
rect 231 441 234 444 
rect 231 444 234 447 
rect 231 447 234 450 
rect 231 450 234 453 
rect 231 453 234 456 
rect 231 456 234 459 
rect 231 459 234 462 
rect 231 462 234 465 
rect 231 465 234 468 
rect 231 468 234 471 
rect 231 471 234 474 
rect 231 474 234 477 
rect 231 477 234 480 
rect 231 480 234 483 
rect 231 483 234 486 
rect 231 486 234 489 
rect 231 489 234 492 
rect 231 492 234 495 
rect 231 495 234 498 
rect 231 498 234 501 
rect 231 501 234 504 
rect 231 504 234 507 
rect 231 507 234 510 
rect 234 0 237 3 
rect 234 3 237 6 
rect 234 6 237 9 
rect 234 9 237 12 
rect 234 12 237 15 
rect 234 15 237 18 
rect 234 18 237 21 
rect 234 21 237 24 
rect 234 24 237 27 
rect 234 27 237 30 
rect 234 30 237 33 
rect 234 33 237 36 
rect 234 36 237 39 
rect 234 39 237 42 
rect 234 42 237 45 
rect 234 45 237 48 
rect 234 48 237 51 
rect 234 51 237 54 
rect 234 54 237 57 
rect 234 57 237 60 
rect 234 60 237 63 
rect 234 63 237 66 
rect 234 66 237 69 
rect 234 69 237 72 
rect 234 72 237 75 
rect 234 75 237 78 
rect 234 78 237 81 
rect 234 81 237 84 
rect 234 84 237 87 
rect 234 87 237 90 
rect 234 90 237 93 
rect 234 93 237 96 
rect 234 96 237 99 
rect 234 99 237 102 
rect 234 102 237 105 
rect 234 105 237 108 
rect 234 108 237 111 
rect 234 111 237 114 
rect 234 114 237 117 
rect 234 117 237 120 
rect 234 120 237 123 
rect 234 123 237 126 
rect 234 126 237 129 
rect 234 129 237 132 
rect 234 132 237 135 
rect 234 135 237 138 
rect 234 138 237 141 
rect 234 141 237 144 
rect 234 144 237 147 
rect 234 147 237 150 
rect 234 150 237 153 
rect 234 153 237 156 
rect 234 156 237 159 
rect 234 159 237 162 
rect 234 162 237 165 
rect 234 165 237 168 
rect 234 168 237 171 
rect 234 171 237 174 
rect 234 174 237 177 
rect 234 177 237 180 
rect 234 180 237 183 
rect 234 183 237 186 
rect 234 186 237 189 
rect 234 189 237 192 
rect 234 192 237 195 
rect 234 195 237 198 
rect 234 198 237 201 
rect 234 201 237 204 
rect 234 204 237 207 
rect 234 207 237 210 
rect 234 210 237 213 
rect 234 213 237 216 
rect 234 216 237 219 
rect 234 219 237 222 
rect 234 222 237 225 
rect 234 225 237 228 
rect 234 228 237 231 
rect 234 231 237 234 
rect 234 234 237 237 
rect 234 237 237 240 
rect 234 240 237 243 
rect 234 243 237 246 
rect 234 246 237 249 
rect 234 249 237 252 
rect 234 252 237 255 
rect 234 255 237 258 
rect 234 258 237 261 
rect 234 261 237 264 
rect 234 264 237 267 
rect 234 267 237 270 
rect 234 270 237 273 
rect 234 273 237 276 
rect 234 276 237 279 
rect 234 279 237 282 
rect 234 282 237 285 
rect 234 285 237 288 
rect 234 288 237 291 
rect 234 291 237 294 
rect 234 294 237 297 
rect 234 297 237 300 
rect 234 300 237 303 
rect 234 303 237 306 
rect 234 306 237 309 
rect 234 309 237 312 
rect 234 312 237 315 
rect 234 315 237 318 
rect 234 318 237 321 
rect 234 321 237 324 
rect 234 324 237 327 
rect 234 327 237 330 
rect 234 330 237 333 
rect 234 333 237 336 
rect 234 336 237 339 
rect 234 339 237 342 
rect 234 342 237 345 
rect 234 345 237 348 
rect 234 348 237 351 
rect 234 351 237 354 
rect 234 354 237 357 
rect 234 357 237 360 
rect 234 360 237 363 
rect 234 363 237 366 
rect 234 366 237 369 
rect 234 369 237 372 
rect 234 372 237 375 
rect 234 375 237 378 
rect 234 378 237 381 
rect 234 381 237 384 
rect 234 384 237 387 
rect 234 387 237 390 
rect 234 390 237 393 
rect 234 393 237 396 
rect 234 396 237 399 
rect 234 399 237 402 
rect 234 402 237 405 
rect 234 405 237 408 
rect 234 408 237 411 
rect 234 411 237 414 
rect 234 414 237 417 
rect 234 417 237 420 
rect 234 420 237 423 
rect 234 423 237 426 
rect 234 426 237 429 
rect 234 429 237 432 
rect 234 432 237 435 
rect 234 435 237 438 
rect 234 438 237 441 
rect 234 441 237 444 
rect 234 444 237 447 
rect 234 447 237 450 
rect 234 450 237 453 
rect 234 453 237 456 
rect 234 456 237 459 
rect 234 459 237 462 
rect 234 462 237 465 
rect 234 465 237 468 
rect 234 468 237 471 
rect 234 471 237 474 
rect 234 474 237 477 
rect 234 477 237 480 
rect 234 480 237 483 
rect 234 483 237 486 
rect 234 486 237 489 
rect 234 489 237 492 
rect 234 492 237 495 
rect 234 495 237 498 
rect 234 498 237 501 
rect 234 501 237 504 
rect 234 504 237 507 
rect 234 507 237 510 
rect 237 0 240 3 
rect 237 3 240 6 
rect 237 6 240 9 
rect 237 9 240 12 
rect 237 12 240 15 
rect 237 15 240 18 
rect 237 18 240 21 
rect 237 21 240 24 
rect 237 24 240 27 
rect 237 27 240 30 
rect 237 30 240 33 
rect 237 33 240 36 
rect 237 36 240 39 
rect 237 39 240 42 
rect 237 42 240 45 
rect 237 45 240 48 
rect 237 48 240 51 
rect 237 51 240 54 
rect 237 54 240 57 
rect 237 57 240 60 
rect 237 60 240 63 
rect 237 63 240 66 
rect 237 66 240 69 
rect 237 69 240 72 
rect 237 72 240 75 
rect 237 75 240 78 
rect 237 78 240 81 
rect 237 81 240 84 
rect 237 84 240 87 
rect 237 87 240 90 
rect 237 90 240 93 
rect 237 93 240 96 
rect 237 96 240 99 
rect 237 99 240 102 
rect 237 102 240 105 
rect 237 105 240 108 
rect 237 108 240 111 
rect 237 111 240 114 
rect 237 114 240 117 
rect 237 117 240 120 
rect 237 120 240 123 
rect 237 123 240 126 
rect 237 126 240 129 
rect 237 129 240 132 
rect 237 132 240 135 
rect 237 135 240 138 
rect 237 138 240 141 
rect 237 141 240 144 
rect 237 144 240 147 
rect 237 147 240 150 
rect 237 150 240 153 
rect 237 153 240 156 
rect 237 156 240 159 
rect 237 159 240 162 
rect 237 162 240 165 
rect 237 165 240 168 
rect 237 168 240 171 
rect 237 171 240 174 
rect 237 174 240 177 
rect 237 177 240 180 
rect 237 180 240 183 
rect 237 183 240 186 
rect 237 186 240 189 
rect 237 189 240 192 
rect 237 192 240 195 
rect 237 195 240 198 
rect 237 198 240 201 
rect 237 201 240 204 
rect 237 204 240 207 
rect 237 207 240 210 
rect 237 210 240 213 
rect 237 213 240 216 
rect 237 216 240 219 
rect 237 219 240 222 
rect 237 222 240 225 
rect 237 225 240 228 
rect 237 228 240 231 
rect 237 231 240 234 
rect 237 234 240 237 
rect 237 237 240 240 
rect 237 240 240 243 
rect 237 243 240 246 
rect 237 246 240 249 
rect 237 249 240 252 
rect 237 252 240 255 
rect 237 255 240 258 
rect 237 258 240 261 
rect 237 261 240 264 
rect 237 264 240 267 
rect 237 267 240 270 
rect 237 270 240 273 
rect 237 273 240 276 
rect 237 276 240 279 
rect 237 279 240 282 
rect 237 282 240 285 
rect 237 285 240 288 
rect 237 288 240 291 
rect 237 291 240 294 
rect 237 294 240 297 
rect 237 297 240 300 
rect 237 300 240 303 
rect 237 303 240 306 
rect 237 306 240 309 
rect 237 309 240 312 
rect 237 312 240 315 
rect 237 315 240 318 
rect 237 318 240 321 
rect 237 321 240 324 
rect 237 324 240 327 
rect 237 327 240 330 
rect 237 330 240 333 
rect 237 333 240 336 
rect 237 336 240 339 
rect 237 339 240 342 
rect 237 342 240 345 
rect 237 345 240 348 
rect 237 348 240 351 
rect 237 351 240 354 
rect 237 354 240 357 
rect 237 357 240 360 
rect 237 360 240 363 
rect 237 363 240 366 
rect 237 366 240 369 
rect 237 369 240 372 
rect 237 372 240 375 
rect 237 375 240 378 
rect 237 378 240 381 
rect 237 381 240 384 
rect 237 384 240 387 
rect 237 387 240 390 
rect 237 390 240 393 
rect 237 393 240 396 
rect 237 396 240 399 
rect 237 399 240 402 
rect 237 402 240 405 
rect 237 405 240 408 
rect 237 408 240 411 
rect 237 411 240 414 
rect 237 414 240 417 
rect 237 417 240 420 
rect 237 420 240 423 
rect 237 423 240 426 
rect 237 426 240 429 
rect 237 429 240 432 
rect 237 432 240 435 
rect 237 435 240 438 
rect 237 438 240 441 
rect 237 441 240 444 
rect 237 444 240 447 
rect 237 447 240 450 
rect 237 450 240 453 
rect 237 453 240 456 
rect 237 456 240 459 
rect 237 459 240 462 
rect 237 462 240 465 
rect 237 465 240 468 
rect 237 468 240 471 
rect 237 471 240 474 
rect 237 474 240 477 
rect 237 477 240 480 
rect 237 480 240 483 
rect 237 483 240 486 
rect 237 486 240 489 
rect 237 489 240 492 
rect 237 492 240 495 
rect 237 495 240 498 
rect 237 498 240 501 
rect 237 501 240 504 
rect 237 504 240 507 
rect 237 507 240 510 
rect 240 0 243 3 
rect 240 3 243 6 
rect 240 6 243 9 
rect 240 9 243 12 
rect 240 12 243 15 
rect 240 15 243 18 
rect 240 18 243 21 
rect 240 21 243 24 
rect 240 24 243 27 
rect 240 27 243 30 
rect 240 30 243 33 
rect 240 33 243 36 
rect 240 36 243 39 
rect 240 39 243 42 
rect 240 42 243 45 
rect 240 45 243 48 
rect 240 48 243 51 
rect 240 51 243 54 
rect 240 54 243 57 
rect 240 57 243 60 
rect 240 60 243 63 
rect 240 63 243 66 
rect 240 66 243 69 
rect 240 69 243 72 
rect 240 72 243 75 
rect 240 75 243 78 
rect 240 78 243 81 
rect 240 81 243 84 
rect 240 84 243 87 
rect 240 87 243 90 
rect 240 90 243 93 
rect 240 93 243 96 
rect 240 96 243 99 
rect 240 99 243 102 
rect 240 102 243 105 
rect 240 105 243 108 
rect 240 108 243 111 
rect 240 111 243 114 
rect 240 114 243 117 
rect 240 117 243 120 
rect 240 120 243 123 
rect 240 123 243 126 
rect 240 126 243 129 
rect 240 129 243 132 
rect 240 132 243 135 
rect 240 135 243 138 
rect 240 138 243 141 
rect 240 141 243 144 
rect 240 144 243 147 
rect 240 147 243 150 
rect 240 150 243 153 
rect 240 153 243 156 
rect 240 156 243 159 
rect 240 159 243 162 
rect 240 162 243 165 
rect 240 165 243 168 
rect 240 168 243 171 
rect 240 171 243 174 
rect 240 174 243 177 
rect 240 177 243 180 
rect 240 180 243 183 
rect 240 183 243 186 
rect 240 186 243 189 
rect 240 189 243 192 
rect 240 192 243 195 
rect 240 195 243 198 
rect 240 198 243 201 
rect 240 201 243 204 
rect 240 204 243 207 
rect 240 207 243 210 
rect 240 210 243 213 
rect 240 213 243 216 
rect 240 216 243 219 
rect 240 219 243 222 
rect 240 222 243 225 
rect 240 225 243 228 
rect 240 228 243 231 
rect 240 231 243 234 
rect 240 234 243 237 
rect 240 237 243 240 
rect 240 240 243 243 
rect 240 243 243 246 
rect 240 246 243 249 
rect 240 249 243 252 
rect 240 252 243 255 
rect 240 255 243 258 
rect 240 258 243 261 
rect 240 261 243 264 
rect 240 264 243 267 
rect 240 267 243 270 
rect 240 270 243 273 
rect 240 273 243 276 
rect 240 276 243 279 
rect 240 279 243 282 
rect 240 282 243 285 
rect 240 285 243 288 
rect 240 288 243 291 
rect 240 291 243 294 
rect 240 294 243 297 
rect 240 297 243 300 
rect 240 300 243 303 
rect 240 303 243 306 
rect 240 306 243 309 
rect 240 309 243 312 
rect 240 312 243 315 
rect 240 315 243 318 
rect 240 318 243 321 
rect 240 321 243 324 
rect 240 324 243 327 
rect 240 327 243 330 
rect 240 330 243 333 
rect 240 333 243 336 
rect 240 336 243 339 
rect 240 339 243 342 
rect 240 342 243 345 
rect 240 345 243 348 
rect 240 348 243 351 
rect 240 351 243 354 
rect 240 354 243 357 
rect 240 357 243 360 
rect 240 360 243 363 
rect 240 363 243 366 
rect 240 366 243 369 
rect 240 369 243 372 
rect 240 372 243 375 
rect 240 375 243 378 
rect 240 378 243 381 
rect 240 381 243 384 
rect 240 384 243 387 
rect 240 387 243 390 
rect 240 390 243 393 
rect 240 393 243 396 
rect 240 396 243 399 
rect 240 399 243 402 
rect 240 402 243 405 
rect 240 405 243 408 
rect 240 408 243 411 
rect 240 411 243 414 
rect 240 414 243 417 
rect 240 417 243 420 
rect 240 420 243 423 
rect 240 423 243 426 
rect 240 426 243 429 
rect 240 429 243 432 
rect 240 432 243 435 
rect 240 435 243 438 
rect 240 438 243 441 
rect 240 441 243 444 
rect 240 444 243 447 
rect 240 447 243 450 
rect 240 450 243 453 
rect 240 453 243 456 
rect 240 456 243 459 
rect 240 459 243 462 
rect 240 462 243 465 
rect 240 465 243 468 
rect 240 468 243 471 
rect 240 471 243 474 
rect 240 474 243 477 
rect 240 477 243 480 
rect 240 480 243 483 
rect 240 483 243 486 
rect 240 486 243 489 
rect 240 489 243 492 
rect 240 492 243 495 
rect 240 495 243 498 
rect 240 498 243 501 
rect 240 501 243 504 
rect 240 504 243 507 
rect 240 507 243 510 
rect 243 0 246 3 
rect 243 3 246 6 
rect 243 6 246 9 
rect 243 9 246 12 
rect 243 12 246 15 
rect 243 15 246 18 
rect 243 18 246 21 
rect 243 21 246 24 
rect 243 24 246 27 
rect 243 27 246 30 
rect 243 30 246 33 
rect 243 33 246 36 
rect 243 36 246 39 
rect 243 39 246 42 
rect 243 42 246 45 
rect 243 45 246 48 
rect 243 48 246 51 
rect 243 51 246 54 
rect 243 54 246 57 
rect 243 57 246 60 
rect 243 60 246 63 
rect 243 63 246 66 
rect 243 66 246 69 
rect 243 69 246 72 
rect 243 72 246 75 
rect 243 75 246 78 
rect 243 78 246 81 
rect 243 81 246 84 
rect 243 84 246 87 
rect 243 87 246 90 
rect 243 90 246 93 
rect 243 93 246 96 
rect 243 96 246 99 
rect 243 99 246 102 
rect 243 102 246 105 
rect 243 105 246 108 
rect 243 108 246 111 
rect 243 111 246 114 
rect 243 114 246 117 
rect 243 117 246 120 
rect 243 120 246 123 
rect 243 123 246 126 
rect 243 126 246 129 
rect 243 129 246 132 
rect 243 132 246 135 
rect 243 135 246 138 
rect 243 138 246 141 
rect 243 141 246 144 
rect 243 144 246 147 
rect 243 147 246 150 
rect 243 150 246 153 
rect 243 153 246 156 
rect 243 156 246 159 
rect 243 159 246 162 
rect 243 162 246 165 
rect 243 165 246 168 
rect 243 168 246 171 
rect 243 171 246 174 
rect 243 174 246 177 
rect 243 177 246 180 
rect 243 180 246 183 
rect 243 183 246 186 
rect 243 186 246 189 
rect 243 189 246 192 
rect 243 192 246 195 
rect 243 195 246 198 
rect 243 198 246 201 
rect 243 201 246 204 
rect 243 204 246 207 
rect 243 207 246 210 
rect 243 210 246 213 
rect 243 213 246 216 
rect 243 216 246 219 
rect 243 219 246 222 
rect 243 222 246 225 
rect 243 225 246 228 
rect 243 228 246 231 
rect 243 231 246 234 
rect 243 234 246 237 
rect 243 237 246 240 
rect 243 240 246 243 
rect 243 243 246 246 
rect 243 246 246 249 
rect 243 249 246 252 
rect 243 252 246 255 
rect 243 255 246 258 
rect 243 258 246 261 
rect 243 261 246 264 
rect 243 264 246 267 
rect 243 267 246 270 
rect 243 270 246 273 
rect 243 273 246 276 
rect 243 276 246 279 
rect 243 279 246 282 
rect 243 282 246 285 
rect 243 285 246 288 
rect 243 288 246 291 
rect 243 291 246 294 
rect 243 294 246 297 
rect 243 297 246 300 
rect 243 300 246 303 
rect 243 303 246 306 
rect 243 306 246 309 
rect 243 309 246 312 
rect 243 312 246 315 
rect 243 315 246 318 
rect 243 318 246 321 
rect 243 321 246 324 
rect 243 324 246 327 
rect 243 327 246 330 
rect 243 330 246 333 
rect 243 333 246 336 
rect 243 336 246 339 
rect 243 339 246 342 
rect 243 342 246 345 
rect 243 345 246 348 
rect 243 348 246 351 
rect 243 351 246 354 
rect 243 354 246 357 
rect 243 357 246 360 
rect 243 360 246 363 
rect 243 363 246 366 
rect 243 366 246 369 
rect 243 369 246 372 
rect 243 372 246 375 
rect 243 375 246 378 
rect 243 378 246 381 
rect 243 381 246 384 
rect 243 384 246 387 
rect 243 387 246 390 
rect 243 390 246 393 
rect 243 393 246 396 
rect 243 396 246 399 
rect 243 399 246 402 
rect 243 402 246 405 
rect 243 405 246 408 
rect 243 408 246 411 
rect 243 411 246 414 
rect 243 414 246 417 
rect 243 417 246 420 
rect 243 420 246 423 
rect 243 423 246 426 
rect 243 426 246 429 
rect 243 429 246 432 
rect 243 432 246 435 
rect 243 435 246 438 
rect 243 438 246 441 
rect 243 441 246 444 
rect 243 444 246 447 
rect 243 447 246 450 
rect 243 450 246 453 
rect 243 453 246 456 
rect 243 456 246 459 
rect 243 459 246 462 
rect 243 462 246 465 
rect 243 465 246 468 
rect 243 468 246 471 
rect 243 471 246 474 
rect 243 474 246 477 
rect 243 477 246 480 
rect 243 480 246 483 
rect 243 483 246 486 
rect 243 486 246 489 
rect 243 489 246 492 
rect 243 492 246 495 
rect 243 495 246 498 
rect 243 498 246 501 
rect 243 501 246 504 
rect 243 504 246 507 
rect 243 507 246 510 
rect 246 0 249 3 
rect 246 3 249 6 
rect 246 6 249 9 
rect 246 9 249 12 
rect 246 12 249 15 
rect 246 15 249 18 
rect 246 18 249 21 
rect 246 21 249 24 
rect 246 24 249 27 
rect 246 27 249 30 
rect 246 30 249 33 
rect 246 33 249 36 
rect 246 36 249 39 
rect 246 39 249 42 
rect 246 42 249 45 
rect 246 45 249 48 
rect 246 48 249 51 
rect 246 51 249 54 
rect 246 54 249 57 
rect 246 57 249 60 
rect 246 60 249 63 
rect 246 63 249 66 
rect 246 66 249 69 
rect 246 69 249 72 
rect 246 72 249 75 
rect 246 75 249 78 
rect 246 78 249 81 
rect 246 81 249 84 
rect 246 84 249 87 
rect 246 87 249 90 
rect 246 90 249 93 
rect 246 93 249 96 
rect 246 96 249 99 
rect 246 99 249 102 
rect 246 102 249 105 
rect 246 105 249 108 
rect 246 108 249 111 
rect 246 111 249 114 
rect 246 114 249 117 
rect 246 117 249 120 
rect 246 120 249 123 
rect 246 123 249 126 
rect 246 126 249 129 
rect 246 129 249 132 
rect 246 132 249 135 
rect 246 135 249 138 
rect 246 138 249 141 
rect 246 141 249 144 
rect 246 144 249 147 
rect 246 147 249 150 
rect 246 150 249 153 
rect 246 153 249 156 
rect 246 156 249 159 
rect 246 159 249 162 
rect 246 162 249 165 
rect 246 165 249 168 
rect 246 168 249 171 
rect 246 171 249 174 
rect 246 174 249 177 
rect 246 177 249 180 
rect 246 180 249 183 
rect 246 183 249 186 
rect 246 186 249 189 
rect 246 189 249 192 
rect 246 192 249 195 
rect 246 195 249 198 
rect 246 198 249 201 
rect 246 201 249 204 
rect 246 204 249 207 
rect 246 207 249 210 
rect 246 210 249 213 
rect 246 213 249 216 
rect 246 216 249 219 
rect 246 219 249 222 
rect 246 222 249 225 
rect 246 225 249 228 
rect 246 228 249 231 
rect 246 231 249 234 
rect 246 234 249 237 
rect 246 237 249 240 
rect 246 240 249 243 
rect 246 243 249 246 
rect 246 246 249 249 
rect 246 249 249 252 
rect 246 252 249 255 
rect 246 255 249 258 
rect 246 258 249 261 
rect 246 261 249 264 
rect 246 264 249 267 
rect 246 267 249 270 
rect 246 270 249 273 
rect 246 273 249 276 
rect 246 276 249 279 
rect 246 279 249 282 
rect 246 282 249 285 
rect 246 285 249 288 
rect 246 288 249 291 
rect 246 291 249 294 
rect 246 294 249 297 
rect 246 297 249 300 
rect 246 300 249 303 
rect 246 303 249 306 
rect 246 306 249 309 
rect 246 309 249 312 
rect 246 312 249 315 
rect 246 315 249 318 
rect 246 318 249 321 
rect 246 321 249 324 
rect 246 324 249 327 
rect 246 327 249 330 
rect 246 330 249 333 
rect 246 333 249 336 
rect 246 336 249 339 
rect 246 339 249 342 
rect 246 342 249 345 
rect 246 345 249 348 
rect 246 348 249 351 
rect 246 351 249 354 
rect 246 354 249 357 
rect 246 357 249 360 
rect 246 360 249 363 
rect 246 363 249 366 
rect 246 366 249 369 
rect 246 369 249 372 
rect 246 372 249 375 
rect 246 375 249 378 
rect 246 378 249 381 
rect 246 381 249 384 
rect 246 384 249 387 
rect 246 387 249 390 
rect 246 390 249 393 
rect 246 393 249 396 
rect 246 396 249 399 
rect 246 399 249 402 
rect 246 402 249 405 
rect 246 405 249 408 
rect 246 408 249 411 
rect 246 411 249 414 
rect 246 414 249 417 
rect 246 417 249 420 
rect 246 420 249 423 
rect 246 423 249 426 
rect 246 426 249 429 
rect 246 429 249 432 
rect 246 432 249 435 
rect 246 435 249 438 
rect 246 438 249 441 
rect 246 441 249 444 
rect 246 444 249 447 
rect 246 447 249 450 
rect 246 450 249 453 
rect 246 453 249 456 
rect 246 456 249 459 
rect 246 459 249 462 
rect 246 462 249 465 
rect 246 465 249 468 
rect 246 468 249 471 
rect 246 471 249 474 
rect 246 474 249 477 
rect 246 477 249 480 
rect 246 480 249 483 
rect 246 483 249 486 
rect 246 486 249 489 
rect 246 489 249 492 
rect 246 492 249 495 
rect 246 495 249 498 
rect 246 498 249 501 
rect 246 501 249 504 
rect 246 504 249 507 
rect 246 507 249 510 
rect 249 0 252 3 
rect 249 3 252 6 
rect 249 6 252 9 
rect 249 9 252 12 
rect 249 12 252 15 
rect 249 15 252 18 
rect 249 18 252 21 
rect 249 21 252 24 
rect 249 24 252 27 
rect 249 27 252 30 
rect 249 30 252 33 
rect 249 33 252 36 
rect 249 36 252 39 
rect 249 39 252 42 
rect 249 42 252 45 
rect 249 45 252 48 
rect 249 48 252 51 
rect 249 51 252 54 
rect 249 54 252 57 
rect 249 57 252 60 
rect 249 60 252 63 
rect 249 63 252 66 
rect 249 66 252 69 
rect 249 69 252 72 
rect 249 72 252 75 
rect 249 75 252 78 
rect 249 78 252 81 
rect 249 81 252 84 
rect 249 84 252 87 
rect 249 87 252 90 
rect 249 90 252 93 
rect 249 93 252 96 
rect 249 96 252 99 
rect 249 99 252 102 
rect 249 102 252 105 
rect 249 105 252 108 
rect 249 108 252 111 
rect 249 111 252 114 
rect 249 114 252 117 
rect 249 117 252 120 
rect 249 120 252 123 
rect 249 123 252 126 
rect 249 126 252 129 
rect 249 129 252 132 
rect 249 132 252 135 
rect 249 135 252 138 
rect 249 138 252 141 
rect 249 141 252 144 
rect 249 144 252 147 
rect 249 147 252 150 
rect 249 150 252 153 
rect 249 153 252 156 
rect 249 156 252 159 
rect 249 159 252 162 
rect 249 162 252 165 
rect 249 165 252 168 
rect 249 168 252 171 
rect 249 171 252 174 
rect 249 174 252 177 
rect 249 177 252 180 
rect 249 180 252 183 
rect 249 183 252 186 
rect 249 186 252 189 
rect 249 189 252 192 
rect 249 192 252 195 
rect 249 195 252 198 
rect 249 198 252 201 
rect 249 201 252 204 
rect 249 204 252 207 
rect 249 207 252 210 
rect 249 210 252 213 
rect 249 213 252 216 
rect 249 216 252 219 
rect 249 219 252 222 
rect 249 222 252 225 
rect 249 225 252 228 
rect 249 228 252 231 
rect 249 231 252 234 
rect 249 234 252 237 
rect 249 237 252 240 
rect 249 240 252 243 
rect 249 243 252 246 
rect 249 246 252 249 
rect 249 249 252 252 
rect 249 252 252 255 
rect 249 255 252 258 
rect 249 258 252 261 
rect 249 261 252 264 
rect 249 264 252 267 
rect 249 267 252 270 
rect 249 270 252 273 
rect 249 273 252 276 
rect 249 276 252 279 
rect 249 279 252 282 
rect 249 282 252 285 
rect 249 285 252 288 
rect 249 288 252 291 
rect 249 291 252 294 
rect 249 294 252 297 
rect 249 297 252 300 
rect 249 300 252 303 
rect 249 303 252 306 
rect 249 306 252 309 
rect 249 309 252 312 
rect 249 312 252 315 
rect 249 315 252 318 
rect 249 318 252 321 
rect 249 321 252 324 
rect 249 324 252 327 
rect 249 327 252 330 
rect 249 330 252 333 
rect 249 333 252 336 
rect 249 336 252 339 
rect 249 339 252 342 
rect 249 342 252 345 
rect 249 345 252 348 
rect 249 348 252 351 
rect 249 351 252 354 
rect 249 354 252 357 
rect 249 357 252 360 
rect 249 360 252 363 
rect 249 363 252 366 
rect 249 366 252 369 
rect 249 369 252 372 
rect 249 372 252 375 
rect 249 375 252 378 
rect 249 378 252 381 
rect 249 381 252 384 
rect 249 384 252 387 
rect 249 387 252 390 
rect 249 390 252 393 
rect 249 393 252 396 
rect 249 396 252 399 
rect 249 399 252 402 
rect 249 402 252 405 
rect 249 405 252 408 
rect 249 408 252 411 
rect 249 411 252 414 
rect 249 414 252 417 
rect 249 417 252 420 
rect 249 420 252 423 
rect 249 423 252 426 
rect 249 426 252 429 
rect 249 429 252 432 
rect 249 432 252 435 
rect 249 435 252 438 
rect 249 438 252 441 
rect 249 441 252 444 
rect 249 444 252 447 
rect 249 447 252 450 
rect 249 450 252 453 
rect 249 453 252 456 
rect 249 456 252 459 
rect 249 459 252 462 
rect 249 462 252 465 
rect 249 465 252 468 
rect 249 468 252 471 
rect 249 471 252 474 
rect 249 474 252 477 
rect 249 477 252 480 
rect 249 480 252 483 
rect 249 483 252 486 
rect 249 486 252 489 
rect 249 489 252 492 
rect 249 492 252 495 
rect 249 495 252 498 
rect 249 498 252 501 
rect 249 501 252 504 
rect 249 504 252 507 
rect 249 507 252 510 
rect 252 0 255 3 
rect 252 3 255 6 
rect 252 6 255 9 
rect 252 9 255 12 
rect 252 12 255 15 
rect 252 15 255 18 
rect 252 18 255 21 
rect 252 21 255 24 
rect 252 24 255 27 
rect 252 27 255 30 
rect 252 30 255 33 
rect 252 33 255 36 
rect 252 36 255 39 
rect 252 39 255 42 
rect 252 42 255 45 
rect 252 45 255 48 
rect 252 48 255 51 
rect 252 51 255 54 
rect 252 54 255 57 
rect 252 57 255 60 
rect 252 60 255 63 
rect 252 63 255 66 
rect 252 66 255 69 
rect 252 69 255 72 
rect 252 72 255 75 
rect 252 75 255 78 
rect 252 78 255 81 
rect 252 81 255 84 
rect 252 84 255 87 
rect 252 87 255 90 
rect 252 90 255 93 
rect 252 93 255 96 
rect 252 96 255 99 
rect 252 99 255 102 
rect 252 102 255 105 
rect 252 105 255 108 
rect 252 108 255 111 
rect 252 111 255 114 
rect 252 114 255 117 
rect 252 117 255 120 
rect 252 120 255 123 
rect 252 123 255 126 
rect 252 126 255 129 
rect 252 129 255 132 
rect 252 132 255 135 
rect 252 135 255 138 
rect 252 138 255 141 
rect 252 141 255 144 
rect 252 144 255 147 
rect 252 147 255 150 
rect 252 150 255 153 
rect 252 153 255 156 
rect 252 156 255 159 
rect 252 159 255 162 
rect 252 162 255 165 
rect 252 165 255 168 
rect 252 168 255 171 
rect 252 171 255 174 
rect 252 174 255 177 
rect 252 177 255 180 
rect 252 180 255 183 
rect 252 183 255 186 
rect 252 186 255 189 
rect 252 189 255 192 
rect 252 192 255 195 
rect 252 195 255 198 
rect 252 198 255 201 
rect 252 201 255 204 
rect 252 204 255 207 
rect 252 207 255 210 
rect 252 210 255 213 
rect 252 213 255 216 
rect 252 216 255 219 
rect 252 219 255 222 
rect 252 222 255 225 
rect 252 225 255 228 
rect 252 228 255 231 
rect 252 231 255 234 
rect 252 234 255 237 
rect 252 237 255 240 
rect 252 240 255 243 
rect 252 243 255 246 
rect 252 246 255 249 
rect 252 249 255 252 
rect 252 252 255 255 
rect 252 255 255 258 
rect 252 258 255 261 
rect 252 261 255 264 
rect 252 264 255 267 
rect 252 267 255 270 
rect 252 270 255 273 
rect 252 273 255 276 
rect 252 276 255 279 
rect 252 279 255 282 
rect 252 282 255 285 
rect 252 285 255 288 
rect 252 288 255 291 
rect 252 291 255 294 
rect 252 294 255 297 
rect 252 297 255 300 
rect 252 300 255 303 
rect 252 303 255 306 
rect 252 306 255 309 
rect 252 309 255 312 
rect 252 312 255 315 
rect 252 315 255 318 
rect 252 318 255 321 
rect 252 321 255 324 
rect 252 324 255 327 
rect 252 327 255 330 
rect 252 330 255 333 
rect 252 333 255 336 
rect 252 336 255 339 
rect 252 339 255 342 
rect 252 342 255 345 
rect 252 345 255 348 
rect 252 348 255 351 
rect 252 351 255 354 
rect 252 354 255 357 
rect 252 357 255 360 
rect 252 360 255 363 
rect 252 363 255 366 
rect 252 366 255 369 
rect 252 369 255 372 
rect 252 372 255 375 
rect 252 375 255 378 
rect 252 378 255 381 
rect 252 381 255 384 
rect 252 384 255 387 
rect 252 387 255 390 
rect 252 390 255 393 
rect 252 393 255 396 
rect 252 396 255 399 
rect 252 399 255 402 
rect 252 402 255 405 
rect 252 405 255 408 
rect 252 408 255 411 
rect 252 411 255 414 
rect 252 414 255 417 
rect 252 417 255 420 
rect 252 420 255 423 
rect 252 423 255 426 
rect 252 426 255 429 
rect 252 429 255 432 
rect 252 432 255 435 
rect 252 435 255 438 
rect 252 438 255 441 
rect 252 441 255 444 
rect 252 444 255 447 
rect 252 447 255 450 
rect 252 450 255 453 
rect 252 453 255 456 
rect 252 456 255 459 
rect 252 459 255 462 
rect 252 462 255 465 
rect 252 465 255 468 
rect 252 468 255 471 
rect 252 471 255 474 
rect 252 474 255 477 
rect 252 477 255 480 
rect 252 480 255 483 
rect 252 483 255 486 
rect 252 486 255 489 
rect 252 489 255 492 
rect 252 492 255 495 
rect 252 495 255 498 
rect 252 498 255 501 
rect 252 501 255 504 
rect 252 504 255 507 
rect 252 507 255 510 
rect 255 0 258 3 
rect 255 3 258 6 
rect 255 6 258 9 
rect 255 9 258 12 
rect 255 12 258 15 
rect 255 15 258 18 
rect 255 18 258 21 
rect 255 21 258 24 
rect 255 24 258 27 
rect 255 27 258 30 
rect 255 30 258 33 
rect 255 33 258 36 
rect 255 36 258 39 
rect 255 39 258 42 
rect 255 42 258 45 
rect 255 45 258 48 
rect 255 48 258 51 
rect 255 51 258 54 
rect 255 54 258 57 
rect 255 57 258 60 
rect 255 60 258 63 
rect 255 63 258 66 
rect 255 66 258 69 
rect 255 69 258 72 
rect 255 72 258 75 
rect 255 75 258 78 
rect 255 78 258 81 
rect 255 81 258 84 
rect 255 84 258 87 
rect 255 87 258 90 
rect 255 90 258 93 
rect 255 93 258 96 
rect 255 96 258 99 
rect 255 99 258 102 
rect 255 102 258 105 
rect 255 105 258 108 
rect 255 108 258 111 
rect 255 111 258 114 
rect 255 114 258 117 
rect 255 117 258 120 
rect 255 120 258 123 
rect 255 123 258 126 
rect 255 126 258 129 
rect 255 129 258 132 
rect 255 132 258 135 
rect 255 135 258 138 
rect 255 138 258 141 
rect 255 141 258 144 
rect 255 144 258 147 
rect 255 147 258 150 
rect 255 150 258 153 
rect 255 153 258 156 
rect 255 156 258 159 
rect 255 159 258 162 
rect 255 162 258 165 
rect 255 165 258 168 
rect 255 168 258 171 
rect 255 171 258 174 
rect 255 174 258 177 
rect 255 177 258 180 
rect 255 180 258 183 
rect 255 183 258 186 
rect 255 186 258 189 
rect 255 189 258 192 
rect 255 192 258 195 
rect 255 195 258 198 
rect 255 198 258 201 
rect 255 201 258 204 
rect 255 204 258 207 
rect 255 207 258 210 
rect 255 210 258 213 
rect 255 213 258 216 
rect 255 216 258 219 
rect 255 219 258 222 
rect 255 222 258 225 
rect 255 225 258 228 
rect 255 228 258 231 
rect 255 231 258 234 
rect 255 234 258 237 
rect 255 237 258 240 
rect 255 240 258 243 
rect 255 243 258 246 
rect 255 246 258 249 
rect 255 249 258 252 
rect 255 252 258 255 
rect 255 255 258 258 
rect 255 258 258 261 
rect 255 261 258 264 
rect 255 264 258 267 
rect 255 267 258 270 
rect 255 270 258 273 
rect 255 273 258 276 
rect 255 276 258 279 
rect 255 279 258 282 
rect 255 282 258 285 
rect 255 285 258 288 
rect 255 288 258 291 
rect 255 291 258 294 
rect 255 294 258 297 
rect 255 297 258 300 
rect 255 300 258 303 
rect 255 303 258 306 
rect 255 306 258 309 
rect 255 309 258 312 
rect 255 312 258 315 
rect 255 315 258 318 
rect 255 318 258 321 
rect 255 321 258 324 
rect 255 324 258 327 
rect 255 327 258 330 
rect 255 330 258 333 
rect 255 333 258 336 
rect 255 336 258 339 
rect 255 339 258 342 
rect 255 342 258 345 
rect 255 345 258 348 
rect 255 348 258 351 
rect 255 351 258 354 
rect 255 354 258 357 
rect 255 357 258 360 
rect 255 360 258 363 
rect 255 363 258 366 
rect 255 366 258 369 
rect 255 369 258 372 
rect 255 372 258 375 
rect 255 375 258 378 
rect 255 378 258 381 
rect 255 381 258 384 
rect 255 384 258 387 
rect 255 387 258 390 
rect 255 390 258 393 
rect 255 393 258 396 
rect 255 396 258 399 
rect 255 399 258 402 
rect 255 402 258 405 
rect 255 405 258 408 
rect 255 408 258 411 
rect 255 411 258 414 
rect 255 414 258 417 
rect 255 417 258 420 
rect 255 420 258 423 
rect 255 423 258 426 
rect 255 426 258 429 
rect 255 429 258 432 
rect 255 432 258 435 
rect 255 435 258 438 
rect 255 438 258 441 
rect 255 441 258 444 
rect 255 444 258 447 
rect 255 447 258 450 
rect 255 450 258 453 
rect 255 453 258 456 
rect 255 456 258 459 
rect 255 459 258 462 
rect 255 462 258 465 
rect 255 465 258 468 
rect 255 468 258 471 
rect 255 471 258 474 
rect 255 474 258 477 
rect 255 477 258 480 
rect 255 480 258 483 
rect 255 483 258 486 
rect 255 486 258 489 
rect 255 489 258 492 
rect 255 492 258 495 
rect 255 495 258 498 
rect 255 498 258 501 
rect 255 501 258 504 
rect 255 504 258 507 
rect 255 507 258 510 
rect 258 0 261 3 
rect 258 3 261 6 
rect 258 6 261 9 
rect 258 9 261 12 
rect 258 12 261 15 
rect 258 15 261 18 
rect 258 18 261 21 
rect 258 21 261 24 
rect 258 24 261 27 
rect 258 27 261 30 
rect 258 30 261 33 
rect 258 33 261 36 
rect 258 36 261 39 
rect 258 39 261 42 
rect 258 42 261 45 
rect 258 45 261 48 
rect 258 48 261 51 
rect 258 51 261 54 
rect 258 54 261 57 
rect 258 57 261 60 
rect 258 60 261 63 
rect 258 63 261 66 
rect 258 66 261 69 
rect 258 69 261 72 
rect 258 72 261 75 
rect 258 75 261 78 
rect 258 78 261 81 
rect 258 81 261 84 
rect 258 84 261 87 
rect 258 87 261 90 
rect 258 90 261 93 
rect 258 93 261 96 
rect 258 96 261 99 
rect 258 99 261 102 
rect 258 102 261 105 
rect 258 105 261 108 
rect 258 108 261 111 
rect 258 111 261 114 
rect 258 114 261 117 
rect 258 117 261 120 
rect 258 120 261 123 
rect 258 123 261 126 
rect 258 126 261 129 
rect 258 129 261 132 
rect 258 132 261 135 
rect 258 135 261 138 
rect 258 138 261 141 
rect 258 141 261 144 
rect 258 144 261 147 
rect 258 147 261 150 
rect 258 150 261 153 
rect 258 153 261 156 
rect 258 156 261 159 
rect 258 159 261 162 
rect 258 162 261 165 
rect 258 165 261 168 
rect 258 168 261 171 
rect 258 171 261 174 
rect 258 174 261 177 
rect 258 177 261 180 
rect 258 180 261 183 
rect 258 183 261 186 
rect 258 186 261 189 
rect 258 189 261 192 
rect 258 192 261 195 
rect 258 195 261 198 
rect 258 198 261 201 
rect 258 201 261 204 
rect 258 204 261 207 
rect 258 207 261 210 
rect 258 210 261 213 
rect 258 213 261 216 
rect 258 216 261 219 
rect 258 219 261 222 
rect 258 222 261 225 
rect 258 225 261 228 
rect 258 228 261 231 
rect 258 231 261 234 
rect 258 234 261 237 
rect 258 237 261 240 
rect 258 240 261 243 
rect 258 243 261 246 
rect 258 246 261 249 
rect 258 249 261 252 
rect 258 252 261 255 
rect 258 255 261 258 
rect 258 258 261 261 
rect 258 261 261 264 
rect 258 264 261 267 
rect 258 267 261 270 
rect 258 270 261 273 
rect 258 273 261 276 
rect 258 276 261 279 
rect 258 279 261 282 
rect 258 282 261 285 
rect 258 285 261 288 
rect 258 288 261 291 
rect 258 291 261 294 
rect 258 294 261 297 
rect 258 297 261 300 
rect 258 300 261 303 
rect 258 303 261 306 
rect 258 306 261 309 
rect 258 309 261 312 
rect 258 312 261 315 
rect 258 315 261 318 
rect 258 318 261 321 
rect 258 321 261 324 
rect 258 324 261 327 
rect 258 327 261 330 
rect 258 330 261 333 
rect 258 333 261 336 
rect 258 336 261 339 
rect 258 339 261 342 
rect 258 342 261 345 
rect 258 345 261 348 
rect 258 348 261 351 
rect 258 351 261 354 
rect 258 354 261 357 
rect 258 357 261 360 
rect 258 360 261 363 
rect 258 363 261 366 
rect 258 366 261 369 
rect 258 369 261 372 
rect 258 372 261 375 
rect 258 375 261 378 
rect 258 378 261 381 
rect 258 381 261 384 
rect 258 384 261 387 
rect 258 387 261 390 
rect 258 390 261 393 
rect 258 393 261 396 
rect 258 396 261 399 
rect 258 399 261 402 
rect 258 402 261 405 
rect 258 405 261 408 
rect 258 408 261 411 
rect 258 411 261 414 
rect 258 414 261 417 
rect 258 417 261 420 
rect 258 420 261 423 
rect 258 423 261 426 
rect 258 426 261 429 
rect 258 429 261 432 
rect 258 432 261 435 
rect 258 435 261 438 
rect 258 438 261 441 
rect 258 441 261 444 
rect 258 444 261 447 
rect 258 447 261 450 
rect 258 450 261 453 
rect 258 453 261 456 
rect 258 456 261 459 
rect 258 459 261 462 
rect 258 462 261 465 
rect 258 465 261 468 
rect 258 468 261 471 
rect 258 471 261 474 
rect 258 474 261 477 
rect 258 477 261 480 
rect 258 480 261 483 
rect 258 483 261 486 
rect 258 486 261 489 
rect 258 489 261 492 
rect 258 492 261 495 
rect 258 495 261 498 
rect 258 498 261 501 
rect 258 501 261 504 
rect 258 504 261 507 
rect 258 507 261 510 
rect 261 0 264 3 
rect 261 3 264 6 
rect 261 6 264 9 
rect 261 9 264 12 
rect 261 12 264 15 
rect 261 15 264 18 
rect 261 18 264 21 
rect 261 21 264 24 
rect 261 24 264 27 
rect 261 27 264 30 
rect 261 30 264 33 
rect 261 33 264 36 
rect 261 36 264 39 
rect 261 39 264 42 
rect 261 42 264 45 
rect 261 45 264 48 
rect 261 48 264 51 
rect 261 51 264 54 
rect 261 54 264 57 
rect 261 57 264 60 
rect 261 60 264 63 
rect 261 63 264 66 
rect 261 66 264 69 
rect 261 69 264 72 
rect 261 72 264 75 
rect 261 75 264 78 
rect 261 78 264 81 
rect 261 81 264 84 
rect 261 84 264 87 
rect 261 87 264 90 
rect 261 90 264 93 
rect 261 93 264 96 
rect 261 96 264 99 
rect 261 99 264 102 
rect 261 102 264 105 
rect 261 105 264 108 
rect 261 108 264 111 
rect 261 111 264 114 
rect 261 114 264 117 
rect 261 117 264 120 
rect 261 120 264 123 
rect 261 123 264 126 
rect 261 126 264 129 
rect 261 129 264 132 
rect 261 132 264 135 
rect 261 135 264 138 
rect 261 138 264 141 
rect 261 141 264 144 
rect 261 144 264 147 
rect 261 147 264 150 
rect 261 150 264 153 
rect 261 153 264 156 
rect 261 156 264 159 
rect 261 159 264 162 
rect 261 162 264 165 
rect 261 165 264 168 
rect 261 168 264 171 
rect 261 171 264 174 
rect 261 174 264 177 
rect 261 177 264 180 
rect 261 180 264 183 
rect 261 183 264 186 
rect 261 186 264 189 
rect 261 189 264 192 
rect 261 192 264 195 
rect 261 195 264 198 
rect 261 198 264 201 
rect 261 201 264 204 
rect 261 204 264 207 
rect 261 207 264 210 
rect 261 210 264 213 
rect 261 213 264 216 
rect 261 216 264 219 
rect 261 219 264 222 
rect 261 222 264 225 
rect 261 225 264 228 
rect 261 228 264 231 
rect 261 231 264 234 
rect 261 234 264 237 
rect 261 237 264 240 
rect 261 240 264 243 
rect 261 243 264 246 
rect 261 246 264 249 
rect 261 249 264 252 
rect 261 252 264 255 
rect 261 255 264 258 
rect 261 258 264 261 
rect 261 261 264 264 
rect 261 264 264 267 
rect 261 267 264 270 
rect 261 270 264 273 
rect 261 273 264 276 
rect 261 276 264 279 
rect 261 279 264 282 
rect 261 282 264 285 
rect 261 285 264 288 
rect 261 288 264 291 
rect 261 291 264 294 
rect 261 294 264 297 
rect 261 297 264 300 
rect 261 300 264 303 
rect 261 303 264 306 
rect 261 306 264 309 
rect 261 309 264 312 
rect 261 312 264 315 
rect 261 315 264 318 
rect 261 318 264 321 
rect 261 321 264 324 
rect 261 324 264 327 
rect 261 327 264 330 
rect 261 330 264 333 
rect 261 333 264 336 
rect 261 336 264 339 
rect 261 339 264 342 
rect 261 342 264 345 
rect 261 345 264 348 
rect 261 348 264 351 
rect 261 351 264 354 
rect 261 354 264 357 
rect 261 357 264 360 
rect 261 360 264 363 
rect 261 363 264 366 
rect 261 366 264 369 
rect 261 369 264 372 
rect 261 372 264 375 
rect 261 375 264 378 
rect 261 378 264 381 
rect 261 381 264 384 
rect 261 384 264 387 
rect 261 387 264 390 
rect 261 390 264 393 
rect 261 393 264 396 
rect 261 396 264 399 
rect 261 399 264 402 
rect 261 402 264 405 
rect 261 405 264 408 
rect 261 408 264 411 
rect 261 411 264 414 
rect 261 414 264 417 
rect 261 417 264 420 
rect 261 420 264 423 
rect 261 423 264 426 
rect 261 426 264 429 
rect 261 429 264 432 
rect 261 432 264 435 
rect 261 435 264 438 
rect 261 438 264 441 
rect 261 441 264 444 
rect 261 444 264 447 
rect 261 447 264 450 
rect 261 450 264 453 
rect 261 453 264 456 
rect 261 456 264 459 
rect 261 459 264 462 
rect 261 462 264 465 
rect 261 465 264 468 
rect 261 468 264 471 
rect 261 471 264 474 
rect 261 474 264 477 
rect 261 477 264 480 
rect 261 480 264 483 
rect 261 483 264 486 
rect 261 486 264 489 
rect 261 489 264 492 
rect 261 492 264 495 
rect 261 495 264 498 
rect 261 498 264 501 
rect 261 501 264 504 
rect 261 504 264 507 
rect 261 507 264 510 
rect 264 0 267 3 
rect 264 3 267 6 
rect 264 6 267 9 
rect 264 9 267 12 
rect 264 12 267 15 
rect 264 15 267 18 
rect 264 18 267 21 
rect 264 21 267 24 
rect 264 24 267 27 
rect 264 27 267 30 
rect 264 30 267 33 
rect 264 33 267 36 
rect 264 36 267 39 
rect 264 39 267 42 
rect 264 42 267 45 
rect 264 45 267 48 
rect 264 48 267 51 
rect 264 51 267 54 
rect 264 54 267 57 
rect 264 57 267 60 
rect 264 60 267 63 
rect 264 63 267 66 
rect 264 66 267 69 
rect 264 69 267 72 
rect 264 72 267 75 
rect 264 75 267 78 
rect 264 78 267 81 
rect 264 81 267 84 
rect 264 84 267 87 
rect 264 87 267 90 
rect 264 90 267 93 
rect 264 93 267 96 
rect 264 96 267 99 
rect 264 99 267 102 
rect 264 102 267 105 
rect 264 105 267 108 
rect 264 108 267 111 
rect 264 111 267 114 
rect 264 114 267 117 
rect 264 117 267 120 
rect 264 120 267 123 
rect 264 123 267 126 
rect 264 126 267 129 
rect 264 129 267 132 
rect 264 132 267 135 
rect 264 135 267 138 
rect 264 138 267 141 
rect 264 141 267 144 
rect 264 144 267 147 
rect 264 147 267 150 
rect 264 150 267 153 
rect 264 153 267 156 
rect 264 156 267 159 
rect 264 159 267 162 
rect 264 162 267 165 
rect 264 165 267 168 
rect 264 168 267 171 
rect 264 171 267 174 
rect 264 174 267 177 
rect 264 177 267 180 
rect 264 180 267 183 
rect 264 183 267 186 
rect 264 186 267 189 
rect 264 189 267 192 
rect 264 192 267 195 
rect 264 195 267 198 
rect 264 198 267 201 
rect 264 201 267 204 
rect 264 204 267 207 
rect 264 207 267 210 
rect 264 210 267 213 
rect 264 213 267 216 
rect 264 216 267 219 
rect 264 219 267 222 
rect 264 222 267 225 
rect 264 225 267 228 
rect 264 228 267 231 
rect 264 231 267 234 
rect 264 234 267 237 
rect 264 237 267 240 
rect 264 240 267 243 
rect 264 243 267 246 
rect 264 246 267 249 
rect 264 249 267 252 
rect 264 252 267 255 
rect 264 255 267 258 
rect 264 258 267 261 
rect 264 261 267 264 
rect 264 264 267 267 
rect 264 267 267 270 
rect 264 270 267 273 
rect 264 273 267 276 
rect 264 276 267 279 
rect 264 279 267 282 
rect 264 282 267 285 
rect 264 285 267 288 
rect 264 288 267 291 
rect 264 291 267 294 
rect 264 294 267 297 
rect 264 297 267 300 
rect 264 300 267 303 
rect 264 303 267 306 
rect 264 306 267 309 
rect 264 309 267 312 
rect 264 312 267 315 
rect 264 315 267 318 
rect 264 318 267 321 
rect 264 321 267 324 
rect 264 324 267 327 
rect 264 327 267 330 
rect 264 330 267 333 
rect 264 333 267 336 
rect 264 336 267 339 
rect 264 339 267 342 
rect 264 342 267 345 
rect 264 345 267 348 
rect 264 348 267 351 
rect 264 351 267 354 
rect 264 354 267 357 
rect 264 357 267 360 
rect 264 360 267 363 
rect 264 363 267 366 
rect 264 366 267 369 
rect 264 369 267 372 
rect 264 372 267 375 
rect 264 375 267 378 
rect 264 378 267 381 
rect 264 381 267 384 
rect 264 384 267 387 
rect 264 387 267 390 
rect 264 390 267 393 
rect 264 393 267 396 
rect 264 396 267 399 
rect 264 399 267 402 
rect 264 402 267 405 
rect 264 405 267 408 
rect 264 408 267 411 
rect 264 411 267 414 
rect 264 414 267 417 
rect 264 417 267 420 
rect 264 420 267 423 
rect 264 423 267 426 
rect 264 426 267 429 
rect 264 429 267 432 
rect 264 432 267 435 
rect 264 435 267 438 
rect 264 438 267 441 
rect 264 441 267 444 
rect 264 444 267 447 
rect 264 447 267 450 
rect 264 450 267 453 
rect 264 453 267 456 
rect 264 456 267 459 
rect 264 459 267 462 
rect 264 462 267 465 
rect 264 465 267 468 
rect 264 468 267 471 
rect 264 471 267 474 
rect 264 474 267 477 
rect 264 477 267 480 
rect 264 480 267 483 
rect 264 483 267 486 
rect 264 486 267 489 
rect 264 489 267 492 
rect 264 492 267 495 
rect 264 495 267 498 
rect 264 498 267 501 
rect 264 501 267 504 
rect 264 504 267 507 
rect 264 507 267 510 
rect 267 0 270 3 
rect 267 3 270 6 
rect 267 6 270 9 
rect 267 9 270 12 
rect 267 12 270 15 
rect 267 15 270 18 
rect 267 18 270 21 
rect 267 21 270 24 
rect 267 24 270 27 
rect 267 27 270 30 
rect 267 30 270 33 
rect 267 33 270 36 
rect 267 36 270 39 
rect 267 39 270 42 
rect 267 42 270 45 
rect 267 45 270 48 
rect 267 48 270 51 
rect 267 51 270 54 
rect 267 54 270 57 
rect 267 57 270 60 
rect 267 60 270 63 
rect 267 63 270 66 
rect 267 66 270 69 
rect 267 69 270 72 
rect 267 72 270 75 
rect 267 75 270 78 
rect 267 78 270 81 
rect 267 81 270 84 
rect 267 84 270 87 
rect 267 87 270 90 
rect 267 90 270 93 
rect 267 93 270 96 
rect 267 96 270 99 
rect 267 99 270 102 
rect 267 102 270 105 
rect 267 105 270 108 
rect 267 108 270 111 
rect 267 111 270 114 
rect 267 114 270 117 
rect 267 117 270 120 
rect 267 120 270 123 
rect 267 123 270 126 
rect 267 126 270 129 
rect 267 129 270 132 
rect 267 132 270 135 
rect 267 135 270 138 
rect 267 138 270 141 
rect 267 141 270 144 
rect 267 144 270 147 
rect 267 147 270 150 
rect 267 150 270 153 
rect 267 153 270 156 
rect 267 156 270 159 
rect 267 159 270 162 
rect 267 162 270 165 
rect 267 165 270 168 
rect 267 168 270 171 
rect 267 171 270 174 
rect 267 174 270 177 
rect 267 177 270 180 
rect 267 180 270 183 
rect 267 183 270 186 
rect 267 186 270 189 
rect 267 189 270 192 
rect 267 192 270 195 
rect 267 195 270 198 
rect 267 198 270 201 
rect 267 201 270 204 
rect 267 204 270 207 
rect 267 207 270 210 
rect 267 210 270 213 
rect 267 213 270 216 
rect 267 216 270 219 
rect 267 219 270 222 
rect 267 222 270 225 
rect 267 225 270 228 
rect 267 228 270 231 
rect 267 231 270 234 
rect 267 234 270 237 
rect 267 237 270 240 
rect 267 240 270 243 
rect 267 243 270 246 
rect 267 246 270 249 
rect 267 249 270 252 
rect 267 252 270 255 
rect 267 255 270 258 
rect 267 258 270 261 
rect 267 261 270 264 
rect 267 264 270 267 
rect 267 267 270 270 
rect 267 270 270 273 
rect 267 273 270 276 
rect 267 276 270 279 
rect 267 279 270 282 
rect 267 282 270 285 
rect 267 285 270 288 
rect 267 288 270 291 
rect 267 291 270 294 
rect 267 294 270 297 
rect 267 297 270 300 
rect 267 300 270 303 
rect 267 303 270 306 
rect 267 306 270 309 
rect 267 309 270 312 
rect 267 312 270 315 
rect 267 315 270 318 
rect 267 318 270 321 
rect 267 321 270 324 
rect 267 324 270 327 
rect 267 327 270 330 
rect 267 330 270 333 
rect 267 333 270 336 
rect 267 336 270 339 
rect 267 339 270 342 
rect 267 342 270 345 
rect 267 345 270 348 
rect 267 348 270 351 
rect 267 351 270 354 
rect 267 354 270 357 
rect 267 357 270 360 
rect 267 360 270 363 
rect 267 363 270 366 
rect 267 366 270 369 
rect 267 369 270 372 
rect 267 372 270 375 
rect 267 375 270 378 
rect 267 378 270 381 
rect 267 381 270 384 
rect 267 384 270 387 
rect 267 387 270 390 
rect 267 390 270 393 
rect 267 393 270 396 
rect 267 396 270 399 
rect 267 399 270 402 
rect 267 402 270 405 
rect 267 405 270 408 
rect 267 408 270 411 
rect 267 411 270 414 
rect 267 414 270 417 
rect 267 417 270 420 
rect 267 420 270 423 
rect 267 423 270 426 
rect 267 426 270 429 
rect 267 429 270 432 
rect 267 432 270 435 
rect 267 435 270 438 
rect 267 438 270 441 
rect 267 441 270 444 
rect 267 444 270 447 
rect 267 447 270 450 
rect 267 450 270 453 
rect 267 453 270 456 
rect 267 456 270 459 
rect 267 459 270 462 
rect 267 462 270 465 
rect 267 465 270 468 
rect 267 468 270 471 
rect 267 471 270 474 
rect 267 474 270 477 
rect 267 477 270 480 
rect 267 480 270 483 
rect 267 483 270 486 
rect 267 486 270 489 
rect 267 489 270 492 
rect 267 492 270 495 
rect 267 495 270 498 
rect 267 498 270 501 
rect 267 501 270 504 
rect 267 504 270 507 
rect 267 507 270 510 
rect 270 0 273 3 
rect 270 3 273 6 
rect 270 6 273 9 
rect 270 9 273 12 
rect 270 12 273 15 
rect 270 15 273 18 
rect 270 18 273 21 
rect 270 21 273 24 
rect 270 24 273 27 
rect 270 27 273 30 
rect 270 30 273 33 
rect 270 33 273 36 
rect 270 36 273 39 
rect 270 39 273 42 
rect 270 42 273 45 
rect 270 45 273 48 
rect 270 48 273 51 
rect 270 51 273 54 
rect 270 54 273 57 
rect 270 57 273 60 
rect 270 60 273 63 
rect 270 63 273 66 
rect 270 66 273 69 
rect 270 69 273 72 
rect 270 72 273 75 
rect 270 75 273 78 
rect 270 78 273 81 
rect 270 81 273 84 
rect 270 84 273 87 
rect 270 87 273 90 
rect 270 90 273 93 
rect 270 93 273 96 
rect 270 96 273 99 
rect 270 99 273 102 
rect 270 102 273 105 
rect 270 105 273 108 
rect 270 108 273 111 
rect 270 111 273 114 
rect 270 114 273 117 
rect 270 117 273 120 
rect 270 120 273 123 
rect 270 123 273 126 
rect 270 126 273 129 
rect 270 129 273 132 
rect 270 132 273 135 
rect 270 135 273 138 
rect 270 138 273 141 
rect 270 141 273 144 
rect 270 144 273 147 
rect 270 147 273 150 
rect 270 150 273 153 
rect 270 153 273 156 
rect 270 156 273 159 
rect 270 159 273 162 
rect 270 162 273 165 
rect 270 165 273 168 
rect 270 168 273 171 
rect 270 171 273 174 
rect 270 174 273 177 
rect 270 177 273 180 
rect 270 180 273 183 
rect 270 183 273 186 
rect 270 186 273 189 
rect 270 189 273 192 
rect 270 192 273 195 
rect 270 195 273 198 
rect 270 198 273 201 
rect 270 201 273 204 
rect 270 204 273 207 
rect 270 207 273 210 
rect 270 210 273 213 
rect 270 213 273 216 
rect 270 216 273 219 
rect 270 219 273 222 
rect 270 222 273 225 
rect 270 225 273 228 
rect 270 228 273 231 
rect 270 231 273 234 
rect 270 234 273 237 
rect 270 237 273 240 
rect 270 240 273 243 
rect 270 243 273 246 
rect 270 246 273 249 
rect 270 249 273 252 
rect 270 252 273 255 
rect 270 255 273 258 
rect 270 258 273 261 
rect 270 261 273 264 
rect 270 264 273 267 
rect 270 267 273 270 
rect 270 270 273 273 
rect 270 273 273 276 
rect 270 276 273 279 
rect 270 279 273 282 
rect 270 282 273 285 
rect 270 285 273 288 
rect 270 288 273 291 
rect 270 291 273 294 
rect 270 294 273 297 
rect 270 297 273 300 
rect 270 300 273 303 
rect 270 303 273 306 
rect 270 306 273 309 
rect 270 309 273 312 
rect 270 312 273 315 
rect 270 315 273 318 
rect 270 318 273 321 
rect 270 321 273 324 
rect 270 324 273 327 
rect 270 327 273 330 
rect 270 330 273 333 
rect 270 333 273 336 
rect 270 336 273 339 
rect 270 339 273 342 
rect 270 342 273 345 
rect 270 345 273 348 
rect 270 348 273 351 
rect 270 351 273 354 
rect 270 354 273 357 
rect 270 357 273 360 
rect 270 360 273 363 
rect 270 363 273 366 
rect 270 366 273 369 
rect 270 369 273 372 
rect 270 372 273 375 
rect 270 375 273 378 
rect 270 378 273 381 
rect 270 381 273 384 
rect 270 384 273 387 
rect 270 387 273 390 
rect 270 390 273 393 
rect 270 393 273 396 
rect 270 396 273 399 
rect 270 399 273 402 
rect 270 402 273 405 
rect 270 405 273 408 
rect 270 408 273 411 
rect 270 411 273 414 
rect 270 414 273 417 
rect 270 417 273 420 
rect 270 420 273 423 
rect 270 423 273 426 
rect 270 426 273 429 
rect 270 429 273 432 
rect 270 432 273 435 
rect 270 435 273 438 
rect 270 438 273 441 
rect 270 441 273 444 
rect 270 444 273 447 
rect 270 447 273 450 
rect 270 450 273 453 
rect 270 453 273 456 
rect 270 456 273 459 
rect 270 459 273 462 
rect 270 462 273 465 
rect 270 465 273 468 
rect 270 468 273 471 
rect 270 471 273 474 
rect 270 474 273 477 
rect 270 477 273 480 
rect 270 480 273 483 
rect 270 483 273 486 
rect 270 486 273 489 
rect 270 489 273 492 
rect 270 492 273 495 
rect 270 495 273 498 
rect 270 498 273 501 
rect 270 501 273 504 
rect 270 504 273 507 
rect 270 507 273 510 
rect 273 0 276 3 
rect 273 3 276 6 
rect 273 6 276 9 
rect 273 9 276 12 
rect 273 12 276 15 
rect 273 15 276 18 
rect 273 18 276 21 
rect 273 21 276 24 
rect 273 24 276 27 
rect 273 27 276 30 
rect 273 30 276 33 
rect 273 33 276 36 
rect 273 36 276 39 
rect 273 39 276 42 
rect 273 42 276 45 
rect 273 45 276 48 
rect 273 48 276 51 
rect 273 51 276 54 
rect 273 54 276 57 
rect 273 57 276 60 
rect 273 60 276 63 
rect 273 63 276 66 
rect 273 66 276 69 
rect 273 69 276 72 
rect 273 72 276 75 
rect 273 75 276 78 
rect 273 78 276 81 
rect 273 81 276 84 
rect 273 84 276 87 
rect 273 87 276 90 
rect 273 90 276 93 
rect 273 93 276 96 
rect 273 96 276 99 
rect 273 99 276 102 
rect 273 102 276 105 
rect 273 105 276 108 
rect 273 108 276 111 
rect 273 111 276 114 
rect 273 114 276 117 
rect 273 117 276 120 
rect 273 120 276 123 
rect 273 123 276 126 
rect 273 126 276 129 
rect 273 129 276 132 
rect 273 132 276 135 
rect 273 135 276 138 
rect 273 138 276 141 
rect 273 141 276 144 
rect 273 144 276 147 
rect 273 147 276 150 
rect 273 150 276 153 
rect 273 153 276 156 
rect 273 156 276 159 
rect 273 159 276 162 
rect 273 162 276 165 
rect 273 165 276 168 
rect 273 168 276 171 
rect 273 171 276 174 
rect 273 174 276 177 
rect 273 177 276 180 
rect 273 180 276 183 
rect 273 183 276 186 
rect 273 186 276 189 
rect 273 189 276 192 
rect 273 192 276 195 
rect 273 195 276 198 
rect 273 198 276 201 
rect 273 201 276 204 
rect 273 204 276 207 
rect 273 207 276 210 
rect 273 210 276 213 
rect 273 213 276 216 
rect 273 216 276 219 
rect 273 219 276 222 
rect 273 222 276 225 
rect 273 225 276 228 
rect 273 228 276 231 
rect 273 231 276 234 
rect 273 234 276 237 
rect 273 237 276 240 
rect 273 240 276 243 
rect 273 243 276 246 
rect 273 246 276 249 
rect 273 249 276 252 
rect 273 252 276 255 
rect 273 255 276 258 
rect 273 258 276 261 
rect 273 261 276 264 
rect 273 264 276 267 
rect 273 267 276 270 
rect 273 270 276 273 
rect 273 273 276 276 
rect 273 276 276 279 
rect 273 279 276 282 
rect 273 282 276 285 
rect 273 285 276 288 
rect 273 288 276 291 
rect 273 291 276 294 
rect 273 294 276 297 
rect 273 297 276 300 
rect 273 300 276 303 
rect 273 303 276 306 
rect 273 306 276 309 
rect 273 309 276 312 
rect 273 312 276 315 
rect 273 315 276 318 
rect 273 318 276 321 
rect 273 321 276 324 
rect 273 324 276 327 
rect 273 327 276 330 
rect 273 330 276 333 
rect 273 333 276 336 
rect 273 336 276 339 
rect 273 339 276 342 
rect 273 342 276 345 
rect 273 345 276 348 
rect 273 348 276 351 
rect 273 351 276 354 
rect 273 354 276 357 
rect 273 357 276 360 
rect 273 360 276 363 
rect 273 363 276 366 
rect 273 366 276 369 
rect 273 369 276 372 
rect 273 372 276 375 
rect 273 375 276 378 
rect 273 378 276 381 
rect 273 381 276 384 
rect 273 384 276 387 
rect 273 387 276 390 
rect 273 390 276 393 
rect 273 393 276 396 
rect 273 396 276 399 
rect 273 399 276 402 
rect 273 402 276 405 
rect 273 405 276 408 
rect 273 408 276 411 
rect 273 411 276 414 
rect 273 414 276 417 
rect 273 417 276 420 
rect 273 420 276 423 
rect 273 423 276 426 
rect 273 426 276 429 
rect 273 429 276 432 
rect 273 432 276 435 
rect 273 435 276 438 
rect 273 438 276 441 
rect 273 441 276 444 
rect 273 444 276 447 
rect 273 447 276 450 
rect 273 450 276 453 
rect 273 453 276 456 
rect 273 456 276 459 
rect 273 459 276 462 
rect 273 462 276 465 
rect 273 465 276 468 
rect 273 468 276 471 
rect 273 471 276 474 
rect 273 474 276 477 
rect 273 477 276 480 
rect 273 480 276 483 
rect 273 483 276 486 
rect 273 486 276 489 
rect 273 489 276 492 
rect 273 492 276 495 
rect 273 495 276 498 
rect 273 498 276 501 
rect 273 501 276 504 
rect 273 504 276 507 
rect 273 507 276 510 
rect 276 0 279 3 
rect 276 3 279 6 
rect 276 6 279 9 
rect 276 9 279 12 
rect 276 12 279 15 
rect 276 15 279 18 
rect 276 18 279 21 
rect 276 21 279 24 
rect 276 24 279 27 
rect 276 27 279 30 
rect 276 30 279 33 
rect 276 33 279 36 
rect 276 36 279 39 
rect 276 39 279 42 
rect 276 42 279 45 
rect 276 45 279 48 
rect 276 48 279 51 
rect 276 51 279 54 
rect 276 54 279 57 
rect 276 57 279 60 
rect 276 60 279 63 
rect 276 63 279 66 
rect 276 66 279 69 
rect 276 69 279 72 
rect 276 72 279 75 
rect 276 75 279 78 
rect 276 78 279 81 
rect 276 81 279 84 
rect 276 84 279 87 
rect 276 87 279 90 
rect 276 90 279 93 
rect 276 93 279 96 
rect 276 96 279 99 
rect 276 99 279 102 
rect 276 102 279 105 
rect 276 105 279 108 
rect 276 108 279 111 
rect 276 111 279 114 
rect 276 114 279 117 
rect 276 117 279 120 
rect 276 120 279 123 
rect 276 123 279 126 
rect 276 126 279 129 
rect 276 129 279 132 
rect 276 132 279 135 
rect 276 135 279 138 
rect 276 138 279 141 
rect 276 141 279 144 
rect 276 144 279 147 
rect 276 147 279 150 
rect 276 150 279 153 
rect 276 153 279 156 
rect 276 156 279 159 
rect 276 159 279 162 
rect 276 162 279 165 
rect 276 165 279 168 
rect 276 168 279 171 
rect 276 171 279 174 
rect 276 174 279 177 
rect 276 177 279 180 
rect 276 180 279 183 
rect 276 183 279 186 
rect 276 186 279 189 
rect 276 189 279 192 
rect 276 192 279 195 
rect 276 195 279 198 
rect 276 198 279 201 
rect 276 201 279 204 
rect 276 204 279 207 
rect 276 207 279 210 
rect 276 210 279 213 
rect 276 213 279 216 
rect 276 216 279 219 
rect 276 219 279 222 
rect 276 222 279 225 
rect 276 225 279 228 
rect 276 228 279 231 
rect 276 231 279 234 
rect 276 234 279 237 
rect 276 237 279 240 
rect 276 240 279 243 
rect 276 243 279 246 
rect 276 246 279 249 
rect 276 249 279 252 
rect 276 252 279 255 
rect 276 255 279 258 
rect 276 258 279 261 
rect 276 261 279 264 
rect 276 264 279 267 
rect 276 267 279 270 
rect 276 270 279 273 
rect 276 273 279 276 
rect 276 276 279 279 
rect 276 279 279 282 
rect 276 282 279 285 
rect 276 285 279 288 
rect 276 288 279 291 
rect 276 291 279 294 
rect 276 294 279 297 
rect 276 297 279 300 
rect 276 300 279 303 
rect 276 303 279 306 
rect 276 306 279 309 
rect 276 309 279 312 
rect 276 312 279 315 
rect 276 315 279 318 
rect 276 318 279 321 
rect 276 321 279 324 
rect 276 324 279 327 
rect 276 327 279 330 
rect 276 330 279 333 
rect 276 333 279 336 
rect 276 336 279 339 
rect 276 339 279 342 
rect 276 342 279 345 
rect 276 345 279 348 
rect 276 348 279 351 
rect 276 351 279 354 
rect 276 354 279 357 
rect 276 357 279 360 
rect 276 360 279 363 
rect 276 363 279 366 
rect 276 366 279 369 
rect 276 369 279 372 
rect 276 372 279 375 
rect 276 375 279 378 
rect 276 378 279 381 
rect 276 381 279 384 
rect 276 384 279 387 
rect 276 387 279 390 
rect 276 390 279 393 
rect 276 393 279 396 
rect 276 396 279 399 
rect 276 399 279 402 
rect 276 402 279 405 
rect 276 405 279 408 
rect 276 408 279 411 
rect 276 411 279 414 
rect 276 414 279 417 
rect 276 417 279 420 
rect 276 420 279 423 
rect 276 423 279 426 
rect 276 426 279 429 
rect 276 429 279 432 
rect 276 432 279 435 
rect 276 435 279 438 
rect 276 438 279 441 
rect 276 441 279 444 
rect 276 444 279 447 
rect 276 447 279 450 
rect 276 450 279 453 
rect 276 453 279 456 
rect 276 456 279 459 
rect 276 459 279 462 
rect 276 462 279 465 
rect 276 465 279 468 
rect 276 468 279 471 
rect 276 471 279 474 
rect 276 474 279 477 
rect 276 477 279 480 
rect 276 480 279 483 
rect 276 483 279 486 
rect 276 486 279 489 
rect 276 489 279 492 
rect 276 492 279 495 
rect 276 495 279 498 
rect 276 498 279 501 
rect 276 501 279 504 
rect 276 504 279 507 
rect 276 507 279 510 
rect 279 0 282 3 
rect 279 3 282 6 
rect 279 6 282 9 
rect 279 9 282 12 
rect 279 12 282 15 
rect 279 15 282 18 
rect 279 18 282 21 
rect 279 21 282 24 
rect 279 24 282 27 
rect 279 27 282 30 
rect 279 30 282 33 
rect 279 33 282 36 
rect 279 36 282 39 
rect 279 39 282 42 
rect 279 42 282 45 
rect 279 45 282 48 
rect 279 48 282 51 
rect 279 51 282 54 
rect 279 54 282 57 
rect 279 57 282 60 
rect 279 60 282 63 
rect 279 63 282 66 
rect 279 66 282 69 
rect 279 69 282 72 
rect 279 72 282 75 
rect 279 75 282 78 
rect 279 78 282 81 
rect 279 81 282 84 
rect 279 84 282 87 
rect 279 87 282 90 
rect 279 90 282 93 
rect 279 93 282 96 
rect 279 96 282 99 
rect 279 99 282 102 
rect 279 102 282 105 
rect 279 105 282 108 
rect 279 108 282 111 
rect 279 111 282 114 
rect 279 114 282 117 
rect 279 117 282 120 
rect 279 120 282 123 
rect 279 123 282 126 
rect 279 126 282 129 
rect 279 129 282 132 
rect 279 132 282 135 
rect 279 135 282 138 
rect 279 138 282 141 
rect 279 141 282 144 
rect 279 144 282 147 
rect 279 147 282 150 
rect 279 150 282 153 
rect 279 153 282 156 
rect 279 156 282 159 
rect 279 159 282 162 
rect 279 162 282 165 
rect 279 165 282 168 
rect 279 168 282 171 
rect 279 171 282 174 
rect 279 174 282 177 
rect 279 177 282 180 
rect 279 180 282 183 
rect 279 183 282 186 
rect 279 186 282 189 
rect 279 189 282 192 
rect 279 192 282 195 
rect 279 195 282 198 
rect 279 198 282 201 
rect 279 201 282 204 
rect 279 204 282 207 
rect 279 207 282 210 
rect 279 210 282 213 
rect 279 213 282 216 
rect 279 216 282 219 
rect 279 219 282 222 
rect 279 222 282 225 
rect 279 225 282 228 
rect 279 228 282 231 
rect 279 231 282 234 
rect 279 234 282 237 
rect 279 237 282 240 
rect 279 240 282 243 
rect 279 243 282 246 
rect 279 246 282 249 
rect 279 249 282 252 
rect 279 252 282 255 
rect 279 255 282 258 
rect 279 258 282 261 
rect 279 261 282 264 
rect 279 264 282 267 
rect 279 267 282 270 
rect 279 270 282 273 
rect 279 273 282 276 
rect 279 276 282 279 
rect 279 279 282 282 
rect 279 282 282 285 
rect 279 285 282 288 
rect 279 288 282 291 
rect 279 291 282 294 
rect 279 294 282 297 
rect 279 297 282 300 
rect 279 300 282 303 
rect 279 303 282 306 
rect 279 306 282 309 
rect 279 309 282 312 
rect 279 312 282 315 
rect 279 315 282 318 
rect 279 318 282 321 
rect 279 321 282 324 
rect 279 324 282 327 
rect 279 327 282 330 
rect 279 330 282 333 
rect 279 333 282 336 
rect 279 336 282 339 
rect 279 339 282 342 
rect 279 342 282 345 
rect 279 345 282 348 
rect 279 348 282 351 
rect 279 351 282 354 
rect 279 354 282 357 
rect 279 357 282 360 
rect 279 360 282 363 
rect 279 363 282 366 
rect 279 366 282 369 
rect 279 369 282 372 
rect 279 372 282 375 
rect 279 375 282 378 
rect 279 378 282 381 
rect 279 381 282 384 
rect 279 384 282 387 
rect 279 387 282 390 
rect 279 390 282 393 
rect 279 393 282 396 
rect 279 396 282 399 
rect 279 399 282 402 
rect 279 402 282 405 
rect 279 405 282 408 
rect 279 408 282 411 
rect 279 411 282 414 
rect 279 414 282 417 
rect 279 417 282 420 
rect 279 420 282 423 
rect 279 423 282 426 
rect 279 426 282 429 
rect 279 429 282 432 
rect 279 432 282 435 
rect 279 435 282 438 
rect 279 438 282 441 
rect 279 441 282 444 
rect 279 444 282 447 
rect 279 447 282 450 
rect 279 450 282 453 
rect 279 453 282 456 
rect 279 456 282 459 
rect 279 459 282 462 
rect 279 462 282 465 
rect 279 465 282 468 
rect 279 468 282 471 
rect 279 471 282 474 
rect 279 474 282 477 
rect 279 477 282 480 
rect 279 480 282 483 
rect 279 483 282 486 
rect 279 486 282 489 
rect 279 489 282 492 
rect 279 492 282 495 
rect 279 495 282 498 
rect 279 498 282 501 
rect 279 501 282 504 
rect 279 504 282 507 
rect 279 507 282 510 
rect 282 0 285 3 
rect 282 3 285 6 
rect 282 6 285 9 
rect 282 9 285 12 
rect 282 12 285 15 
rect 282 15 285 18 
rect 282 18 285 21 
rect 282 21 285 24 
rect 282 24 285 27 
rect 282 27 285 30 
rect 282 30 285 33 
rect 282 33 285 36 
rect 282 36 285 39 
rect 282 39 285 42 
rect 282 42 285 45 
rect 282 45 285 48 
rect 282 48 285 51 
rect 282 51 285 54 
rect 282 54 285 57 
rect 282 57 285 60 
rect 282 60 285 63 
rect 282 63 285 66 
rect 282 66 285 69 
rect 282 69 285 72 
rect 282 72 285 75 
rect 282 75 285 78 
rect 282 78 285 81 
rect 282 81 285 84 
rect 282 84 285 87 
rect 282 87 285 90 
rect 282 90 285 93 
rect 282 93 285 96 
rect 282 96 285 99 
rect 282 99 285 102 
rect 282 102 285 105 
rect 282 105 285 108 
rect 282 108 285 111 
rect 282 111 285 114 
rect 282 114 285 117 
rect 282 117 285 120 
rect 282 120 285 123 
rect 282 123 285 126 
rect 282 126 285 129 
rect 282 129 285 132 
rect 282 132 285 135 
rect 282 135 285 138 
rect 282 138 285 141 
rect 282 141 285 144 
rect 282 144 285 147 
rect 282 147 285 150 
rect 282 150 285 153 
rect 282 153 285 156 
rect 282 156 285 159 
rect 282 159 285 162 
rect 282 162 285 165 
rect 282 165 285 168 
rect 282 168 285 171 
rect 282 171 285 174 
rect 282 174 285 177 
rect 282 177 285 180 
rect 282 180 285 183 
rect 282 183 285 186 
rect 282 186 285 189 
rect 282 189 285 192 
rect 282 192 285 195 
rect 282 195 285 198 
rect 282 198 285 201 
rect 282 201 285 204 
rect 282 204 285 207 
rect 282 207 285 210 
rect 282 210 285 213 
rect 282 213 285 216 
rect 282 216 285 219 
rect 282 219 285 222 
rect 282 222 285 225 
rect 282 225 285 228 
rect 282 228 285 231 
rect 282 231 285 234 
rect 282 234 285 237 
rect 282 237 285 240 
rect 282 240 285 243 
rect 282 243 285 246 
rect 282 246 285 249 
rect 282 249 285 252 
rect 282 252 285 255 
rect 282 255 285 258 
rect 282 258 285 261 
rect 282 261 285 264 
rect 282 264 285 267 
rect 282 267 285 270 
rect 282 270 285 273 
rect 282 273 285 276 
rect 282 276 285 279 
rect 282 279 285 282 
rect 282 282 285 285 
rect 282 285 285 288 
rect 282 288 285 291 
rect 282 291 285 294 
rect 282 294 285 297 
rect 282 297 285 300 
rect 282 300 285 303 
rect 282 303 285 306 
rect 282 306 285 309 
rect 282 309 285 312 
rect 282 312 285 315 
rect 282 315 285 318 
rect 282 318 285 321 
rect 282 321 285 324 
rect 282 324 285 327 
rect 282 327 285 330 
rect 282 330 285 333 
rect 282 333 285 336 
rect 282 336 285 339 
rect 282 339 285 342 
rect 282 342 285 345 
rect 282 345 285 348 
rect 282 348 285 351 
rect 282 351 285 354 
rect 282 354 285 357 
rect 282 357 285 360 
rect 282 360 285 363 
rect 282 363 285 366 
rect 282 366 285 369 
rect 282 369 285 372 
rect 282 372 285 375 
rect 282 375 285 378 
rect 282 378 285 381 
rect 282 381 285 384 
rect 282 384 285 387 
rect 282 387 285 390 
rect 282 390 285 393 
rect 282 393 285 396 
rect 282 396 285 399 
rect 282 399 285 402 
rect 282 402 285 405 
rect 282 405 285 408 
rect 282 408 285 411 
rect 282 411 285 414 
rect 282 414 285 417 
rect 282 417 285 420 
rect 282 420 285 423 
rect 282 423 285 426 
rect 282 426 285 429 
rect 282 429 285 432 
rect 282 432 285 435 
rect 282 435 285 438 
rect 282 438 285 441 
rect 282 441 285 444 
rect 282 444 285 447 
rect 282 447 285 450 
rect 282 450 285 453 
rect 282 453 285 456 
rect 282 456 285 459 
rect 282 459 285 462 
rect 282 462 285 465 
rect 282 465 285 468 
rect 282 468 285 471 
rect 282 471 285 474 
rect 282 474 285 477 
rect 282 477 285 480 
rect 282 480 285 483 
rect 282 483 285 486 
rect 282 486 285 489 
rect 282 489 285 492 
rect 282 492 285 495 
rect 282 495 285 498 
rect 282 498 285 501 
rect 282 501 285 504 
rect 282 504 285 507 
rect 282 507 285 510 
rect 285 0 288 3 
rect 285 3 288 6 
rect 285 6 288 9 
rect 285 9 288 12 
rect 285 12 288 15 
rect 285 15 288 18 
rect 285 18 288 21 
rect 285 21 288 24 
rect 285 24 288 27 
rect 285 27 288 30 
rect 285 30 288 33 
rect 285 33 288 36 
rect 285 36 288 39 
rect 285 39 288 42 
rect 285 42 288 45 
rect 285 45 288 48 
rect 285 48 288 51 
rect 285 51 288 54 
rect 285 54 288 57 
rect 285 57 288 60 
rect 285 60 288 63 
rect 285 63 288 66 
rect 285 66 288 69 
rect 285 69 288 72 
rect 285 72 288 75 
rect 285 75 288 78 
rect 285 78 288 81 
rect 285 81 288 84 
rect 285 84 288 87 
rect 285 87 288 90 
rect 285 90 288 93 
rect 285 93 288 96 
rect 285 96 288 99 
rect 285 99 288 102 
rect 285 102 288 105 
rect 285 105 288 108 
rect 285 108 288 111 
rect 285 111 288 114 
rect 285 114 288 117 
rect 285 117 288 120 
rect 285 120 288 123 
rect 285 123 288 126 
rect 285 126 288 129 
rect 285 129 288 132 
rect 285 132 288 135 
rect 285 135 288 138 
rect 285 138 288 141 
rect 285 141 288 144 
rect 285 144 288 147 
rect 285 147 288 150 
rect 285 150 288 153 
rect 285 153 288 156 
rect 285 156 288 159 
rect 285 159 288 162 
rect 285 162 288 165 
rect 285 165 288 168 
rect 285 168 288 171 
rect 285 171 288 174 
rect 285 174 288 177 
rect 285 177 288 180 
rect 285 180 288 183 
rect 285 183 288 186 
rect 285 186 288 189 
rect 285 189 288 192 
rect 285 192 288 195 
rect 285 195 288 198 
rect 285 198 288 201 
rect 285 201 288 204 
rect 285 204 288 207 
rect 285 207 288 210 
rect 285 210 288 213 
rect 285 213 288 216 
rect 285 216 288 219 
rect 285 219 288 222 
rect 285 222 288 225 
rect 285 225 288 228 
rect 285 228 288 231 
rect 285 231 288 234 
rect 285 234 288 237 
rect 285 237 288 240 
rect 285 240 288 243 
rect 285 243 288 246 
rect 285 246 288 249 
rect 285 249 288 252 
rect 285 252 288 255 
rect 285 255 288 258 
rect 285 258 288 261 
rect 285 261 288 264 
rect 285 264 288 267 
rect 285 267 288 270 
rect 285 270 288 273 
rect 285 273 288 276 
rect 285 276 288 279 
rect 285 279 288 282 
rect 285 282 288 285 
rect 285 285 288 288 
rect 285 288 288 291 
rect 285 291 288 294 
rect 285 294 288 297 
rect 285 297 288 300 
rect 285 300 288 303 
rect 285 303 288 306 
rect 285 306 288 309 
rect 285 309 288 312 
rect 285 312 288 315 
rect 285 315 288 318 
rect 285 318 288 321 
rect 285 321 288 324 
rect 285 324 288 327 
rect 285 327 288 330 
rect 285 330 288 333 
rect 285 333 288 336 
rect 285 336 288 339 
rect 285 339 288 342 
rect 285 342 288 345 
rect 285 345 288 348 
rect 285 348 288 351 
rect 285 351 288 354 
rect 285 354 288 357 
rect 285 357 288 360 
rect 285 360 288 363 
rect 285 363 288 366 
rect 285 366 288 369 
rect 285 369 288 372 
rect 285 372 288 375 
rect 285 375 288 378 
rect 285 378 288 381 
rect 285 381 288 384 
rect 285 384 288 387 
rect 285 387 288 390 
rect 285 390 288 393 
rect 285 393 288 396 
rect 285 396 288 399 
rect 285 399 288 402 
rect 285 402 288 405 
rect 285 405 288 408 
rect 285 408 288 411 
rect 285 411 288 414 
rect 285 414 288 417 
rect 285 417 288 420 
rect 285 420 288 423 
rect 285 423 288 426 
rect 285 426 288 429 
rect 285 429 288 432 
rect 285 432 288 435 
rect 285 435 288 438 
rect 285 438 288 441 
rect 285 441 288 444 
rect 285 444 288 447 
rect 285 447 288 450 
rect 285 450 288 453 
rect 285 453 288 456 
rect 285 456 288 459 
rect 285 459 288 462 
rect 285 462 288 465 
rect 285 465 288 468 
rect 285 468 288 471 
rect 285 471 288 474 
rect 285 474 288 477 
rect 285 477 288 480 
rect 285 480 288 483 
rect 285 483 288 486 
rect 285 486 288 489 
rect 285 489 288 492 
rect 285 492 288 495 
rect 285 495 288 498 
rect 285 498 288 501 
rect 285 501 288 504 
rect 285 504 288 507 
rect 285 507 288 510 
rect 288 0 291 3 
rect 288 3 291 6 
rect 288 6 291 9 
rect 288 9 291 12 
rect 288 12 291 15 
rect 288 15 291 18 
rect 288 18 291 21 
rect 288 21 291 24 
rect 288 24 291 27 
rect 288 27 291 30 
rect 288 30 291 33 
rect 288 33 291 36 
rect 288 36 291 39 
rect 288 39 291 42 
rect 288 42 291 45 
rect 288 45 291 48 
rect 288 48 291 51 
rect 288 51 291 54 
rect 288 54 291 57 
rect 288 57 291 60 
rect 288 60 291 63 
rect 288 63 291 66 
rect 288 66 291 69 
rect 288 69 291 72 
rect 288 72 291 75 
rect 288 75 291 78 
rect 288 78 291 81 
rect 288 81 291 84 
rect 288 84 291 87 
rect 288 87 291 90 
rect 288 90 291 93 
rect 288 93 291 96 
rect 288 96 291 99 
rect 288 99 291 102 
rect 288 102 291 105 
rect 288 105 291 108 
rect 288 108 291 111 
rect 288 111 291 114 
rect 288 114 291 117 
rect 288 117 291 120 
rect 288 120 291 123 
rect 288 123 291 126 
rect 288 126 291 129 
rect 288 129 291 132 
rect 288 132 291 135 
rect 288 135 291 138 
rect 288 138 291 141 
rect 288 141 291 144 
rect 288 144 291 147 
rect 288 147 291 150 
rect 288 150 291 153 
rect 288 153 291 156 
rect 288 156 291 159 
rect 288 159 291 162 
rect 288 162 291 165 
rect 288 165 291 168 
rect 288 168 291 171 
rect 288 171 291 174 
rect 288 174 291 177 
rect 288 177 291 180 
rect 288 180 291 183 
rect 288 183 291 186 
rect 288 186 291 189 
rect 288 189 291 192 
rect 288 192 291 195 
rect 288 195 291 198 
rect 288 198 291 201 
rect 288 201 291 204 
rect 288 204 291 207 
rect 288 207 291 210 
rect 288 210 291 213 
rect 288 213 291 216 
rect 288 216 291 219 
rect 288 219 291 222 
rect 288 222 291 225 
rect 288 225 291 228 
rect 288 228 291 231 
rect 288 231 291 234 
rect 288 234 291 237 
rect 288 237 291 240 
rect 288 240 291 243 
rect 288 243 291 246 
rect 288 246 291 249 
rect 288 249 291 252 
rect 288 252 291 255 
rect 288 255 291 258 
rect 288 258 291 261 
rect 288 261 291 264 
rect 288 264 291 267 
rect 288 267 291 270 
rect 288 270 291 273 
rect 288 273 291 276 
rect 288 276 291 279 
rect 288 279 291 282 
rect 288 282 291 285 
rect 288 285 291 288 
rect 288 288 291 291 
rect 288 291 291 294 
rect 288 294 291 297 
rect 288 297 291 300 
rect 288 300 291 303 
rect 288 303 291 306 
rect 288 306 291 309 
rect 288 309 291 312 
rect 288 312 291 315 
rect 288 315 291 318 
rect 288 318 291 321 
rect 288 321 291 324 
rect 288 324 291 327 
rect 288 327 291 330 
rect 288 330 291 333 
rect 288 333 291 336 
rect 288 336 291 339 
rect 288 339 291 342 
rect 288 342 291 345 
rect 288 345 291 348 
rect 288 348 291 351 
rect 288 351 291 354 
rect 288 354 291 357 
rect 288 357 291 360 
rect 288 360 291 363 
rect 288 363 291 366 
rect 288 366 291 369 
rect 288 369 291 372 
rect 288 372 291 375 
rect 288 375 291 378 
rect 288 378 291 381 
rect 288 381 291 384 
rect 288 384 291 387 
rect 288 387 291 390 
rect 288 390 291 393 
rect 288 393 291 396 
rect 288 396 291 399 
rect 288 399 291 402 
rect 288 402 291 405 
rect 288 405 291 408 
rect 288 408 291 411 
rect 288 411 291 414 
rect 288 414 291 417 
rect 288 417 291 420 
rect 288 420 291 423 
rect 288 423 291 426 
rect 288 426 291 429 
rect 288 429 291 432 
rect 288 432 291 435 
rect 288 435 291 438 
rect 288 438 291 441 
rect 288 441 291 444 
rect 288 444 291 447 
rect 288 447 291 450 
rect 288 450 291 453 
rect 288 453 291 456 
rect 288 456 291 459 
rect 288 459 291 462 
rect 288 462 291 465 
rect 288 465 291 468 
rect 288 468 291 471 
rect 288 471 291 474 
rect 288 474 291 477 
rect 288 477 291 480 
rect 288 480 291 483 
rect 288 483 291 486 
rect 288 486 291 489 
rect 288 489 291 492 
rect 288 492 291 495 
rect 288 495 291 498 
rect 288 498 291 501 
rect 288 501 291 504 
rect 288 504 291 507 
rect 288 507 291 510 
rect 291 0 294 3 
rect 291 3 294 6 
rect 291 6 294 9 
rect 291 9 294 12 
rect 291 12 294 15 
rect 291 15 294 18 
rect 291 18 294 21 
rect 291 21 294 24 
rect 291 24 294 27 
rect 291 27 294 30 
rect 291 30 294 33 
rect 291 33 294 36 
rect 291 36 294 39 
rect 291 39 294 42 
rect 291 42 294 45 
rect 291 45 294 48 
rect 291 48 294 51 
rect 291 51 294 54 
rect 291 54 294 57 
rect 291 57 294 60 
rect 291 60 294 63 
rect 291 63 294 66 
rect 291 66 294 69 
rect 291 69 294 72 
rect 291 72 294 75 
rect 291 75 294 78 
rect 291 78 294 81 
rect 291 81 294 84 
rect 291 84 294 87 
rect 291 87 294 90 
rect 291 90 294 93 
rect 291 93 294 96 
rect 291 96 294 99 
rect 291 99 294 102 
rect 291 102 294 105 
rect 291 105 294 108 
rect 291 108 294 111 
rect 291 111 294 114 
rect 291 114 294 117 
rect 291 117 294 120 
rect 291 120 294 123 
rect 291 123 294 126 
rect 291 126 294 129 
rect 291 129 294 132 
rect 291 132 294 135 
rect 291 135 294 138 
rect 291 138 294 141 
rect 291 141 294 144 
rect 291 144 294 147 
rect 291 147 294 150 
rect 291 150 294 153 
rect 291 153 294 156 
rect 291 156 294 159 
rect 291 159 294 162 
rect 291 162 294 165 
rect 291 165 294 168 
rect 291 168 294 171 
rect 291 171 294 174 
rect 291 174 294 177 
rect 291 177 294 180 
rect 291 180 294 183 
rect 291 183 294 186 
rect 291 186 294 189 
rect 291 189 294 192 
rect 291 192 294 195 
rect 291 195 294 198 
rect 291 198 294 201 
rect 291 201 294 204 
rect 291 204 294 207 
rect 291 207 294 210 
rect 291 210 294 213 
rect 291 213 294 216 
rect 291 216 294 219 
rect 291 219 294 222 
rect 291 222 294 225 
rect 291 225 294 228 
rect 291 228 294 231 
rect 291 231 294 234 
rect 291 234 294 237 
rect 291 237 294 240 
rect 291 240 294 243 
rect 291 243 294 246 
rect 291 246 294 249 
rect 291 249 294 252 
rect 291 252 294 255 
rect 291 255 294 258 
rect 291 258 294 261 
rect 291 261 294 264 
rect 291 264 294 267 
rect 291 267 294 270 
rect 291 270 294 273 
rect 291 273 294 276 
rect 291 276 294 279 
rect 291 279 294 282 
rect 291 282 294 285 
rect 291 285 294 288 
rect 291 288 294 291 
rect 291 291 294 294 
rect 291 294 294 297 
rect 291 297 294 300 
rect 291 300 294 303 
rect 291 303 294 306 
rect 291 306 294 309 
rect 291 309 294 312 
rect 291 312 294 315 
rect 291 315 294 318 
rect 291 318 294 321 
rect 291 321 294 324 
rect 291 324 294 327 
rect 291 327 294 330 
rect 291 330 294 333 
rect 291 333 294 336 
rect 291 336 294 339 
rect 291 339 294 342 
rect 291 342 294 345 
rect 291 345 294 348 
rect 291 348 294 351 
rect 291 351 294 354 
rect 291 354 294 357 
rect 291 357 294 360 
rect 291 360 294 363 
rect 291 363 294 366 
rect 291 366 294 369 
rect 291 369 294 372 
rect 291 372 294 375 
rect 291 375 294 378 
rect 291 378 294 381 
rect 291 381 294 384 
rect 291 384 294 387 
rect 291 387 294 390 
rect 291 390 294 393 
rect 291 393 294 396 
rect 291 396 294 399 
rect 291 399 294 402 
rect 291 402 294 405 
rect 291 405 294 408 
rect 291 408 294 411 
rect 291 411 294 414 
rect 291 414 294 417 
rect 291 417 294 420 
rect 291 420 294 423 
rect 291 423 294 426 
rect 291 426 294 429 
rect 291 429 294 432 
rect 291 432 294 435 
rect 291 435 294 438 
rect 291 438 294 441 
rect 291 441 294 444 
rect 291 444 294 447 
rect 291 447 294 450 
rect 291 450 294 453 
rect 291 453 294 456 
rect 291 456 294 459 
rect 291 459 294 462 
rect 291 462 294 465 
rect 291 465 294 468 
rect 291 468 294 471 
rect 291 471 294 474 
rect 291 474 294 477 
rect 291 477 294 480 
rect 291 480 294 483 
rect 291 483 294 486 
rect 291 486 294 489 
rect 291 489 294 492 
rect 291 492 294 495 
rect 291 495 294 498 
rect 291 498 294 501 
rect 291 501 294 504 
rect 291 504 294 507 
rect 291 507 294 510 
rect 294 0 297 3 
rect 294 3 297 6 
rect 294 6 297 9 
rect 294 9 297 12 
rect 294 12 297 15 
rect 294 15 297 18 
rect 294 18 297 21 
rect 294 21 297 24 
rect 294 24 297 27 
rect 294 27 297 30 
rect 294 30 297 33 
rect 294 33 297 36 
rect 294 36 297 39 
rect 294 39 297 42 
rect 294 42 297 45 
rect 294 45 297 48 
rect 294 48 297 51 
rect 294 51 297 54 
rect 294 54 297 57 
rect 294 57 297 60 
rect 294 60 297 63 
rect 294 63 297 66 
rect 294 66 297 69 
rect 294 69 297 72 
rect 294 72 297 75 
rect 294 75 297 78 
rect 294 78 297 81 
rect 294 81 297 84 
rect 294 84 297 87 
rect 294 87 297 90 
rect 294 90 297 93 
rect 294 93 297 96 
rect 294 96 297 99 
rect 294 99 297 102 
rect 294 102 297 105 
rect 294 105 297 108 
rect 294 108 297 111 
rect 294 111 297 114 
rect 294 114 297 117 
rect 294 117 297 120 
rect 294 120 297 123 
rect 294 123 297 126 
rect 294 126 297 129 
rect 294 129 297 132 
rect 294 132 297 135 
rect 294 135 297 138 
rect 294 138 297 141 
rect 294 141 297 144 
rect 294 144 297 147 
rect 294 147 297 150 
rect 294 150 297 153 
rect 294 153 297 156 
rect 294 156 297 159 
rect 294 159 297 162 
rect 294 162 297 165 
rect 294 165 297 168 
rect 294 168 297 171 
rect 294 171 297 174 
rect 294 174 297 177 
rect 294 177 297 180 
rect 294 180 297 183 
rect 294 183 297 186 
rect 294 186 297 189 
rect 294 189 297 192 
rect 294 192 297 195 
rect 294 195 297 198 
rect 294 198 297 201 
rect 294 201 297 204 
rect 294 204 297 207 
rect 294 207 297 210 
rect 294 210 297 213 
rect 294 213 297 216 
rect 294 216 297 219 
rect 294 219 297 222 
rect 294 222 297 225 
rect 294 225 297 228 
rect 294 228 297 231 
rect 294 231 297 234 
rect 294 234 297 237 
rect 294 237 297 240 
rect 294 240 297 243 
rect 294 243 297 246 
rect 294 246 297 249 
rect 294 249 297 252 
rect 294 252 297 255 
rect 294 255 297 258 
rect 294 258 297 261 
rect 294 261 297 264 
rect 294 264 297 267 
rect 294 267 297 270 
rect 294 270 297 273 
rect 294 273 297 276 
rect 294 276 297 279 
rect 294 279 297 282 
rect 294 282 297 285 
rect 294 285 297 288 
rect 294 288 297 291 
rect 294 291 297 294 
rect 294 294 297 297 
rect 294 297 297 300 
rect 294 300 297 303 
rect 294 303 297 306 
rect 294 306 297 309 
rect 294 309 297 312 
rect 294 312 297 315 
rect 294 315 297 318 
rect 294 318 297 321 
rect 294 321 297 324 
rect 294 324 297 327 
rect 294 327 297 330 
rect 294 330 297 333 
rect 294 333 297 336 
rect 294 336 297 339 
rect 294 339 297 342 
rect 294 342 297 345 
rect 294 345 297 348 
rect 294 348 297 351 
rect 294 351 297 354 
rect 294 354 297 357 
rect 294 357 297 360 
rect 294 360 297 363 
rect 294 363 297 366 
rect 294 366 297 369 
rect 294 369 297 372 
rect 294 372 297 375 
rect 294 375 297 378 
rect 294 378 297 381 
rect 294 381 297 384 
rect 294 384 297 387 
rect 294 387 297 390 
rect 294 390 297 393 
rect 294 393 297 396 
rect 294 396 297 399 
rect 294 399 297 402 
rect 294 402 297 405 
rect 294 405 297 408 
rect 294 408 297 411 
rect 294 411 297 414 
rect 294 414 297 417 
rect 294 417 297 420 
rect 294 420 297 423 
rect 294 423 297 426 
rect 294 426 297 429 
rect 294 429 297 432 
rect 294 432 297 435 
rect 294 435 297 438 
rect 294 438 297 441 
rect 294 441 297 444 
rect 294 444 297 447 
rect 294 447 297 450 
rect 294 450 297 453 
rect 294 453 297 456 
rect 294 456 297 459 
rect 294 459 297 462 
rect 294 462 297 465 
rect 294 465 297 468 
rect 294 468 297 471 
rect 294 471 297 474 
rect 294 474 297 477 
rect 294 477 297 480 
rect 294 480 297 483 
rect 294 483 297 486 
rect 294 486 297 489 
rect 294 489 297 492 
rect 294 492 297 495 
rect 294 495 297 498 
rect 294 498 297 501 
rect 294 501 297 504 
rect 294 504 297 507 
rect 294 507 297 510 
rect 297 0 300 3 
rect 297 3 300 6 
rect 297 6 300 9 
rect 297 9 300 12 
rect 297 12 300 15 
rect 297 15 300 18 
rect 297 18 300 21 
rect 297 21 300 24 
rect 297 24 300 27 
rect 297 27 300 30 
rect 297 30 300 33 
rect 297 33 300 36 
rect 297 36 300 39 
rect 297 39 300 42 
rect 297 42 300 45 
rect 297 45 300 48 
rect 297 48 300 51 
rect 297 51 300 54 
rect 297 54 300 57 
rect 297 57 300 60 
rect 297 60 300 63 
rect 297 63 300 66 
rect 297 66 300 69 
rect 297 69 300 72 
rect 297 72 300 75 
rect 297 75 300 78 
rect 297 78 300 81 
rect 297 81 300 84 
rect 297 84 300 87 
rect 297 87 300 90 
rect 297 90 300 93 
rect 297 93 300 96 
rect 297 96 300 99 
rect 297 99 300 102 
rect 297 102 300 105 
rect 297 105 300 108 
rect 297 108 300 111 
rect 297 111 300 114 
rect 297 114 300 117 
rect 297 117 300 120 
rect 297 120 300 123 
rect 297 123 300 126 
rect 297 126 300 129 
rect 297 129 300 132 
rect 297 132 300 135 
rect 297 135 300 138 
rect 297 138 300 141 
rect 297 141 300 144 
rect 297 144 300 147 
rect 297 147 300 150 
rect 297 150 300 153 
rect 297 153 300 156 
rect 297 156 300 159 
rect 297 159 300 162 
rect 297 162 300 165 
rect 297 165 300 168 
rect 297 168 300 171 
rect 297 171 300 174 
rect 297 174 300 177 
rect 297 177 300 180 
rect 297 180 300 183 
rect 297 183 300 186 
rect 297 186 300 189 
rect 297 189 300 192 
rect 297 192 300 195 
rect 297 195 300 198 
rect 297 198 300 201 
rect 297 201 300 204 
rect 297 204 300 207 
rect 297 207 300 210 
rect 297 210 300 213 
rect 297 213 300 216 
rect 297 216 300 219 
rect 297 219 300 222 
rect 297 222 300 225 
rect 297 225 300 228 
rect 297 228 300 231 
rect 297 231 300 234 
rect 297 234 300 237 
rect 297 237 300 240 
rect 297 240 300 243 
rect 297 243 300 246 
rect 297 246 300 249 
rect 297 249 300 252 
rect 297 252 300 255 
rect 297 255 300 258 
rect 297 258 300 261 
rect 297 261 300 264 
rect 297 264 300 267 
rect 297 267 300 270 
rect 297 270 300 273 
rect 297 273 300 276 
rect 297 276 300 279 
rect 297 279 300 282 
rect 297 282 300 285 
rect 297 285 300 288 
rect 297 288 300 291 
rect 297 291 300 294 
rect 297 294 300 297 
rect 297 297 300 300 
rect 297 300 300 303 
rect 297 303 300 306 
rect 297 306 300 309 
rect 297 309 300 312 
rect 297 312 300 315 
rect 297 315 300 318 
rect 297 318 300 321 
rect 297 321 300 324 
rect 297 324 300 327 
rect 297 327 300 330 
rect 297 330 300 333 
rect 297 333 300 336 
rect 297 336 300 339 
rect 297 339 300 342 
rect 297 342 300 345 
rect 297 345 300 348 
rect 297 348 300 351 
rect 297 351 300 354 
rect 297 354 300 357 
rect 297 357 300 360 
rect 297 360 300 363 
rect 297 363 300 366 
rect 297 366 300 369 
rect 297 369 300 372 
rect 297 372 300 375 
rect 297 375 300 378 
rect 297 378 300 381 
rect 297 381 300 384 
rect 297 384 300 387 
rect 297 387 300 390 
rect 297 390 300 393 
rect 297 393 300 396 
rect 297 396 300 399 
rect 297 399 300 402 
rect 297 402 300 405 
rect 297 405 300 408 
rect 297 408 300 411 
rect 297 411 300 414 
rect 297 414 300 417 
rect 297 417 300 420 
rect 297 420 300 423 
rect 297 423 300 426 
rect 297 426 300 429 
rect 297 429 300 432 
rect 297 432 300 435 
rect 297 435 300 438 
rect 297 438 300 441 
rect 297 441 300 444 
rect 297 444 300 447 
rect 297 447 300 450 
rect 297 450 300 453 
rect 297 453 300 456 
rect 297 456 300 459 
rect 297 459 300 462 
rect 297 462 300 465 
rect 297 465 300 468 
rect 297 468 300 471 
rect 297 471 300 474 
rect 297 474 300 477 
rect 297 477 300 480 
rect 297 480 300 483 
rect 297 483 300 486 
rect 297 486 300 489 
rect 297 489 300 492 
rect 297 492 300 495 
rect 297 495 300 498 
rect 297 498 300 501 
rect 297 501 300 504 
rect 297 504 300 507 
rect 297 507 300 510 
rect 300 0 303 3 
rect 300 3 303 6 
rect 300 6 303 9 
rect 300 9 303 12 
rect 300 12 303 15 
rect 300 15 303 18 
rect 300 18 303 21 
rect 300 21 303 24 
rect 300 24 303 27 
rect 300 27 303 30 
rect 300 30 303 33 
rect 300 33 303 36 
rect 300 36 303 39 
rect 300 39 303 42 
rect 300 42 303 45 
rect 300 45 303 48 
rect 300 48 303 51 
rect 300 51 303 54 
rect 300 54 303 57 
rect 300 57 303 60 
rect 300 60 303 63 
rect 300 63 303 66 
rect 300 66 303 69 
rect 300 69 303 72 
rect 300 72 303 75 
rect 300 75 303 78 
rect 300 78 303 81 
rect 300 81 303 84 
rect 300 84 303 87 
rect 300 87 303 90 
rect 300 90 303 93 
rect 300 93 303 96 
rect 300 96 303 99 
rect 300 99 303 102 
rect 300 102 303 105 
rect 300 105 303 108 
rect 300 108 303 111 
rect 300 111 303 114 
rect 300 114 303 117 
rect 300 117 303 120 
rect 300 120 303 123 
rect 300 123 303 126 
rect 300 126 303 129 
rect 300 129 303 132 
rect 300 132 303 135 
rect 300 135 303 138 
rect 300 138 303 141 
rect 300 141 303 144 
rect 300 144 303 147 
rect 300 147 303 150 
rect 300 150 303 153 
rect 300 153 303 156 
rect 300 156 303 159 
rect 300 159 303 162 
rect 300 162 303 165 
rect 300 165 303 168 
rect 300 168 303 171 
rect 300 171 303 174 
rect 300 174 303 177 
rect 300 177 303 180 
rect 300 180 303 183 
rect 300 183 303 186 
rect 300 186 303 189 
rect 300 189 303 192 
rect 300 192 303 195 
rect 300 195 303 198 
rect 300 198 303 201 
rect 300 201 303 204 
rect 300 204 303 207 
rect 300 207 303 210 
rect 300 210 303 213 
rect 300 213 303 216 
rect 300 216 303 219 
rect 300 219 303 222 
rect 300 222 303 225 
rect 300 225 303 228 
rect 300 228 303 231 
rect 300 231 303 234 
rect 300 234 303 237 
rect 300 237 303 240 
rect 300 240 303 243 
rect 300 243 303 246 
rect 300 246 303 249 
rect 300 249 303 252 
rect 300 252 303 255 
rect 300 255 303 258 
rect 300 258 303 261 
rect 300 261 303 264 
rect 300 264 303 267 
rect 300 267 303 270 
rect 300 270 303 273 
rect 300 273 303 276 
rect 300 276 303 279 
rect 300 279 303 282 
rect 300 282 303 285 
rect 300 285 303 288 
rect 300 288 303 291 
rect 300 291 303 294 
rect 300 294 303 297 
rect 300 297 303 300 
rect 300 300 303 303 
rect 300 303 303 306 
rect 300 306 303 309 
rect 300 309 303 312 
rect 300 312 303 315 
rect 300 315 303 318 
rect 300 318 303 321 
rect 300 321 303 324 
rect 300 324 303 327 
rect 300 327 303 330 
rect 300 330 303 333 
rect 300 333 303 336 
rect 300 336 303 339 
rect 300 339 303 342 
rect 300 342 303 345 
rect 300 345 303 348 
rect 300 348 303 351 
rect 300 351 303 354 
rect 300 354 303 357 
rect 300 357 303 360 
rect 300 360 303 363 
rect 300 363 303 366 
rect 300 366 303 369 
rect 300 369 303 372 
rect 300 372 303 375 
rect 300 375 303 378 
rect 300 378 303 381 
rect 300 381 303 384 
rect 300 384 303 387 
rect 300 387 303 390 
rect 300 390 303 393 
rect 300 393 303 396 
rect 300 396 303 399 
rect 300 399 303 402 
rect 300 402 303 405 
rect 300 405 303 408 
rect 300 408 303 411 
rect 300 411 303 414 
rect 300 414 303 417 
rect 300 417 303 420 
rect 300 420 303 423 
rect 300 423 303 426 
rect 300 426 303 429 
rect 300 429 303 432 
rect 300 432 303 435 
rect 300 435 303 438 
rect 300 438 303 441 
rect 300 441 303 444 
rect 300 444 303 447 
rect 300 447 303 450 
rect 300 450 303 453 
rect 300 453 303 456 
rect 300 456 303 459 
rect 300 459 303 462 
rect 300 462 303 465 
rect 300 465 303 468 
rect 300 468 303 471 
rect 300 471 303 474 
rect 300 474 303 477 
rect 300 477 303 480 
rect 300 480 303 483 
rect 300 483 303 486 
rect 300 486 303 489 
rect 300 489 303 492 
rect 300 492 303 495 
rect 300 495 303 498 
rect 300 498 303 501 
rect 300 501 303 504 
rect 300 504 303 507 
rect 300 507 303 510 
rect 303 0 306 3 
rect 303 3 306 6 
rect 303 6 306 9 
rect 303 9 306 12 
rect 303 12 306 15 
rect 303 15 306 18 
rect 303 18 306 21 
rect 303 21 306 24 
rect 303 24 306 27 
rect 303 27 306 30 
rect 303 30 306 33 
rect 303 33 306 36 
rect 303 36 306 39 
rect 303 39 306 42 
rect 303 42 306 45 
rect 303 45 306 48 
rect 303 48 306 51 
rect 303 51 306 54 
rect 303 54 306 57 
rect 303 57 306 60 
rect 303 60 306 63 
rect 303 63 306 66 
rect 303 66 306 69 
rect 303 69 306 72 
rect 303 72 306 75 
rect 303 75 306 78 
rect 303 78 306 81 
rect 303 81 306 84 
rect 303 84 306 87 
rect 303 87 306 90 
rect 303 90 306 93 
rect 303 93 306 96 
rect 303 96 306 99 
rect 303 99 306 102 
rect 303 102 306 105 
rect 303 105 306 108 
rect 303 108 306 111 
rect 303 111 306 114 
rect 303 114 306 117 
rect 303 117 306 120 
rect 303 120 306 123 
rect 303 123 306 126 
rect 303 126 306 129 
rect 303 129 306 132 
rect 303 132 306 135 
rect 303 135 306 138 
rect 303 138 306 141 
rect 303 141 306 144 
rect 303 144 306 147 
rect 303 147 306 150 
rect 303 150 306 153 
rect 303 153 306 156 
rect 303 156 306 159 
rect 303 159 306 162 
rect 303 162 306 165 
rect 303 165 306 168 
rect 303 168 306 171 
rect 303 171 306 174 
rect 303 174 306 177 
rect 303 177 306 180 
rect 303 180 306 183 
rect 303 183 306 186 
rect 303 186 306 189 
rect 303 189 306 192 
rect 303 192 306 195 
rect 303 195 306 198 
rect 303 198 306 201 
rect 303 201 306 204 
rect 303 204 306 207 
rect 303 207 306 210 
rect 303 210 306 213 
rect 303 213 306 216 
rect 303 216 306 219 
rect 303 219 306 222 
rect 303 222 306 225 
rect 303 225 306 228 
rect 303 228 306 231 
rect 303 231 306 234 
rect 303 234 306 237 
rect 303 237 306 240 
rect 303 240 306 243 
rect 303 243 306 246 
rect 303 246 306 249 
rect 303 249 306 252 
rect 303 252 306 255 
rect 303 255 306 258 
rect 303 258 306 261 
rect 303 261 306 264 
rect 303 264 306 267 
rect 303 267 306 270 
rect 303 270 306 273 
rect 303 273 306 276 
rect 303 276 306 279 
rect 303 279 306 282 
rect 303 282 306 285 
rect 303 285 306 288 
rect 303 288 306 291 
rect 303 291 306 294 
rect 303 294 306 297 
rect 303 297 306 300 
rect 303 300 306 303 
rect 303 303 306 306 
rect 303 306 306 309 
rect 303 309 306 312 
rect 303 312 306 315 
rect 303 315 306 318 
rect 303 318 306 321 
rect 303 321 306 324 
rect 303 324 306 327 
rect 303 327 306 330 
rect 303 330 306 333 
rect 303 333 306 336 
rect 303 336 306 339 
rect 303 339 306 342 
rect 303 342 306 345 
rect 303 345 306 348 
rect 303 348 306 351 
rect 303 351 306 354 
rect 303 354 306 357 
rect 303 357 306 360 
rect 303 360 306 363 
rect 303 363 306 366 
rect 303 366 306 369 
rect 303 369 306 372 
rect 303 372 306 375 
rect 303 375 306 378 
rect 303 378 306 381 
rect 303 381 306 384 
rect 303 384 306 387 
rect 303 387 306 390 
rect 303 390 306 393 
rect 303 393 306 396 
rect 303 396 306 399 
rect 303 399 306 402 
rect 303 402 306 405 
rect 303 405 306 408 
rect 303 408 306 411 
rect 303 411 306 414 
rect 303 414 306 417 
rect 303 417 306 420 
rect 303 420 306 423 
rect 303 423 306 426 
rect 303 426 306 429 
rect 303 429 306 432 
rect 303 432 306 435 
rect 303 435 306 438 
rect 303 438 306 441 
rect 303 441 306 444 
rect 303 444 306 447 
rect 303 447 306 450 
rect 303 450 306 453 
rect 303 453 306 456 
rect 303 456 306 459 
rect 303 459 306 462 
rect 303 462 306 465 
rect 303 465 306 468 
rect 303 468 306 471 
rect 303 471 306 474 
rect 303 474 306 477 
rect 303 477 306 480 
rect 303 480 306 483 
rect 303 483 306 486 
rect 303 486 306 489 
rect 303 489 306 492 
rect 303 492 306 495 
rect 303 495 306 498 
rect 303 498 306 501 
rect 303 501 306 504 
rect 303 504 306 507 
rect 303 507 306 510 
rect 306 0 309 3 
rect 306 3 309 6 
rect 306 6 309 9 
rect 306 9 309 12 
rect 306 12 309 15 
rect 306 15 309 18 
rect 306 18 309 21 
rect 306 21 309 24 
rect 306 24 309 27 
rect 306 27 309 30 
rect 306 30 309 33 
rect 306 33 309 36 
rect 306 36 309 39 
rect 306 39 309 42 
rect 306 42 309 45 
rect 306 45 309 48 
rect 306 48 309 51 
rect 306 51 309 54 
rect 306 54 309 57 
rect 306 57 309 60 
rect 306 60 309 63 
rect 306 63 309 66 
rect 306 66 309 69 
rect 306 69 309 72 
rect 306 72 309 75 
rect 306 75 309 78 
rect 306 78 309 81 
rect 306 81 309 84 
rect 306 84 309 87 
rect 306 87 309 90 
rect 306 90 309 93 
rect 306 93 309 96 
rect 306 96 309 99 
rect 306 99 309 102 
rect 306 102 309 105 
rect 306 105 309 108 
rect 306 108 309 111 
rect 306 111 309 114 
rect 306 114 309 117 
rect 306 117 309 120 
rect 306 120 309 123 
rect 306 123 309 126 
rect 306 126 309 129 
rect 306 129 309 132 
rect 306 132 309 135 
rect 306 135 309 138 
rect 306 138 309 141 
rect 306 141 309 144 
rect 306 144 309 147 
rect 306 147 309 150 
rect 306 150 309 153 
rect 306 153 309 156 
rect 306 156 309 159 
rect 306 159 309 162 
rect 306 162 309 165 
rect 306 165 309 168 
rect 306 168 309 171 
rect 306 171 309 174 
rect 306 174 309 177 
rect 306 177 309 180 
rect 306 180 309 183 
rect 306 183 309 186 
rect 306 186 309 189 
rect 306 189 309 192 
rect 306 192 309 195 
rect 306 195 309 198 
rect 306 198 309 201 
rect 306 201 309 204 
rect 306 204 309 207 
rect 306 207 309 210 
rect 306 210 309 213 
rect 306 213 309 216 
rect 306 216 309 219 
rect 306 219 309 222 
rect 306 222 309 225 
rect 306 225 309 228 
rect 306 228 309 231 
rect 306 231 309 234 
rect 306 234 309 237 
rect 306 237 309 240 
rect 306 240 309 243 
rect 306 243 309 246 
rect 306 246 309 249 
rect 306 249 309 252 
rect 306 252 309 255 
rect 306 255 309 258 
rect 306 258 309 261 
rect 306 261 309 264 
rect 306 264 309 267 
rect 306 267 309 270 
rect 306 270 309 273 
rect 306 273 309 276 
rect 306 276 309 279 
rect 306 279 309 282 
rect 306 282 309 285 
rect 306 285 309 288 
rect 306 288 309 291 
rect 306 291 309 294 
rect 306 294 309 297 
rect 306 297 309 300 
rect 306 300 309 303 
rect 306 303 309 306 
rect 306 306 309 309 
rect 306 309 309 312 
rect 306 312 309 315 
rect 306 315 309 318 
rect 306 318 309 321 
rect 306 321 309 324 
rect 306 324 309 327 
rect 306 327 309 330 
rect 306 330 309 333 
rect 306 333 309 336 
rect 306 336 309 339 
rect 306 339 309 342 
rect 306 342 309 345 
rect 306 345 309 348 
rect 306 348 309 351 
rect 306 351 309 354 
rect 306 354 309 357 
rect 306 357 309 360 
rect 306 360 309 363 
rect 306 363 309 366 
rect 306 366 309 369 
rect 306 369 309 372 
rect 306 372 309 375 
rect 306 375 309 378 
rect 306 378 309 381 
rect 306 381 309 384 
rect 306 384 309 387 
rect 306 387 309 390 
rect 306 390 309 393 
rect 306 393 309 396 
rect 306 396 309 399 
rect 306 399 309 402 
rect 306 402 309 405 
rect 306 405 309 408 
rect 306 408 309 411 
rect 306 411 309 414 
rect 306 414 309 417 
rect 306 417 309 420 
rect 306 420 309 423 
rect 306 423 309 426 
rect 306 426 309 429 
rect 306 429 309 432 
rect 306 432 309 435 
rect 306 435 309 438 
rect 306 438 309 441 
rect 306 441 309 444 
rect 306 444 309 447 
rect 306 447 309 450 
rect 306 450 309 453 
rect 306 453 309 456 
rect 306 456 309 459 
rect 306 459 309 462 
rect 306 462 309 465 
rect 306 465 309 468 
rect 306 468 309 471 
rect 306 471 309 474 
rect 306 474 309 477 
rect 306 477 309 480 
rect 306 480 309 483 
rect 306 483 309 486 
rect 306 486 309 489 
rect 306 489 309 492 
rect 306 492 309 495 
rect 306 495 309 498 
rect 306 498 309 501 
rect 306 501 309 504 
rect 306 504 309 507 
rect 306 507 309 510 
rect 309 0 312 3 
rect 309 3 312 6 
rect 309 6 312 9 
rect 309 9 312 12 
rect 309 12 312 15 
rect 309 15 312 18 
rect 309 18 312 21 
rect 309 21 312 24 
rect 309 24 312 27 
rect 309 27 312 30 
rect 309 30 312 33 
rect 309 33 312 36 
rect 309 36 312 39 
rect 309 39 312 42 
rect 309 42 312 45 
rect 309 45 312 48 
rect 309 48 312 51 
rect 309 51 312 54 
rect 309 54 312 57 
rect 309 57 312 60 
rect 309 60 312 63 
rect 309 63 312 66 
rect 309 66 312 69 
rect 309 69 312 72 
rect 309 72 312 75 
rect 309 75 312 78 
rect 309 78 312 81 
rect 309 81 312 84 
rect 309 84 312 87 
rect 309 87 312 90 
rect 309 90 312 93 
rect 309 93 312 96 
rect 309 96 312 99 
rect 309 99 312 102 
rect 309 102 312 105 
rect 309 105 312 108 
rect 309 108 312 111 
rect 309 111 312 114 
rect 309 114 312 117 
rect 309 117 312 120 
rect 309 120 312 123 
rect 309 123 312 126 
rect 309 126 312 129 
rect 309 129 312 132 
rect 309 132 312 135 
rect 309 135 312 138 
rect 309 138 312 141 
rect 309 141 312 144 
rect 309 144 312 147 
rect 309 147 312 150 
rect 309 150 312 153 
rect 309 153 312 156 
rect 309 156 312 159 
rect 309 159 312 162 
rect 309 162 312 165 
rect 309 165 312 168 
rect 309 168 312 171 
rect 309 171 312 174 
rect 309 174 312 177 
rect 309 177 312 180 
rect 309 180 312 183 
rect 309 183 312 186 
rect 309 186 312 189 
rect 309 189 312 192 
rect 309 192 312 195 
rect 309 195 312 198 
rect 309 198 312 201 
rect 309 201 312 204 
rect 309 204 312 207 
rect 309 207 312 210 
rect 309 210 312 213 
rect 309 213 312 216 
rect 309 216 312 219 
rect 309 219 312 222 
rect 309 222 312 225 
rect 309 225 312 228 
rect 309 228 312 231 
rect 309 231 312 234 
rect 309 234 312 237 
rect 309 237 312 240 
rect 309 240 312 243 
rect 309 243 312 246 
rect 309 246 312 249 
rect 309 249 312 252 
rect 309 252 312 255 
rect 309 255 312 258 
rect 309 258 312 261 
rect 309 261 312 264 
rect 309 264 312 267 
rect 309 267 312 270 
rect 309 270 312 273 
rect 309 273 312 276 
rect 309 276 312 279 
rect 309 279 312 282 
rect 309 282 312 285 
rect 309 285 312 288 
rect 309 288 312 291 
rect 309 291 312 294 
rect 309 294 312 297 
rect 309 297 312 300 
rect 309 300 312 303 
rect 309 303 312 306 
rect 309 306 312 309 
rect 309 309 312 312 
rect 309 312 312 315 
rect 309 315 312 318 
rect 309 318 312 321 
rect 309 321 312 324 
rect 309 324 312 327 
rect 309 327 312 330 
rect 309 330 312 333 
rect 309 333 312 336 
rect 309 336 312 339 
rect 309 339 312 342 
rect 309 342 312 345 
rect 309 345 312 348 
rect 309 348 312 351 
rect 309 351 312 354 
rect 309 354 312 357 
rect 309 357 312 360 
rect 309 360 312 363 
rect 309 363 312 366 
rect 309 366 312 369 
rect 309 369 312 372 
rect 309 372 312 375 
rect 309 375 312 378 
rect 309 378 312 381 
rect 309 381 312 384 
rect 309 384 312 387 
rect 309 387 312 390 
rect 309 390 312 393 
rect 309 393 312 396 
rect 309 396 312 399 
rect 309 399 312 402 
rect 309 402 312 405 
rect 309 405 312 408 
rect 309 408 312 411 
rect 309 411 312 414 
rect 309 414 312 417 
rect 309 417 312 420 
rect 309 420 312 423 
rect 309 423 312 426 
rect 309 426 312 429 
rect 309 429 312 432 
rect 309 432 312 435 
rect 309 435 312 438 
rect 309 438 312 441 
rect 309 441 312 444 
rect 309 444 312 447 
rect 309 447 312 450 
rect 309 450 312 453 
rect 309 453 312 456 
rect 309 456 312 459 
rect 309 459 312 462 
rect 309 462 312 465 
rect 309 465 312 468 
rect 309 468 312 471 
rect 309 471 312 474 
rect 309 474 312 477 
rect 309 477 312 480 
rect 309 480 312 483 
rect 309 483 312 486 
rect 309 486 312 489 
rect 309 489 312 492 
rect 309 492 312 495 
rect 309 495 312 498 
rect 309 498 312 501 
rect 309 501 312 504 
rect 309 504 312 507 
rect 309 507 312 510 
rect 312 0 315 3 
rect 312 3 315 6 
rect 312 6 315 9 
rect 312 9 315 12 
rect 312 12 315 15 
rect 312 15 315 18 
rect 312 18 315 21 
rect 312 21 315 24 
rect 312 24 315 27 
rect 312 27 315 30 
rect 312 30 315 33 
rect 312 33 315 36 
rect 312 36 315 39 
rect 312 39 315 42 
rect 312 42 315 45 
rect 312 45 315 48 
rect 312 48 315 51 
rect 312 51 315 54 
rect 312 54 315 57 
rect 312 57 315 60 
rect 312 60 315 63 
rect 312 63 315 66 
rect 312 66 315 69 
rect 312 69 315 72 
rect 312 72 315 75 
rect 312 75 315 78 
rect 312 78 315 81 
rect 312 81 315 84 
rect 312 84 315 87 
rect 312 87 315 90 
rect 312 90 315 93 
rect 312 93 315 96 
rect 312 96 315 99 
rect 312 99 315 102 
rect 312 102 315 105 
rect 312 105 315 108 
rect 312 108 315 111 
rect 312 111 315 114 
rect 312 114 315 117 
rect 312 117 315 120 
rect 312 120 315 123 
rect 312 123 315 126 
rect 312 126 315 129 
rect 312 129 315 132 
rect 312 132 315 135 
rect 312 135 315 138 
rect 312 138 315 141 
rect 312 141 315 144 
rect 312 144 315 147 
rect 312 147 315 150 
rect 312 150 315 153 
rect 312 153 315 156 
rect 312 156 315 159 
rect 312 159 315 162 
rect 312 162 315 165 
rect 312 165 315 168 
rect 312 168 315 171 
rect 312 171 315 174 
rect 312 174 315 177 
rect 312 177 315 180 
rect 312 180 315 183 
rect 312 183 315 186 
rect 312 186 315 189 
rect 312 189 315 192 
rect 312 192 315 195 
rect 312 195 315 198 
rect 312 198 315 201 
rect 312 201 315 204 
rect 312 204 315 207 
rect 312 207 315 210 
rect 312 210 315 213 
rect 312 213 315 216 
rect 312 216 315 219 
rect 312 219 315 222 
rect 312 222 315 225 
rect 312 225 315 228 
rect 312 228 315 231 
rect 312 231 315 234 
rect 312 234 315 237 
rect 312 237 315 240 
rect 312 240 315 243 
rect 312 243 315 246 
rect 312 246 315 249 
rect 312 249 315 252 
rect 312 252 315 255 
rect 312 255 315 258 
rect 312 258 315 261 
rect 312 261 315 264 
rect 312 264 315 267 
rect 312 267 315 270 
rect 312 270 315 273 
rect 312 273 315 276 
rect 312 276 315 279 
rect 312 279 315 282 
rect 312 282 315 285 
rect 312 285 315 288 
rect 312 288 315 291 
rect 312 291 315 294 
rect 312 294 315 297 
rect 312 297 315 300 
rect 312 300 315 303 
rect 312 303 315 306 
rect 312 306 315 309 
rect 312 309 315 312 
rect 312 312 315 315 
rect 312 315 315 318 
rect 312 318 315 321 
rect 312 321 315 324 
rect 312 324 315 327 
rect 312 327 315 330 
rect 312 330 315 333 
rect 312 333 315 336 
rect 312 336 315 339 
rect 312 339 315 342 
rect 312 342 315 345 
rect 312 345 315 348 
rect 312 348 315 351 
rect 312 351 315 354 
rect 312 354 315 357 
rect 312 357 315 360 
rect 312 360 315 363 
rect 312 363 315 366 
rect 312 366 315 369 
rect 312 369 315 372 
rect 312 372 315 375 
rect 312 375 315 378 
rect 312 378 315 381 
rect 312 381 315 384 
rect 312 384 315 387 
rect 312 387 315 390 
rect 312 390 315 393 
rect 312 393 315 396 
rect 312 396 315 399 
rect 312 399 315 402 
rect 312 402 315 405 
rect 312 405 315 408 
rect 312 408 315 411 
rect 312 411 315 414 
rect 312 414 315 417 
rect 312 417 315 420 
rect 312 420 315 423 
rect 312 423 315 426 
rect 312 426 315 429 
rect 312 429 315 432 
rect 312 432 315 435 
rect 312 435 315 438 
rect 312 438 315 441 
rect 312 441 315 444 
rect 312 444 315 447 
rect 312 447 315 450 
rect 312 450 315 453 
rect 312 453 315 456 
rect 312 456 315 459 
rect 312 459 315 462 
rect 312 462 315 465 
rect 312 465 315 468 
rect 312 468 315 471 
rect 312 471 315 474 
rect 312 474 315 477 
rect 312 477 315 480 
rect 312 480 315 483 
rect 312 483 315 486 
rect 312 486 315 489 
rect 312 489 315 492 
rect 312 492 315 495 
rect 312 495 315 498 
rect 312 498 315 501 
rect 312 501 315 504 
rect 312 504 315 507 
rect 312 507 315 510 
rect 315 0 318 3 
rect 315 3 318 6 
rect 315 6 318 9 
rect 315 9 318 12 
rect 315 12 318 15 
rect 315 15 318 18 
rect 315 18 318 21 
rect 315 21 318 24 
rect 315 24 318 27 
rect 315 27 318 30 
rect 315 30 318 33 
rect 315 33 318 36 
rect 315 36 318 39 
rect 315 39 318 42 
rect 315 42 318 45 
rect 315 45 318 48 
rect 315 48 318 51 
rect 315 51 318 54 
rect 315 54 318 57 
rect 315 57 318 60 
rect 315 60 318 63 
rect 315 63 318 66 
rect 315 66 318 69 
rect 315 69 318 72 
rect 315 72 318 75 
rect 315 75 318 78 
rect 315 78 318 81 
rect 315 81 318 84 
rect 315 84 318 87 
rect 315 87 318 90 
rect 315 90 318 93 
rect 315 93 318 96 
rect 315 96 318 99 
rect 315 99 318 102 
rect 315 102 318 105 
rect 315 105 318 108 
rect 315 108 318 111 
rect 315 111 318 114 
rect 315 114 318 117 
rect 315 117 318 120 
rect 315 120 318 123 
rect 315 123 318 126 
rect 315 126 318 129 
rect 315 129 318 132 
rect 315 132 318 135 
rect 315 135 318 138 
rect 315 138 318 141 
rect 315 141 318 144 
rect 315 144 318 147 
rect 315 147 318 150 
rect 315 150 318 153 
rect 315 153 318 156 
rect 315 156 318 159 
rect 315 159 318 162 
rect 315 162 318 165 
rect 315 165 318 168 
rect 315 168 318 171 
rect 315 171 318 174 
rect 315 174 318 177 
rect 315 177 318 180 
rect 315 180 318 183 
rect 315 183 318 186 
rect 315 186 318 189 
rect 315 189 318 192 
rect 315 192 318 195 
rect 315 195 318 198 
rect 315 198 318 201 
rect 315 201 318 204 
rect 315 204 318 207 
rect 315 207 318 210 
rect 315 210 318 213 
rect 315 213 318 216 
rect 315 216 318 219 
rect 315 219 318 222 
rect 315 222 318 225 
rect 315 225 318 228 
rect 315 228 318 231 
rect 315 231 318 234 
rect 315 234 318 237 
rect 315 237 318 240 
rect 315 240 318 243 
rect 315 243 318 246 
rect 315 246 318 249 
rect 315 249 318 252 
rect 315 252 318 255 
rect 315 255 318 258 
rect 315 258 318 261 
rect 315 261 318 264 
rect 315 264 318 267 
rect 315 267 318 270 
rect 315 270 318 273 
rect 315 273 318 276 
rect 315 276 318 279 
rect 315 279 318 282 
rect 315 282 318 285 
rect 315 285 318 288 
rect 315 288 318 291 
rect 315 291 318 294 
rect 315 294 318 297 
rect 315 297 318 300 
rect 315 300 318 303 
rect 315 303 318 306 
rect 315 306 318 309 
rect 315 309 318 312 
rect 315 312 318 315 
rect 315 315 318 318 
rect 315 318 318 321 
rect 315 321 318 324 
rect 315 324 318 327 
rect 315 327 318 330 
rect 315 330 318 333 
rect 315 333 318 336 
rect 315 336 318 339 
rect 315 339 318 342 
rect 315 342 318 345 
rect 315 345 318 348 
rect 315 348 318 351 
rect 315 351 318 354 
rect 315 354 318 357 
rect 315 357 318 360 
rect 315 360 318 363 
rect 315 363 318 366 
rect 315 366 318 369 
rect 315 369 318 372 
rect 315 372 318 375 
rect 315 375 318 378 
rect 315 378 318 381 
rect 315 381 318 384 
rect 315 384 318 387 
rect 315 387 318 390 
rect 315 390 318 393 
rect 315 393 318 396 
rect 315 396 318 399 
rect 315 399 318 402 
rect 315 402 318 405 
rect 315 405 318 408 
rect 315 408 318 411 
rect 315 411 318 414 
rect 315 414 318 417 
rect 315 417 318 420 
rect 315 420 318 423 
rect 315 423 318 426 
rect 315 426 318 429 
rect 315 429 318 432 
rect 315 432 318 435 
rect 315 435 318 438 
rect 315 438 318 441 
rect 315 441 318 444 
rect 315 444 318 447 
rect 315 447 318 450 
rect 315 450 318 453 
rect 315 453 318 456 
rect 315 456 318 459 
rect 315 459 318 462 
rect 315 462 318 465 
rect 315 465 318 468 
rect 315 468 318 471 
rect 315 471 318 474 
rect 315 474 318 477 
rect 315 477 318 480 
rect 315 480 318 483 
rect 315 483 318 486 
rect 315 486 318 489 
rect 315 489 318 492 
rect 315 492 318 495 
rect 315 495 318 498 
rect 315 498 318 501 
rect 315 501 318 504 
rect 315 504 318 507 
rect 315 507 318 510 
rect 318 0 321 3 
rect 318 3 321 6 
rect 318 6 321 9 
rect 318 9 321 12 
rect 318 12 321 15 
rect 318 15 321 18 
rect 318 18 321 21 
rect 318 21 321 24 
rect 318 24 321 27 
rect 318 27 321 30 
rect 318 30 321 33 
rect 318 33 321 36 
rect 318 36 321 39 
rect 318 39 321 42 
rect 318 42 321 45 
rect 318 45 321 48 
rect 318 48 321 51 
rect 318 51 321 54 
rect 318 54 321 57 
rect 318 57 321 60 
rect 318 60 321 63 
rect 318 63 321 66 
rect 318 66 321 69 
rect 318 69 321 72 
rect 318 72 321 75 
rect 318 75 321 78 
rect 318 78 321 81 
rect 318 81 321 84 
rect 318 84 321 87 
rect 318 87 321 90 
rect 318 90 321 93 
rect 318 93 321 96 
rect 318 96 321 99 
rect 318 99 321 102 
rect 318 102 321 105 
rect 318 105 321 108 
rect 318 108 321 111 
rect 318 111 321 114 
rect 318 114 321 117 
rect 318 117 321 120 
rect 318 120 321 123 
rect 318 123 321 126 
rect 318 126 321 129 
rect 318 129 321 132 
rect 318 132 321 135 
rect 318 135 321 138 
rect 318 138 321 141 
rect 318 141 321 144 
rect 318 144 321 147 
rect 318 147 321 150 
rect 318 150 321 153 
rect 318 153 321 156 
rect 318 156 321 159 
rect 318 159 321 162 
rect 318 162 321 165 
rect 318 165 321 168 
rect 318 168 321 171 
rect 318 171 321 174 
rect 318 174 321 177 
rect 318 177 321 180 
rect 318 180 321 183 
rect 318 183 321 186 
rect 318 186 321 189 
rect 318 189 321 192 
rect 318 192 321 195 
rect 318 195 321 198 
rect 318 198 321 201 
rect 318 201 321 204 
rect 318 204 321 207 
rect 318 207 321 210 
rect 318 210 321 213 
rect 318 213 321 216 
rect 318 216 321 219 
rect 318 219 321 222 
rect 318 222 321 225 
rect 318 225 321 228 
rect 318 228 321 231 
rect 318 231 321 234 
rect 318 234 321 237 
rect 318 237 321 240 
rect 318 240 321 243 
rect 318 243 321 246 
rect 318 246 321 249 
rect 318 249 321 252 
rect 318 252 321 255 
rect 318 255 321 258 
rect 318 258 321 261 
rect 318 261 321 264 
rect 318 264 321 267 
rect 318 267 321 270 
rect 318 270 321 273 
rect 318 273 321 276 
rect 318 276 321 279 
rect 318 279 321 282 
rect 318 282 321 285 
rect 318 285 321 288 
rect 318 288 321 291 
rect 318 291 321 294 
rect 318 294 321 297 
rect 318 297 321 300 
rect 318 300 321 303 
rect 318 303 321 306 
rect 318 306 321 309 
rect 318 309 321 312 
rect 318 312 321 315 
rect 318 315 321 318 
rect 318 318 321 321 
rect 318 321 321 324 
rect 318 324 321 327 
rect 318 327 321 330 
rect 318 330 321 333 
rect 318 333 321 336 
rect 318 336 321 339 
rect 318 339 321 342 
rect 318 342 321 345 
rect 318 345 321 348 
rect 318 348 321 351 
rect 318 351 321 354 
rect 318 354 321 357 
rect 318 357 321 360 
rect 318 360 321 363 
rect 318 363 321 366 
rect 318 366 321 369 
rect 318 369 321 372 
rect 318 372 321 375 
rect 318 375 321 378 
rect 318 378 321 381 
rect 318 381 321 384 
rect 318 384 321 387 
rect 318 387 321 390 
rect 318 390 321 393 
rect 318 393 321 396 
rect 318 396 321 399 
rect 318 399 321 402 
rect 318 402 321 405 
rect 318 405 321 408 
rect 318 408 321 411 
rect 318 411 321 414 
rect 318 414 321 417 
rect 318 417 321 420 
rect 318 420 321 423 
rect 318 423 321 426 
rect 318 426 321 429 
rect 318 429 321 432 
rect 318 432 321 435 
rect 318 435 321 438 
rect 318 438 321 441 
rect 318 441 321 444 
rect 318 444 321 447 
rect 318 447 321 450 
rect 318 450 321 453 
rect 318 453 321 456 
rect 318 456 321 459 
rect 318 459 321 462 
rect 318 462 321 465 
rect 318 465 321 468 
rect 318 468 321 471 
rect 318 471 321 474 
rect 318 474 321 477 
rect 318 477 321 480 
rect 318 480 321 483 
rect 318 483 321 486 
rect 318 486 321 489 
rect 318 489 321 492 
rect 318 492 321 495 
rect 318 495 321 498 
rect 318 498 321 501 
rect 318 501 321 504 
rect 318 504 321 507 
rect 318 507 321 510 
rect 321 0 324 3 
rect 321 3 324 6 
rect 321 6 324 9 
rect 321 9 324 12 
rect 321 12 324 15 
rect 321 15 324 18 
rect 321 18 324 21 
rect 321 21 324 24 
rect 321 24 324 27 
rect 321 27 324 30 
rect 321 30 324 33 
rect 321 33 324 36 
rect 321 36 324 39 
rect 321 39 324 42 
rect 321 42 324 45 
rect 321 45 324 48 
rect 321 48 324 51 
rect 321 51 324 54 
rect 321 54 324 57 
rect 321 57 324 60 
rect 321 60 324 63 
rect 321 63 324 66 
rect 321 66 324 69 
rect 321 69 324 72 
rect 321 72 324 75 
rect 321 75 324 78 
rect 321 78 324 81 
rect 321 81 324 84 
rect 321 84 324 87 
rect 321 87 324 90 
rect 321 90 324 93 
rect 321 93 324 96 
rect 321 96 324 99 
rect 321 99 324 102 
rect 321 102 324 105 
rect 321 105 324 108 
rect 321 108 324 111 
rect 321 111 324 114 
rect 321 114 324 117 
rect 321 117 324 120 
rect 321 120 324 123 
rect 321 123 324 126 
rect 321 126 324 129 
rect 321 129 324 132 
rect 321 132 324 135 
rect 321 135 324 138 
rect 321 138 324 141 
rect 321 141 324 144 
rect 321 144 324 147 
rect 321 147 324 150 
rect 321 150 324 153 
rect 321 153 324 156 
rect 321 156 324 159 
rect 321 159 324 162 
rect 321 162 324 165 
rect 321 165 324 168 
rect 321 168 324 171 
rect 321 171 324 174 
rect 321 174 324 177 
rect 321 177 324 180 
rect 321 180 324 183 
rect 321 183 324 186 
rect 321 186 324 189 
rect 321 189 324 192 
rect 321 192 324 195 
rect 321 195 324 198 
rect 321 198 324 201 
rect 321 201 324 204 
rect 321 204 324 207 
rect 321 207 324 210 
rect 321 210 324 213 
rect 321 213 324 216 
rect 321 216 324 219 
rect 321 219 324 222 
rect 321 222 324 225 
rect 321 225 324 228 
rect 321 228 324 231 
rect 321 231 324 234 
rect 321 234 324 237 
rect 321 237 324 240 
rect 321 240 324 243 
rect 321 243 324 246 
rect 321 246 324 249 
rect 321 249 324 252 
rect 321 252 324 255 
rect 321 255 324 258 
rect 321 258 324 261 
rect 321 261 324 264 
rect 321 264 324 267 
rect 321 267 324 270 
rect 321 270 324 273 
rect 321 273 324 276 
rect 321 276 324 279 
rect 321 279 324 282 
rect 321 282 324 285 
rect 321 285 324 288 
rect 321 288 324 291 
rect 321 291 324 294 
rect 321 294 324 297 
rect 321 297 324 300 
rect 321 300 324 303 
rect 321 303 324 306 
rect 321 306 324 309 
rect 321 309 324 312 
rect 321 312 324 315 
rect 321 315 324 318 
rect 321 318 324 321 
rect 321 321 324 324 
rect 321 324 324 327 
rect 321 327 324 330 
rect 321 330 324 333 
rect 321 333 324 336 
rect 321 336 324 339 
rect 321 339 324 342 
rect 321 342 324 345 
rect 321 345 324 348 
rect 321 348 324 351 
rect 321 351 324 354 
rect 321 354 324 357 
rect 321 357 324 360 
rect 321 360 324 363 
rect 321 363 324 366 
rect 321 366 324 369 
rect 321 369 324 372 
rect 321 372 324 375 
rect 321 375 324 378 
rect 321 378 324 381 
rect 321 381 324 384 
rect 321 384 324 387 
rect 321 387 324 390 
rect 321 390 324 393 
rect 321 393 324 396 
rect 321 396 324 399 
rect 321 399 324 402 
rect 321 402 324 405 
rect 321 405 324 408 
rect 321 408 324 411 
rect 321 411 324 414 
rect 321 414 324 417 
rect 321 417 324 420 
rect 321 420 324 423 
rect 321 423 324 426 
rect 321 426 324 429 
rect 321 429 324 432 
rect 321 432 324 435 
rect 321 435 324 438 
rect 321 438 324 441 
rect 321 441 324 444 
rect 321 444 324 447 
rect 321 447 324 450 
rect 321 450 324 453 
rect 321 453 324 456 
rect 321 456 324 459 
rect 321 459 324 462 
rect 321 462 324 465 
rect 321 465 324 468 
rect 321 468 324 471 
rect 321 471 324 474 
rect 321 474 324 477 
rect 321 477 324 480 
rect 321 480 324 483 
rect 321 483 324 486 
rect 321 486 324 489 
rect 321 489 324 492 
rect 321 492 324 495 
rect 321 495 324 498 
rect 321 498 324 501 
rect 321 501 324 504 
rect 321 504 324 507 
rect 321 507 324 510 
rect 324 0 327 3 
rect 324 3 327 6 
rect 324 6 327 9 
rect 324 9 327 12 
rect 324 12 327 15 
rect 324 15 327 18 
rect 324 18 327 21 
rect 324 21 327 24 
rect 324 24 327 27 
rect 324 27 327 30 
rect 324 30 327 33 
rect 324 33 327 36 
rect 324 36 327 39 
rect 324 39 327 42 
rect 324 42 327 45 
rect 324 45 327 48 
rect 324 48 327 51 
rect 324 51 327 54 
rect 324 54 327 57 
rect 324 57 327 60 
rect 324 60 327 63 
rect 324 63 327 66 
rect 324 66 327 69 
rect 324 69 327 72 
rect 324 72 327 75 
rect 324 75 327 78 
rect 324 78 327 81 
rect 324 81 327 84 
rect 324 84 327 87 
rect 324 87 327 90 
rect 324 90 327 93 
rect 324 93 327 96 
rect 324 96 327 99 
rect 324 99 327 102 
rect 324 102 327 105 
rect 324 105 327 108 
rect 324 108 327 111 
rect 324 111 327 114 
rect 324 114 327 117 
rect 324 117 327 120 
rect 324 120 327 123 
rect 324 123 327 126 
rect 324 126 327 129 
rect 324 129 327 132 
rect 324 132 327 135 
rect 324 135 327 138 
rect 324 138 327 141 
rect 324 141 327 144 
rect 324 144 327 147 
rect 324 147 327 150 
rect 324 150 327 153 
rect 324 153 327 156 
rect 324 156 327 159 
rect 324 159 327 162 
rect 324 162 327 165 
rect 324 165 327 168 
rect 324 168 327 171 
rect 324 171 327 174 
rect 324 174 327 177 
rect 324 177 327 180 
rect 324 180 327 183 
rect 324 183 327 186 
rect 324 186 327 189 
rect 324 189 327 192 
rect 324 192 327 195 
rect 324 195 327 198 
rect 324 198 327 201 
rect 324 201 327 204 
rect 324 204 327 207 
rect 324 207 327 210 
rect 324 210 327 213 
rect 324 213 327 216 
rect 324 216 327 219 
rect 324 219 327 222 
rect 324 222 327 225 
rect 324 225 327 228 
rect 324 228 327 231 
rect 324 231 327 234 
rect 324 234 327 237 
rect 324 237 327 240 
rect 324 240 327 243 
rect 324 243 327 246 
rect 324 246 327 249 
rect 324 249 327 252 
rect 324 252 327 255 
rect 324 255 327 258 
rect 324 258 327 261 
rect 324 261 327 264 
rect 324 264 327 267 
rect 324 267 327 270 
rect 324 270 327 273 
rect 324 273 327 276 
rect 324 276 327 279 
rect 324 279 327 282 
rect 324 282 327 285 
rect 324 285 327 288 
rect 324 288 327 291 
rect 324 291 327 294 
rect 324 294 327 297 
rect 324 297 327 300 
rect 324 300 327 303 
rect 324 303 327 306 
rect 324 306 327 309 
rect 324 309 327 312 
rect 324 312 327 315 
rect 324 315 327 318 
rect 324 318 327 321 
rect 324 321 327 324 
rect 324 324 327 327 
rect 324 327 327 330 
rect 324 330 327 333 
rect 324 333 327 336 
rect 324 336 327 339 
rect 324 339 327 342 
rect 324 342 327 345 
rect 324 345 327 348 
rect 324 348 327 351 
rect 324 351 327 354 
rect 324 354 327 357 
rect 324 357 327 360 
rect 324 360 327 363 
rect 324 363 327 366 
rect 324 366 327 369 
rect 324 369 327 372 
rect 324 372 327 375 
rect 324 375 327 378 
rect 324 378 327 381 
rect 324 381 327 384 
rect 324 384 327 387 
rect 324 387 327 390 
rect 324 390 327 393 
rect 324 393 327 396 
rect 324 396 327 399 
rect 324 399 327 402 
rect 324 402 327 405 
rect 324 405 327 408 
rect 324 408 327 411 
rect 324 411 327 414 
rect 324 414 327 417 
rect 324 417 327 420 
rect 324 420 327 423 
rect 324 423 327 426 
rect 324 426 327 429 
rect 324 429 327 432 
rect 324 432 327 435 
rect 324 435 327 438 
rect 324 438 327 441 
rect 324 441 327 444 
rect 324 444 327 447 
rect 324 447 327 450 
rect 324 450 327 453 
rect 324 453 327 456 
rect 324 456 327 459 
rect 324 459 327 462 
rect 324 462 327 465 
rect 324 465 327 468 
rect 324 468 327 471 
rect 324 471 327 474 
rect 324 474 327 477 
rect 324 477 327 480 
rect 324 480 327 483 
rect 324 483 327 486 
rect 324 486 327 489 
rect 324 489 327 492 
rect 324 492 327 495 
rect 324 495 327 498 
rect 324 498 327 501 
rect 324 501 327 504 
rect 324 504 327 507 
rect 324 507 327 510 
rect 327 0 330 3 
rect 327 3 330 6 
rect 327 6 330 9 
rect 327 9 330 12 
rect 327 12 330 15 
rect 327 15 330 18 
rect 327 18 330 21 
rect 327 21 330 24 
rect 327 24 330 27 
rect 327 27 330 30 
rect 327 30 330 33 
rect 327 33 330 36 
rect 327 36 330 39 
rect 327 39 330 42 
rect 327 42 330 45 
rect 327 45 330 48 
rect 327 48 330 51 
rect 327 51 330 54 
rect 327 54 330 57 
rect 327 57 330 60 
rect 327 60 330 63 
rect 327 63 330 66 
rect 327 66 330 69 
rect 327 69 330 72 
rect 327 72 330 75 
rect 327 75 330 78 
rect 327 78 330 81 
rect 327 81 330 84 
rect 327 84 330 87 
rect 327 87 330 90 
rect 327 90 330 93 
rect 327 93 330 96 
rect 327 96 330 99 
rect 327 99 330 102 
rect 327 102 330 105 
rect 327 105 330 108 
rect 327 108 330 111 
rect 327 111 330 114 
rect 327 114 330 117 
rect 327 117 330 120 
rect 327 120 330 123 
rect 327 123 330 126 
rect 327 126 330 129 
rect 327 129 330 132 
rect 327 132 330 135 
rect 327 135 330 138 
rect 327 138 330 141 
rect 327 141 330 144 
rect 327 144 330 147 
rect 327 147 330 150 
rect 327 150 330 153 
rect 327 153 330 156 
rect 327 156 330 159 
rect 327 159 330 162 
rect 327 162 330 165 
rect 327 165 330 168 
rect 327 168 330 171 
rect 327 171 330 174 
rect 327 174 330 177 
rect 327 177 330 180 
rect 327 180 330 183 
rect 327 183 330 186 
rect 327 186 330 189 
rect 327 189 330 192 
rect 327 192 330 195 
rect 327 195 330 198 
rect 327 198 330 201 
rect 327 201 330 204 
rect 327 204 330 207 
rect 327 207 330 210 
rect 327 210 330 213 
rect 327 213 330 216 
rect 327 216 330 219 
rect 327 219 330 222 
rect 327 222 330 225 
rect 327 225 330 228 
rect 327 228 330 231 
rect 327 231 330 234 
rect 327 234 330 237 
rect 327 237 330 240 
rect 327 240 330 243 
rect 327 243 330 246 
rect 327 246 330 249 
rect 327 249 330 252 
rect 327 252 330 255 
rect 327 255 330 258 
rect 327 258 330 261 
rect 327 261 330 264 
rect 327 264 330 267 
rect 327 267 330 270 
rect 327 270 330 273 
rect 327 273 330 276 
rect 327 276 330 279 
rect 327 279 330 282 
rect 327 282 330 285 
rect 327 285 330 288 
rect 327 288 330 291 
rect 327 291 330 294 
rect 327 294 330 297 
rect 327 297 330 300 
rect 327 300 330 303 
rect 327 303 330 306 
rect 327 306 330 309 
rect 327 309 330 312 
rect 327 312 330 315 
rect 327 315 330 318 
rect 327 318 330 321 
rect 327 321 330 324 
rect 327 324 330 327 
rect 327 327 330 330 
rect 327 330 330 333 
rect 327 333 330 336 
rect 327 336 330 339 
rect 327 339 330 342 
rect 327 342 330 345 
rect 327 345 330 348 
rect 327 348 330 351 
rect 327 351 330 354 
rect 327 354 330 357 
rect 327 357 330 360 
rect 327 360 330 363 
rect 327 363 330 366 
rect 327 366 330 369 
rect 327 369 330 372 
rect 327 372 330 375 
rect 327 375 330 378 
rect 327 378 330 381 
rect 327 381 330 384 
rect 327 384 330 387 
rect 327 387 330 390 
rect 327 390 330 393 
rect 327 393 330 396 
rect 327 396 330 399 
rect 327 399 330 402 
rect 327 402 330 405 
rect 327 405 330 408 
rect 327 408 330 411 
rect 327 411 330 414 
rect 327 414 330 417 
rect 327 417 330 420 
rect 327 420 330 423 
rect 327 423 330 426 
rect 327 426 330 429 
rect 327 429 330 432 
rect 327 432 330 435 
rect 327 435 330 438 
rect 327 438 330 441 
rect 327 441 330 444 
rect 327 444 330 447 
rect 327 447 330 450 
rect 327 450 330 453 
rect 327 453 330 456 
rect 327 456 330 459 
rect 327 459 330 462 
rect 327 462 330 465 
rect 327 465 330 468 
rect 327 468 330 471 
rect 327 471 330 474 
rect 327 474 330 477 
rect 327 477 330 480 
rect 327 480 330 483 
rect 327 483 330 486 
rect 327 486 330 489 
rect 327 489 330 492 
rect 327 492 330 495 
rect 327 495 330 498 
rect 327 498 330 501 
rect 327 501 330 504 
rect 327 504 330 507 
rect 327 507 330 510 
rect 330 0 333 3 
rect 330 3 333 6 
rect 330 6 333 9 
rect 330 9 333 12 
rect 330 12 333 15 
rect 330 15 333 18 
rect 330 18 333 21 
rect 330 21 333 24 
rect 330 24 333 27 
rect 330 27 333 30 
rect 330 30 333 33 
rect 330 33 333 36 
rect 330 36 333 39 
rect 330 39 333 42 
rect 330 42 333 45 
rect 330 45 333 48 
rect 330 48 333 51 
rect 330 51 333 54 
rect 330 54 333 57 
rect 330 57 333 60 
rect 330 60 333 63 
rect 330 63 333 66 
rect 330 66 333 69 
rect 330 69 333 72 
rect 330 72 333 75 
rect 330 75 333 78 
rect 330 78 333 81 
rect 330 81 333 84 
rect 330 84 333 87 
rect 330 87 333 90 
rect 330 90 333 93 
rect 330 93 333 96 
rect 330 96 333 99 
rect 330 99 333 102 
rect 330 102 333 105 
rect 330 105 333 108 
rect 330 108 333 111 
rect 330 111 333 114 
rect 330 114 333 117 
rect 330 117 333 120 
rect 330 120 333 123 
rect 330 123 333 126 
rect 330 126 333 129 
rect 330 129 333 132 
rect 330 132 333 135 
rect 330 135 333 138 
rect 330 138 333 141 
rect 330 141 333 144 
rect 330 144 333 147 
rect 330 147 333 150 
rect 330 150 333 153 
rect 330 153 333 156 
rect 330 156 333 159 
rect 330 159 333 162 
rect 330 162 333 165 
rect 330 165 333 168 
rect 330 168 333 171 
rect 330 171 333 174 
rect 330 174 333 177 
rect 330 177 333 180 
rect 330 180 333 183 
rect 330 183 333 186 
rect 330 186 333 189 
rect 330 189 333 192 
rect 330 192 333 195 
rect 330 195 333 198 
rect 330 198 333 201 
rect 330 201 333 204 
rect 330 204 333 207 
rect 330 207 333 210 
rect 330 210 333 213 
rect 330 213 333 216 
rect 330 216 333 219 
rect 330 219 333 222 
rect 330 222 333 225 
rect 330 225 333 228 
rect 330 228 333 231 
rect 330 231 333 234 
rect 330 234 333 237 
rect 330 237 333 240 
rect 330 240 333 243 
rect 330 243 333 246 
rect 330 246 333 249 
rect 330 249 333 252 
rect 330 252 333 255 
rect 330 255 333 258 
rect 330 258 333 261 
rect 330 261 333 264 
rect 330 264 333 267 
rect 330 267 333 270 
rect 330 270 333 273 
rect 330 273 333 276 
rect 330 276 333 279 
rect 330 279 333 282 
rect 330 282 333 285 
rect 330 285 333 288 
rect 330 288 333 291 
rect 330 291 333 294 
rect 330 294 333 297 
rect 330 297 333 300 
rect 330 300 333 303 
rect 330 303 333 306 
rect 330 306 333 309 
rect 330 309 333 312 
rect 330 312 333 315 
rect 330 315 333 318 
rect 330 318 333 321 
rect 330 321 333 324 
rect 330 324 333 327 
rect 330 327 333 330 
rect 330 330 333 333 
rect 330 333 333 336 
rect 330 336 333 339 
rect 330 339 333 342 
rect 330 342 333 345 
rect 330 345 333 348 
rect 330 348 333 351 
rect 330 351 333 354 
rect 330 354 333 357 
rect 330 357 333 360 
rect 330 360 333 363 
rect 330 363 333 366 
rect 330 366 333 369 
rect 330 369 333 372 
rect 330 372 333 375 
rect 330 375 333 378 
rect 330 378 333 381 
rect 330 381 333 384 
rect 330 384 333 387 
rect 330 387 333 390 
rect 330 390 333 393 
rect 330 393 333 396 
rect 330 396 333 399 
rect 330 399 333 402 
rect 330 402 333 405 
rect 330 405 333 408 
rect 330 408 333 411 
rect 330 411 333 414 
rect 330 414 333 417 
rect 330 417 333 420 
rect 330 420 333 423 
rect 330 423 333 426 
rect 330 426 333 429 
rect 330 429 333 432 
rect 330 432 333 435 
rect 330 435 333 438 
rect 330 438 333 441 
rect 330 441 333 444 
rect 330 444 333 447 
rect 330 447 333 450 
rect 330 450 333 453 
rect 330 453 333 456 
rect 330 456 333 459 
rect 330 459 333 462 
rect 330 462 333 465 
rect 330 465 333 468 
rect 330 468 333 471 
rect 330 471 333 474 
rect 330 474 333 477 
rect 330 477 333 480 
rect 330 480 333 483 
rect 330 483 333 486 
rect 330 486 333 489 
rect 330 489 333 492 
rect 330 492 333 495 
rect 330 495 333 498 
rect 330 498 333 501 
rect 330 501 333 504 
rect 330 504 333 507 
rect 330 507 333 510 
rect 333 0 336 3 
rect 333 3 336 6 
rect 333 6 336 9 
rect 333 9 336 12 
rect 333 12 336 15 
rect 333 15 336 18 
rect 333 18 336 21 
rect 333 21 336 24 
rect 333 24 336 27 
rect 333 27 336 30 
rect 333 30 336 33 
rect 333 33 336 36 
rect 333 36 336 39 
rect 333 39 336 42 
rect 333 42 336 45 
rect 333 45 336 48 
rect 333 48 336 51 
rect 333 51 336 54 
rect 333 54 336 57 
rect 333 57 336 60 
rect 333 60 336 63 
rect 333 63 336 66 
rect 333 66 336 69 
rect 333 69 336 72 
rect 333 72 336 75 
rect 333 75 336 78 
rect 333 78 336 81 
rect 333 81 336 84 
rect 333 84 336 87 
rect 333 87 336 90 
rect 333 90 336 93 
rect 333 93 336 96 
rect 333 96 336 99 
rect 333 99 336 102 
rect 333 102 336 105 
rect 333 105 336 108 
rect 333 108 336 111 
rect 333 111 336 114 
rect 333 114 336 117 
rect 333 117 336 120 
rect 333 120 336 123 
rect 333 123 336 126 
rect 333 126 336 129 
rect 333 129 336 132 
rect 333 132 336 135 
rect 333 135 336 138 
rect 333 138 336 141 
rect 333 141 336 144 
rect 333 144 336 147 
rect 333 147 336 150 
rect 333 150 336 153 
rect 333 153 336 156 
rect 333 156 336 159 
rect 333 159 336 162 
rect 333 162 336 165 
rect 333 165 336 168 
rect 333 168 336 171 
rect 333 171 336 174 
rect 333 174 336 177 
rect 333 177 336 180 
rect 333 180 336 183 
rect 333 183 336 186 
rect 333 186 336 189 
rect 333 189 336 192 
rect 333 192 336 195 
rect 333 195 336 198 
rect 333 198 336 201 
rect 333 201 336 204 
rect 333 204 336 207 
rect 333 207 336 210 
rect 333 210 336 213 
rect 333 213 336 216 
rect 333 216 336 219 
rect 333 219 336 222 
rect 333 222 336 225 
rect 333 225 336 228 
rect 333 228 336 231 
rect 333 231 336 234 
rect 333 234 336 237 
rect 333 237 336 240 
rect 333 240 336 243 
rect 333 243 336 246 
rect 333 246 336 249 
rect 333 249 336 252 
rect 333 252 336 255 
rect 333 255 336 258 
rect 333 258 336 261 
rect 333 261 336 264 
rect 333 264 336 267 
rect 333 267 336 270 
rect 333 270 336 273 
rect 333 273 336 276 
rect 333 276 336 279 
rect 333 279 336 282 
rect 333 282 336 285 
rect 333 285 336 288 
rect 333 288 336 291 
rect 333 291 336 294 
rect 333 294 336 297 
rect 333 297 336 300 
rect 333 300 336 303 
rect 333 303 336 306 
rect 333 306 336 309 
rect 333 309 336 312 
rect 333 312 336 315 
rect 333 315 336 318 
rect 333 318 336 321 
rect 333 321 336 324 
rect 333 324 336 327 
rect 333 327 336 330 
rect 333 330 336 333 
rect 333 333 336 336 
rect 333 336 336 339 
rect 333 339 336 342 
rect 333 342 336 345 
rect 333 345 336 348 
rect 333 348 336 351 
rect 333 351 336 354 
rect 333 354 336 357 
rect 333 357 336 360 
rect 333 360 336 363 
rect 333 363 336 366 
rect 333 366 336 369 
rect 333 369 336 372 
rect 333 372 336 375 
rect 333 375 336 378 
rect 333 378 336 381 
rect 333 381 336 384 
rect 333 384 336 387 
rect 333 387 336 390 
rect 333 390 336 393 
rect 333 393 336 396 
rect 333 396 336 399 
rect 333 399 336 402 
rect 333 402 336 405 
rect 333 405 336 408 
rect 333 408 336 411 
rect 333 411 336 414 
rect 333 414 336 417 
rect 333 417 336 420 
rect 333 420 336 423 
rect 333 423 336 426 
rect 333 426 336 429 
rect 333 429 336 432 
rect 333 432 336 435 
rect 333 435 336 438 
rect 333 438 336 441 
rect 333 441 336 444 
rect 333 444 336 447 
rect 333 447 336 450 
rect 333 450 336 453 
rect 333 453 336 456 
rect 333 456 336 459 
rect 333 459 336 462 
rect 333 462 336 465 
rect 333 465 336 468 
rect 333 468 336 471 
rect 333 471 336 474 
rect 333 474 336 477 
rect 333 477 336 480 
rect 333 480 336 483 
rect 333 483 336 486 
rect 333 486 336 489 
rect 333 489 336 492 
rect 333 492 336 495 
rect 333 495 336 498 
rect 333 498 336 501 
rect 333 501 336 504 
rect 333 504 336 507 
rect 333 507 336 510 
rect 336 0 339 3 
rect 336 3 339 6 
rect 336 6 339 9 
rect 336 9 339 12 
rect 336 12 339 15 
rect 336 15 339 18 
rect 336 18 339 21 
rect 336 21 339 24 
rect 336 24 339 27 
rect 336 27 339 30 
rect 336 30 339 33 
rect 336 33 339 36 
rect 336 36 339 39 
rect 336 39 339 42 
rect 336 42 339 45 
rect 336 45 339 48 
rect 336 48 339 51 
rect 336 51 339 54 
rect 336 54 339 57 
rect 336 57 339 60 
rect 336 60 339 63 
rect 336 63 339 66 
rect 336 66 339 69 
rect 336 69 339 72 
rect 336 72 339 75 
rect 336 75 339 78 
rect 336 78 339 81 
rect 336 81 339 84 
rect 336 84 339 87 
rect 336 87 339 90 
rect 336 90 339 93 
rect 336 93 339 96 
rect 336 96 339 99 
rect 336 99 339 102 
rect 336 102 339 105 
rect 336 105 339 108 
rect 336 108 339 111 
rect 336 111 339 114 
rect 336 114 339 117 
rect 336 117 339 120 
rect 336 120 339 123 
rect 336 123 339 126 
rect 336 126 339 129 
rect 336 129 339 132 
rect 336 132 339 135 
rect 336 135 339 138 
rect 336 138 339 141 
rect 336 141 339 144 
rect 336 144 339 147 
rect 336 147 339 150 
rect 336 150 339 153 
rect 336 153 339 156 
rect 336 156 339 159 
rect 336 159 339 162 
rect 336 162 339 165 
rect 336 165 339 168 
rect 336 168 339 171 
rect 336 171 339 174 
rect 336 174 339 177 
rect 336 177 339 180 
rect 336 180 339 183 
rect 336 183 339 186 
rect 336 186 339 189 
rect 336 189 339 192 
rect 336 192 339 195 
rect 336 195 339 198 
rect 336 198 339 201 
rect 336 201 339 204 
rect 336 204 339 207 
rect 336 207 339 210 
rect 336 210 339 213 
rect 336 213 339 216 
rect 336 216 339 219 
rect 336 219 339 222 
rect 336 222 339 225 
rect 336 225 339 228 
rect 336 228 339 231 
rect 336 231 339 234 
rect 336 234 339 237 
rect 336 237 339 240 
rect 336 240 339 243 
rect 336 243 339 246 
rect 336 246 339 249 
rect 336 249 339 252 
rect 336 252 339 255 
rect 336 255 339 258 
rect 336 258 339 261 
rect 336 261 339 264 
rect 336 264 339 267 
rect 336 267 339 270 
rect 336 270 339 273 
rect 336 273 339 276 
rect 336 276 339 279 
rect 336 279 339 282 
rect 336 282 339 285 
rect 336 285 339 288 
rect 336 288 339 291 
rect 336 291 339 294 
rect 336 294 339 297 
rect 336 297 339 300 
rect 336 300 339 303 
rect 336 303 339 306 
rect 336 306 339 309 
rect 336 309 339 312 
rect 336 312 339 315 
rect 336 315 339 318 
rect 336 318 339 321 
rect 336 321 339 324 
rect 336 324 339 327 
rect 336 327 339 330 
rect 336 330 339 333 
rect 336 333 339 336 
rect 336 336 339 339 
rect 336 339 339 342 
rect 336 342 339 345 
rect 336 345 339 348 
rect 336 348 339 351 
rect 336 351 339 354 
rect 336 354 339 357 
rect 336 357 339 360 
rect 336 360 339 363 
rect 336 363 339 366 
rect 336 366 339 369 
rect 336 369 339 372 
rect 336 372 339 375 
rect 336 375 339 378 
rect 336 378 339 381 
rect 336 381 339 384 
rect 336 384 339 387 
rect 336 387 339 390 
rect 336 390 339 393 
rect 336 393 339 396 
rect 336 396 339 399 
rect 336 399 339 402 
rect 336 402 339 405 
rect 336 405 339 408 
rect 336 408 339 411 
rect 336 411 339 414 
rect 336 414 339 417 
rect 336 417 339 420 
rect 336 420 339 423 
rect 336 423 339 426 
rect 336 426 339 429 
rect 336 429 339 432 
rect 336 432 339 435 
rect 336 435 339 438 
rect 336 438 339 441 
rect 336 441 339 444 
rect 336 444 339 447 
rect 336 447 339 450 
rect 336 450 339 453 
rect 336 453 339 456 
rect 336 456 339 459 
rect 336 459 339 462 
rect 336 462 339 465 
rect 336 465 339 468 
rect 336 468 339 471 
rect 336 471 339 474 
rect 336 474 339 477 
rect 336 477 339 480 
rect 336 480 339 483 
rect 336 483 339 486 
rect 336 486 339 489 
rect 336 489 339 492 
rect 336 492 339 495 
rect 336 495 339 498 
rect 336 498 339 501 
rect 336 501 339 504 
rect 336 504 339 507 
rect 336 507 339 510 
rect 339 0 342 3 
rect 339 3 342 6 
rect 339 6 342 9 
rect 339 9 342 12 
rect 339 12 342 15 
rect 339 15 342 18 
rect 339 18 342 21 
rect 339 21 342 24 
rect 339 24 342 27 
rect 339 27 342 30 
rect 339 30 342 33 
rect 339 33 342 36 
rect 339 36 342 39 
rect 339 39 342 42 
rect 339 42 342 45 
rect 339 45 342 48 
rect 339 48 342 51 
rect 339 51 342 54 
rect 339 54 342 57 
rect 339 57 342 60 
rect 339 60 342 63 
rect 339 63 342 66 
rect 339 66 342 69 
rect 339 69 342 72 
rect 339 72 342 75 
rect 339 75 342 78 
rect 339 78 342 81 
rect 339 81 342 84 
rect 339 84 342 87 
rect 339 87 342 90 
rect 339 90 342 93 
rect 339 93 342 96 
rect 339 96 342 99 
rect 339 99 342 102 
rect 339 102 342 105 
rect 339 105 342 108 
rect 339 108 342 111 
rect 339 111 342 114 
rect 339 114 342 117 
rect 339 117 342 120 
rect 339 120 342 123 
rect 339 123 342 126 
rect 339 126 342 129 
rect 339 129 342 132 
rect 339 132 342 135 
rect 339 135 342 138 
rect 339 138 342 141 
rect 339 141 342 144 
rect 339 144 342 147 
rect 339 147 342 150 
rect 339 150 342 153 
rect 339 153 342 156 
rect 339 156 342 159 
rect 339 159 342 162 
rect 339 162 342 165 
rect 339 165 342 168 
rect 339 168 342 171 
rect 339 171 342 174 
rect 339 174 342 177 
rect 339 177 342 180 
rect 339 180 342 183 
rect 339 183 342 186 
rect 339 186 342 189 
rect 339 189 342 192 
rect 339 192 342 195 
rect 339 195 342 198 
rect 339 198 342 201 
rect 339 201 342 204 
rect 339 204 342 207 
rect 339 207 342 210 
rect 339 210 342 213 
rect 339 213 342 216 
rect 339 216 342 219 
rect 339 219 342 222 
rect 339 222 342 225 
rect 339 225 342 228 
rect 339 228 342 231 
rect 339 231 342 234 
rect 339 234 342 237 
rect 339 237 342 240 
rect 339 240 342 243 
rect 339 243 342 246 
rect 339 246 342 249 
rect 339 249 342 252 
rect 339 252 342 255 
rect 339 255 342 258 
rect 339 258 342 261 
rect 339 261 342 264 
rect 339 264 342 267 
rect 339 267 342 270 
rect 339 270 342 273 
rect 339 273 342 276 
rect 339 276 342 279 
rect 339 279 342 282 
rect 339 282 342 285 
rect 339 285 342 288 
rect 339 288 342 291 
rect 339 291 342 294 
rect 339 294 342 297 
rect 339 297 342 300 
rect 339 300 342 303 
rect 339 303 342 306 
rect 339 306 342 309 
rect 339 309 342 312 
rect 339 312 342 315 
rect 339 315 342 318 
rect 339 318 342 321 
rect 339 321 342 324 
rect 339 324 342 327 
rect 339 327 342 330 
rect 339 330 342 333 
rect 339 333 342 336 
rect 339 336 342 339 
rect 339 339 342 342 
rect 339 342 342 345 
rect 339 345 342 348 
rect 339 348 342 351 
rect 339 351 342 354 
rect 339 354 342 357 
rect 339 357 342 360 
rect 339 360 342 363 
rect 339 363 342 366 
rect 339 366 342 369 
rect 339 369 342 372 
rect 339 372 342 375 
rect 339 375 342 378 
rect 339 378 342 381 
rect 339 381 342 384 
rect 339 384 342 387 
rect 339 387 342 390 
rect 339 390 342 393 
rect 339 393 342 396 
rect 339 396 342 399 
rect 339 399 342 402 
rect 339 402 342 405 
rect 339 405 342 408 
rect 339 408 342 411 
rect 339 411 342 414 
rect 339 414 342 417 
rect 339 417 342 420 
rect 339 420 342 423 
rect 339 423 342 426 
rect 339 426 342 429 
rect 339 429 342 432 
rect 339 432 342 435 
rect 339 435 342 438 
rect 339 438 342 441 
rect 339 441 342 444 
rect 339 444 342 447 
rect 339 447 342 450 
rect 339 450 342 453 
rect 339 453 342 456 
rect 339 456 342 459 
rect 339 459 342 462 
rect 339 462 342 465 
rect 339 465 342 468 
rect 339 468 342 471 
rect 339 471 342 474 
rect 339 474 342 477 
rect 339 477 342 480 
rect 339 480 342 483 
rect 339 483 342 486 
rect 339 486 342 489 
rect 339 489 342 492 
rect 339 492 342 495 
rect 339 495 342 498 
rect 339 498 342 501 
rect 339 501 342 504 
rect 339 504 342 507 
rect 339 507 342 510 
rect 342 0 345 3 
rect 342 3 345 6 
rect 342 6 345 9 
rect 342 9 345 12 
rect 342 12 345 15 
rect 342 15 345 18 
rect 342 18 345 21 
rect 342 21 345 24 
rect 342 24 345 27 
rect 342 27 345 30 
rect 342 30 345 33 
rect 342 33 345 36 
rect 342 36 345 39 
rect 342 39 345 42 
rect 342 42 345 45 
rect 342 45 345 48 
rect 342 48 345 51 
rect 342 51 345 54 
rect 342 54 345 57 
rect 342 57 345 60 
rect 342 60 345 63 
rect 342 63 345 66 
rect 342 66 345 69 
rect 342 69 345 72 
rect 342 72 345 75 
rect 342 75 345 78 
rect 342 78 345 81 
rect 342 81 345 84 
rect 342 84 345 87 
rect 342 87 345 90 
rect 342 90 345 93 
rect 342 93 345 96 
rect 342 96 345 99 
rect 342 99 345 102 
rect 342 102 345 105 
rect 342 105 345 108 
rect 342 108 345 111 
rect 342 111 345 114 
rect 342 114 345 117 
rect 342 117 345 120 
rect 342 120 345 123 
rect 342 123 345 126 
rect 342 126 345 129 
rect 342 129 345 132 
rect 342 132 345 135 
rect 342 135 345 138 
rect 342 138 345 141 
rect 342 141 345 144 
rect 342 144 345 147 
rect 342 147 345 150 
rect 342 150 345 153 
rect 342 153 345 156 
rect 342 156 345 159 
rect 342 159 345 162 
rect 342 162 345 165 
rect 342 165 345 168 
rect 342 168 345 171 
rect 342 171 345 174 
rect 342 174 345 177 
rect 342 177 345 180 
rect 342 180 345 183 
rect 342 183 345 186 
rect 342 186 345 189 
rect 342 189 345 192 
rect 342 192 345 195 
rect 342 195 345 198 
rect 342 198 345 201 
rect 342 201 345 204 
rect 342 204 345 207 
rect 342 207 345 210 
rect 342 210 345 213 
rect 342 213 345 216 
rect 342 216 345 219 
rect 342 219 345 222 
rect 342 222 345 225 
rect 342 225 345 228 
rect 342 228 345 231 
rect 342 231 345 234 
rect 342 234 345 237 
rect 342 237 345 240 
rect 342 240 345 243 
rect 342 243 345 246 
rect 342 246 345 249 
rect 342 249 345 252 
rect 342 252 345 255 
rect 342 255 345 258 
rect 342 258 345 261 
rect 342 261 345 264 
rect 342 264 345 267 
rect 342 267 345 270 
rect 342 270 345 273 
rect 342 273 345 276 
rect 342 276 345 279 
rect 342 279 345 282 
rect 342 282 345 285 
rect 342 285 345 288 
rect 342 288 345 291 
rect 342 291 345 294 
rect 342 294 345 297 
rect 342 297 345 300 
rect 342 300 345 303 
rect 342 303 345 306 
rect 342 306 345 309 
rect 342 309 345 312 
rect 342 312 345 315 
rect 342 315 345 318 
rect 342 318 345 321 
rect 342 321 345 324 
rect 342 324 345 327 
rect 342 327 345 330 
rect 342 330 345 333 
rect 342 333 345 336 
rect 342 336 345 339 
rect 342 339 345 342 
rect 342 342 345 345 
rect 342 345 345 348 
rect 342 348 345 351 
rect 342 351 345 354 
rect 342 354 345 357 
rect 342 357 345 360 
rect 342 360 345 363 
rect 342 363 345 366 
rect 342 366 345 369 
rect 342 369 345 372 
rect 342 372 345 375 
rect 342 375 345 378 
rect 342 378 345 381 
rect 342 381 345 384 
rect 342 384 345 387 
rect 342 387 345 390 
rect 342 390 345 393 
rect 342 393 345 396 
rect 342 396 345 399 
rect 342 399 345 402 
rect 342 402 345 405 
rect 342 405 345 408 
rect 342 408 345 411 
rect 342 411 345 414 
rect 342 414 345 417 
rect 342 417 345 420 
rect 342 420 345 423 
rect 342 423 345 426 
rect 342 426 345 429 
rect 342 429 345 432 
rect 342 432 345 435 
rect 342 435 345 438 
rect 342 438 345 441 
rect 342 441 345 444 
rect 342 444 345 447 
rect 342 447 345 450 
rect 342 450 345 453 
rect 342 453 345 456 
rect 342 456 345 459 
rect 342 459 345 462 
rect 342 462 345 465 
rect 342 465 345 468 
rect 342 468 345 471 
rect 342 471 345 474 
rect 342 474 345 477 
rect 342 477 345 480 
rect 342 480 345 483 
rect 342 483 345 486 
rect 342 486 345 489 
rect 342 489 345 492 
rect 342 492 345 495 
rect 342 495 345 498 
rect 342 498 345 501 
rect 342 501 345 504 
rect 342 504 345 507 
rect 342 507 345 510 
rect 345 0 348 3 
rect 345 3 348 6 
rect 345 6 348 9 
rect 345 9 348 12 
rect 345 12 348 15 
rect 345 15 348 18 
rect 345 18 348 21 
rect 345 21 348 24 
rect 345 24 348 27 
rect 345 27 348 30 
rect 345 30 348 33 
rect 345 33 348 36 
rect 345 36 348 39 
rect 345 39 348 42 
rect 345 42 348 45 
rect 345 45 348 48 
rect 345 48 348 51 
rect 345 51 348 54 
rect 345 54 348 57 
rect 345 57 348 60 
rect 345 60 348 63 
rect 345 63 348 66 
rect 345 66 348 69 
rect 345 69 348 72 
rect 345 72 348 75 
rect 345 75 348 78 
rect 345 78 348 81 
rect 345 81 348 84 
rect 345 84 348 87 
rect 345 87 348 90 
rect 345 90 348 93 
rect 345 93 348 96 
rect 345 96 348 99 
rect 345 99 348 102 
rect 345 102 348 105 
rect 345 105 348 108 
rect 345 108 348 111 
rect 345 111 348 114 
rect 345 114 348 117 
rect 345 117 348 120 
rect 345 120 348 123 
rect 345 123 348 126 
rect 345 126 348 129 
rect 345 129 348 132 
rect 345 132 348 135 
rect 345 135 348 138 
rect 345 138 348 141 
rect 345 141 348 144 
rect 345 144 348 147 
rect 345 147 348 150 
rect 345 150 348 153 
rect 345 153 348 156 
rect 345 156 348 159 
rect 345 159 348 162 
rect 345 162 348 165 
rect 345 165 348 168 
rect 345 168 348 171 
rect 345 171 348 174 
rect 345 174 348 177 
rect 345 177 348 180 
rect 345 180 348 183 
rect 345 183 348 186 
rect 345 186 348 189 
rect 345 189 348 192 
rect 345 192 348 195 
rect 345 195 348 198 
rect 345 198 348 201 
rect 345 201 348 204 
rect 345 204 348 207 
rect 345 207 348 210 
rect 345 210 348 213 
rect 345 213 348 216 
rect 345 216 348 219 
rect 345 219 348 222 
rect 345 222 348 225 
rect 345 225 348 228 
rect 345 228 348 231 
rect 345 231 348 234 
rect 345 234 348 237 
rect 345 237 348 240 
rect 345 240 348 243 
rect 345 243 348 246 
rect 345 246 348 249 
rect 345 249 348 252 
rect 345 252 348 255 
rect 345 255 348 258 
rect 345 258 348 261 
rect 345 261 348 264 
rect 345 264 348 267 
rect 345 267 348 270 
rect 345 270 348 273 
rect 345 273 348 276 
rect 345 276 348 279 
rect 345 279 348 282 
rect 345 282 348 285 
rect 345 285 348 288 
rect 345 288 348 291 
rect 345 291 348 294 
rect 345 294 348 297 
rect 345 297 348 300 
rect 345 300 348 303 
rect 345 303 348 306 
rect 345 306 348 309 
rect 345 309 348 312 
rect 345 312 348 315 
rect 345 315 348 318 
rect 345 318 348 321 
rect 345 321 348 324 
rect 345 324 348 327 
rect 345 327 348 330 
rect 345 330 348 333 
rect 345 333 348 336 
rect 345 336 348 339 
rect 345 339 348 342 
rect 345 342 348 345 
rect 345 345 348 348 
rect 345 348 348 351 
rect 345 351 348 354 
rect 345 354 348 357 
rect 345 357 348 360 
rect 345 360 348 363 
rect 345 363 348 366 
rect 345 366 348 369 
rect 345 369 348 372 
rect 345 372 348 375 
rect 345 375 348 378 
rect 345 378 348 381 
rect 345 381 348 384 
rect 345 384 348 387 
rect 345 387 348 390 
rect 345 390 348 393 
rect 345 393 348 396 
rect 345 396 348 399 
rect 345 399 348 402 
rect 345 402 348 405 
rect 345 405 348 408 
rect 345 408 348 411 
rect 345 411 348 414 
rect 345 414 348 417 
rect 345 417 348 420 
rect 345 420 348 423 
rect 345 423 348 426 
rect 345 426 348 429 
rect 345 429 348 432 
rect 345 432 348 435 
rect 345 435 348 438 
rect 345 438 348 441 
rect 345 441 348 444 
rect 345 444 348 447 
rect 345 447 348 450 
rect 345 450 348 453 
rect 345 453 348 456 
rect 345 456 348 459 
rect 345 459 348 462 
rect 345 462 348 465 
rect 345 465 348 468 
rect 345 468 348 471 
rect 345 471 348 474 
rect 345 474 348 477 
rect 345 477 348 480 
rect 345 480 348 483 
rect 345 483 348 486 
rect 345 486 348 489 
rect 345 489 348 492 
rect 345 492 348 495 
rect 345 495 348 498 
rect 345 498 348 501 
rect 345 501 348 504 
rect 345 504 348 507 
rect 345 507 348 510 
rect 348 0 351 3 
rect 348 3 351 6 
rect 348 6 351 9 
rect 348 9 351 12 
rect 348 12 351 15 
rect 348 15 351 18 
rect 348 18 351 21 
rect 348 21 351 24 
rect 348 24 351 27 
rect 348 27 351 30 
rect 348 30 351 33 
rect 348 33 351 36 
rect 348 36 351 39 
rect 348 39 351 42 
rect 348 42 351 45 
rect 348 45 351 48 
rect 348 48 351 51 
rect 348 51 351 54 
rect 348 54 351 57 
rect 348 57 351 60 
rect 348 60 351 63 
rect 348 63 351 66 
rect 348 66 351 69 
rect 348 69 351 72 
rect 348 72 351 75 
rect 348 75 351 78 
rect 348 78 351 81 
rect 348 81 351 84 
rect 348 84 351 87 
rect 348 87 351 90 
rect 348 90 351 93 
rect 348 93 351 96 
rect 348 96 351 99 
rect 348 99 351 102 
rect 348 102 351 105 
rect 348 105 351 108 
rect 348 108 351 111 
rect 348 111 351 114 
rect 348 114 351 117 
rect 348 117 351 120 
rect 348 120 351 123 
rect 348 123 351 126 
rect 348 126 351 129 
rect 348 129 351 132 
rect 348 132 351 135 
rect 348 135 351 138 
rect 348 138 351 141 
rect 348 141 351 144 
rect 348 144 351 147 
rect 348 147 351 150 
rect 348 150 351 153 
rect 348 153 351 156 
rect 348 156 351 159 
rect 348 159 351 162 
rect 348 162 351 165 
rect 348 165 351 168 
rect 348 168 351 171 
rect 348 171 351 174 
rect 348 174 351 177 
rect 348 177 351 180 
rect 348 180 351 183 
rect 348 183 351 186 
rect 348 186 351 189 
rect 348 189 351 192 
rect 348 192 351 195 
rect 348 195 351 198 
rect 348 198 351 201 
rect 348 201 351 204 
rect 348 204 351 207 
rect 348 207 351 210 
rect 348 210 351 213 
rect 348 213 351 216 
rect 348 216 351 219 
rect 348 219 351 222 
rect 348 222 351 225 
rect 348 225 351 228 
rect 348 228 351 231 
rect 348 231 351 234 
rect 348 234 351 237 
rect 348 237 351 240 
rect 348 240 351 243 
rect 348 243 351 246 
rect 348 246 351 249 
rect 348 249 351 252 
rect 348 252 351 255 
rect 348 255 351 258 
rect 348 258 351 261 
rect 348 261 351 264 
rect 348 264 351 267 
rect 348 267 351 270 
rect 348 270 351 273 
rect 348 273 351 276 
rect 348 276 351 279 
rect 348 279 351 282 
rect 348 282 351 285 
rect 348 285 351 288 
rect 348 288 351 291 
rect 348 291 351 294 
rect 348 294 351 297 
rect 348 297 351 300 
rect 348 300 351 303 
rect 348 303 351 306 
rect 348 306 351 309 
rect 348 309 351 312 
rect 348 312 351 315 
rect 348 315 351 318 
rect 348 318 351 321 
rect 348 321 351 324 
rect 348 324 351 327 
rect 348 327 351 330 
rect 348 330 351 333 
rect 348 333 351 336 
rect 348 336 351 339 
rect 348 339 351 342 
rect 348 342 351 345 
rect 348 345 351 348 
rect 348 348 351 351 
rect 348 351 351 354 
rect 348 354 351 357 
rect 348 357 351 360 
rect 348 360 351 363 
rect 348 363 351 366 
rect 348 366 351 369 
rect 348 369 351 372 
rect 348 372 351 375 
rect 348 375 351 378 
rect 348 378 351 381 
rect 348 381 351 384 
rect 348 384 351 387 
rect 348 387 351 390 
rect 348 390 351 393 
rect 348 393 351 396 
rect 348 396 351 399 
rect 348 399 351 402 
rect 348 402 351 405 
rect 348 405 351 408 
rect 348 408 351 411 
rect 348 411 351 414 
rect 348 414 351 417 
rect 348 417 351 420 
rect 348 420 351 423 
rect 348 423 351 426 
rect 348 426 351 429 
rect 348 429 351 432 
rect 348 432 351 435 
rect 348 435 351 438 
rect 348 438 351 441 
rect 348 441 351 444 
rect 348 444 351 447 
rect 348 447 351 450 
rect 348 450 351 453 
rect 348 453 351 456 
rect 348 456 351 459 
rect 348 459 351 462 
rect 348 462 351 465 
rect 348 465 351 468 
rect 348 468 351 471 
rect 348 471 351 474 
rect 348 474 351 477 
rect 348 477 351 480 
rect 348 480 351 483 
rect 348 483 351 486 
rect 348 486 351 489 
rect 348 489 351 492 
rect 348 492 351 495 
rect 348 495 351 498 
rect 348 498 351 501 
rect 348 501 351 504 
rect 348 504 351 507 
rect 348 507 351 510 
rect 351 0 354 3 
rect 351 3 354 6 
rect 351 6 354 9 
rect 351 9 354 12 
rect 351 12 354 15 
rect 351 15 354 18 
rect 351 18 354 21 
rect 351 21 354 24 
rect 351 24 354 27 
rect 351 27 354 30 
rect 351 30 354 33 
rect 351 33 354 36 
rect 351 36 354 39 
rect 351 39 354 42 
rect 351 42 354 45 
rect 351 45 354 48 
rect 351 48 354 51 
rect 351 51 354 54 
rect 351 54 354 57 
rect 351 57 354 60 
rect 351 60 354 63 
rect 351 63 354 66 
rect 351 66 354 69 
rect 351 69 354 72 
rect 351 72 354 75 
rect 351 75 354 78 
rect 351 78 354 81 
rect 351 81 354 84 
rect 351 84 354 87 
rect 351 87 354 90 
rect 351 90 354 93 
rect 351 93 354 96 
rect 351 96 354 99 
rect 351 99 354 102 
rect 351 102 354 105 
rect 351 105 354 108 
rect 351 108 354 111 
rect 351 111 354 114 
rect 351 114 354 117 
rect 351 117 354 120 
rect 351 120 354 123 
rect 351 123 354 126 
rect 351 126 354 129 
rect 351 129 354 132 
rect 351 132 354 135 
rect 351 135 354 138 
rect 351 138 354 141 
rect 351 141 354 144 
rect 351 144 354 147 
rect 351 147 354 150 
rect 351 150 354 153 
rect 351 153 354 156 
rect 351 156 354 159 
rect 351 159 354 162 
rect 351 162 354 165 
rect 351 165 354 168 
rect 351 168 354 171 
rect 351 171 354 174 
rect 351 174 354 177 
rect 351 177 354 180 
rect 351 180 354 183 
rect 351 183 354 186 
rect 351 186 354 189 
rect 351 189 354 192 
rect 351 192 354 195 
rect 351 195 354 198 
rect 351 198 354 201 
rect 351 201 354 204 
rect 351 204 354 207 
rect 351 207 354 210 
rect 351 210 354 213 
rect 351 213 354 216 
rect 351 216 354 219 
rect 351 219 354 222 
rect 351 222 354 225 
rect 351 225 354 228 
rect 351 228 354 231 
rect 351 231 354 234 
rect 351 234 354 237 
rect 351 237 354 240 
rect 351 240 354 243 
rect 351 243 354 246 
rect 351 246 354 249 
rect 351 249 354 252 
rect 351 252 354 255 
rect 351 255 354 258 
rect 351 258 354 261 
rect 351 261 354 264 
rect 351 264 354 267 
rect 351 267 354 270 
rect 351 270 354 273 
rect 351 273 354 276 
rect 351 276 354 279 
rect 351 279 354 282 
rect 351 282 354 285 
rect 351 285 354 288 
rect 351 288 354 291 
rect 351 291 354 294 
rect 351 294 354 297 
rect 351 297 354 300 
rect 351 300 354 303 
rect 351 303 354 306 
rect 351 306 354 309 
rect 351 309 354 312 
rect 351 312 354 315 
rect 351 315 354 318 
rect 351 318 354 321 
rect 351 321 354 324 
rect 351 324 354 327 
rect 351 327 354 330 
rect 351 330 354 333 
rect 351 333 354 336 
rect 351 336 354 339 
rect 351 339 354 342 
rect 351 342 354 345 
rect 351 345 354 348 
rect 351 348 354 351 
rect 351 351 354 354 
rect 351 354 354 357 
rect 351 357 354 360 
rect 351 360 354 363 
rect 351 363 354 366 
rect 351 366 354 369 
rect 351 369 354 372 
rect 351 372 354 375 
rect 351 375 354 378 
rect 351 378 354 381 
rect 351 381 354 384 
rect 351 384 354 387 
rect 351 387 354 390 
rect 351 390 354 393 
rect 351 393 354 396 
rect 351 396 354 399 
rect 351 399 354 402 
rect 351 402 354 405 
rect 351 405 354 408 
rect 351 408 354 411 
rect 351 411 354 414 
rect 351 414 354 417 
rect 351 417 354 420 
rect 351 420 354 423 
rect 351 423 354 426 
rect 351 426 354 429 
rect 351 429 354 432 
rect 351 432 354 435 
rect 351 435 354 438 
rect 351 438 354 441 
rect 351 441 354 444 
rect 351 444 354 447 
rect 351 447 354 450 
rect 351 450 354 453 
rect 351 453 354 456 
rect 351 456 354 459 
rect 351 459 354 462 
rect 351 462 354 465 
rect 351 465 354 468 
rect 351 468 354 471 
rect 351 471 354 474 
rect 351 474 354 477 
rect 351 477 354 480 
rect 351 480 354 483 
rect 351 483 354 486 
rect 351 486 354 489 
rect 351 489 354 492 
rect 351 492 354 495 
rect 351 495 354 498 
rect 351 498 354 501 
rect 351 501 354 504 
rect 351 504 354 507 
rect 351 507 354 510 
rect 354 0 357 3 
rect 354 3 357 6 
rect 354 6 357 9 
rect 354 9 357 12 
rect 354 12 357 15 
rect 354 15 357 18 
rect 354 18 357 21 
rect 354 21 357 24 
rect 354 24 357 27 
rect 354 27 357 30 
rect 354 30 357 33 
rect 354 33 357 36 
rect 354 36 357 39 
rect 354 39 357 42 
rect 354 42 357 45 
rect 354 45 357 48 
rect 354 48 357 51 
rect 354 51 357 54 
rect 354 54 357 57 
rect 354 57 357 60 
rect 354 60 357 63 
rect 354 63 357 66 
rect 354 66 357 69 
rect 354 69 357 72 
rect 354 72 357 75 
rect 354 75 357 78 
rect 354 78 357 81 
rect 354 81 357 84 
rect 354 84 357 87 
rect 354 87 357 90 
rect 354 90 357 93 
rect 354 93 357 96 
rect 354 96 357 99 
rect 354 99 357 102 
rect 354 102 357 105 
rect 354 105 357 108 
rect 354 108 357 111 
rect 354 111 357 114 
rect 354 114 357 117 
rect 354 117 357 120 
rect 354 120 357 123 
rect 354 123 357 126 
rect 354 126 357 129 
rect 354 129 357 132 
rect 354 132 357 135 
rect 354 135 357 138 
rect 354 138 357 141 
rect 354 141 357 144 
rect 354 144 357 147 
rect 354 147 357 150 
rect 354 150 357 153 
rect 354 153 357 156 
rect 354 156 357 159 
rect 354 159 357 162 
rect 354 162 357 165 
rect 354 165 357 168 
rect 354 168 357 171 
rect 354 171 357 174 
rect 354 174 357 177 
rect 354 177 357 180 
rect 354 180 357 183 
rect 354 183 357 186 
rect 354 186 357 189 
rect 354 189 357 192 
rect 354 192 357 195 
rect 354 195 357 198 
rect 354 198 357 201 
rect 354 201 357 204 
rect 354 204 357 207 
rect 354 207 357 210 
rect 354 210 357 213 
rect 354 213 357 216 
rect 354 216 357 219 
rect 354 219 357 222 
rect 354 222 357 225 
rect 354 225 357 228 
rect 354 228 357 231 
rect 354 231 357 234 
rect 354 234 357 237 
rect 354 237 357 240 
rect 354 240 357 243 
rect 354 243 357 246 
rect 354 246 357 249 
rect 354 249 357 252 
rect 354 252 357 255 
rect 354 255 357 258 
rect 354 258 357 261 
rect 354 261 357 264 
rect 354 264 357 267 
rect 354 267 357 270 
rect 354 270 357 273 
rect 354 273 357 276 
rect 354 276 357 279 
rect 354 279 357 282 
rect 354 282 357 285 
rect 354 285 357 288 
rect 354 288 357 291 
rect 354 291 357 294 
rect 354 294 357 297 
rect 354 297 357 300 
rect 354 300 357 303 
rect 354 303 357 306 
rect 354 306 357 309 
rect 354 309 357 312 
rect 354 312 357 315 
rect 354 315 357 318 
rect 354 318 357 321 
rect 354 321 357 324 
rect 354 324 357 327 
rect 354 327 357 330 
rect 354 330 357 333 
rect 354 333 357 336 
rect 354 336 357 339 
rect 354 339 357 342 
rect 354 342 357 345 
rect 354 345 357 348 
rect 354 348 357 351 
rect 354 351 357 354 
rect 354 354 357 357 
rect 354 357 357 360 
rect 354 360 357 363 
rect 354 363 357 366 
rect 354 366 357 369 
rect 354 369 357 372 
rect 354 372 357 375 
rect 354 375 357 378 
rect 354 378 357 381 
rect 354 381 357 384 
rect 354 384 357 387 
rect 354 387 357 390 
rect 354 390 357 393 
rect 354 393 357 396 
rect 354 396 357 399 
rect 354 399 357 402 
rect 354 402 357 405 
rect 354 405 357 408 
rect 354 408 357 411 
rect 354 411 357 414 
rect 354 414 357 417 
rect 354 417 357 420 
rect 354 420 357 423 
rect 354 423 357 426 
rect 354 426 357 429 
rect 354 429 357 432 
rect 354 432 357 435 
rect 354 435 357 438 
rect 354 438 357 441 
rect 354 441 357 444 
rect 354 444 357 447 
rect 354 447 357 450 
rect 354 450 357 453 
rect 354 453 357 456 
rect 354 456 357 459 
rect 354 459 357 462 
rect 354 462 357 465 
rect 354 465 357 468 
rect 354 468 357 471 
rect 354 471 357 474 
rect 354 474 357 477 
rect 354 477 357 480 
rect 354 480 357 483 
rect 354 483 357 486 
rect 354 486 357 489 
rect 354 489 357 492 
rect 354 492 357 495 
rect 354 495 357 498 
rect 354 498 357 501 
rect 354 501 357 504 
rect 354 504 357 507 
rect 354 507 357 510 
rect 357 0 360 3 
rect 357 3 360 6 
rect 357 6 360 9 
rect 357 9 360 12 
rect 357 12 360 15 
rect 357 15 360 18 
rect 357 18 360 21 
rect 357 21 360 24 
rect 357 24 360 27 
rect 357 27 360 30 
rect 357 30 360 33 
rect 357 33 360 36 
rect 357 36 360 39 
rect 357 39 360 42 
rect 357 42 360 45 
rect 357 45 360 48 
rect 357 48 360 51 
rect 357 51 360 54 
rect 357 54 360 57 
rect 357 57 360 60 
rect 357 60 360 63 
rect 357 63 360 66 
rect 357 66 360 69 
rect 357 69 360 72 
rect 357 72 360 75 
rect 357 75 360 78 
rect 357 78 360 81 
rect 357 81 360 84 
rect 357 84 360 87 
rect 357 87 360 90 
rect 357 90 360 93 
rect 357 93 360 96 
rect 357 96 360 99 
rect 357 99 360 102 
rect 357 102 360 105 
rect 357 105 360 108 
rect 357 108 360 111 
rect 357 111 360 114 
rect 357 114 360 117 
rect 357 117 360 120 
rect 357 120 360 123 
rect 357 123 360 126 
rect 357 126 360 129 
rect 357 129 360 132 
rect 357 132 360 135 
rect 357 135 360 138 
rect 357 138 360 141 
rect 357 141 360 144 
rect 357 144 360 147 
rect 357 147 360 150 
rect 357 150 360 153 
rect 357 153 360 156 
rect 357 156 360 159 
rect 357 159 360 162 
rect 357 162 360 165 
rect 357 165 360 168 
rect 357 168 360 171 
rect 357 171 360 174 
rect 357 174 360 177 
rect 357 177 360 180 
rect 357 180 360 183 
rect 357 183 360 186 
rect 357 186 360 189 
rect 357 189 360 192 
rect 357 192 360 195 
rect 357 195 360 198 
rect 357 198 360 201 
rect 357 201 360 204 
rect 357 204 360 207 
rect 357 207 360 210 
rect 357 210 360 213 
rect 357 213 360 216 
rect 357 216 360 219 
rect 357 219 360 222 
rect 357 222 360 225 
rect 357 225 360 228 
rect 357 228 360 231 
rect 357 231 360 234 
rect 357 234 360 237 
rect 357 237 360 240 
rect 357 240 360 243 
rect 357 243 360 246 
rect 357 246 360 249 
rect 357 249 360 252 
rect 357 252 360 255 
rect 357 255 360 258 
rect 357 258 360 261 
rect 357 261 360 264 
rect 357 264 360 267 
rect 357 267 360 270 
rect 357 270 360 273 
rect 357 273 360 276 
rect 357 276 360 279 
rect 357 279 360 282 
rect 357 282 360 285 
rect 357 285 360 288 
rect 357 288 360 291 
rect 357 291 360 294 
rect 357 294 360 297 
rect 357 297 360 300 
rect 357 300 360 303 
rect 357 303 360 306 
rect 357 306 360 309 
rect 357 309 360 312 
rect 357 312 360 315 
rect 357 315 360 318 
rect 357 318 360 321 
rect 357 321 360 324 
rect 357 324 360 327 
rect 357 327 360 330 
rect 357 330 360 333 
rect 357 333 360 336 
rect 357 336 360 339 
rect 357 339 360 342 
rect 357 342 360 345 
rect 357 345 360 348 
rect 357 348 360 351 
rect 357 351 360 354 
rect 357 354 360 357 
rect 357 357 360 360 
rect 357 360 360 363 
rect 357 363 360 366 
rect 357 366 360 369 
rect 357 369 360 372 
rect 357 372 360 375 
rect 357 375 360 378 
rect 357 378 360 381 
rect 357 381 360 384 
rect 357 384 360 387 
rect 357 387 360 390 
rect 357 390 360 393 
rect 357 393 360 396 
rect 357 396 360 399 
rect 357 399 360 402 
rect 357 402 360 405 
rect 357 405 360 408 
rect 357 408 360 411 
rect 357 411 360 414 
rect 357 414 360 417 
rect 357 417 360 420 
rect 357 420 360 423 
rect 357 423 360 426 
rect 357 426 360 429 
rect 357 429 360 432 
rect 357 432 360 435 
rect 357 435 360 438 
rect 357 438 360 441 
rect 357 441 360 444 
rect 357 444 360 447 
rect 357 447 360 450 
rect 357 450 360 453 
rect 357 453 360 456 
rect 357 456 360 459 
rect 357 459 360 462 
rect 357 462 360 465 
rect 357 465 360 468 
rect 357 468 360 471 
rect 357 471 360 474 
rect 357 474 360 477 
rect 357 477 360 480 
rect 357 480 360 483 
rect 357 483 360 486 
rect 357 486 360 489 
rect 357 489 360 492 
rect 357 492 360 495 
rect 357 495 360 498 
rect 357 498 360 501 
rect 357 501 360 504 
rect 357 504 360 507 
rect 357 507 360 510 
rect 360 0 363 3 
rect 360 3 363 6 
rect 360 6 363 9 
rect 360 9 363 12 
rect 360 12 363 15 
rect 360 15 363 18 
rect 360 18 363 21 
rect 360 21 363 24 
rect 360 24 363 27 
rect 360 27 363 30 
rect 360 30 363 33 
rect 360 33 363 36 
rect 360 36 363 39 
rect 360 39 363 42 
rect 360 42 363 45 
rect 360 45 363 48 
rect 360 48 363 51 
rect 360 51 363 54 
rect 360 54 363 57 
rect 360 57 363 60 
rect 360 60 363 63 
rect 360 63 363 66 
rect 360 66 363 69 
rect 360 69 363 72 
rect 360 72 363 75 
rect 360 75 363 78 
rect 360 78 363 81 
rect 360 81 363 84 
rect 360 84 363 87 
rect 360 87 363 90 
rect 360 90 363 93 
rect 360 93 363 96 
rect 360 96 363 99 
rect 360 99 363 102 
rect 360 102 363 105 
rect 360 105 363 108 
rect 360 108 363 111 
rect 360 111 363 114 
rect 360 114 363 117 
rect 360 117 363 120 
rect 360 120 363 123 
rect 360 123 363 126 
rect 360 126 363 129 
rect 360 129 363 132 
rect 360 132 363 135 
rect 360 135 363 138 
rect 360 138 363 141 
rect 360 141 363 144 
rect 360 144 363 147 
rect 360 147 363 150 
rect 360 150 363 153 
rect 360 153 363 156 
rect 360 156 363 159 
rect 360 159 363 162 
rect 360 162 363 165 
rect 360 165 363 168 
rect 360 168 363 171 
rect 360 171 363 174 
rect 360 174 363 177 
rect 360 177 363 180 
rect 360 180 363 183 
rect 360 183 363 186 
rect 360 186 363 189 
rect 360 189 363 192 
rect 360 192 363 195 
rect 360 195 363 198 
rect 360 198 363 201 
rect 360 201 363 204 
rect 360 204 363 207 
rect 360 207 363 210 
rect 360 210 363 213 
rect 360 213 363 216 
rect 360 216 363 219 
rect 360 219 363 222 
rect 360 222 363 225 
rect 360 225 363 228 
rect 360 228 363 231 
rect 360 231 363 234 
rect 360 234 363 237 
rect 360 237 363 240 
rect 360 240 363 243 
rect 360 243 363 246 
rect 360 246 363 249 
rect 360 249 363 252 
rect 360 252 363 255 
rect 360 255 363 258 
rect 360 258 363 261 
rect 360 261 363 264 
rect 360 264 363 267 
rect 360 267 363 270 
rect 360 270 363 273 
rect 360 273 363 276 
rect 360 276 363 279 
rect 360 279 363 282 
rect 360 282 363 285 
rect 360 285 363 288 
rect 360 288 363 291 
rect 360 291 363 294 
rect 360 294 363 297 
rect 360 297 363 300 
rect 360 300 363 303 
rect 360 303 363 306 
rect 360 306 363 309 
rect 360 309 363 312 
rect 360 312 363 315 
rect 360 315 363 318 
rect 360 318 363 321 
rect 360 321 363 324 
rect 360 324 363 327 
rect 360 327 363 330 
rect 360 330 363 333 
rect 360 333 363 336 
rect 360 336 363 339 
rect 360 339 363 342 
rect 360 342 363 345 
rect 360 345 363 348 
rect 360 348 363 351 
rect 360 351 363 354 
rect 360 354 363 357 
rect 360 357 363 360 
rect 360 360 363 363 
rect 360 363 363 366 
rect 360 366 363 369 
rect 360 369 363 372 
rect 360 372 363 375 
rect 360 375 363 378 
rect 360 378 363 381 
rect 360 381 363 384 
rect 360 384 363 387 
rect 360 387 363 390 
rect 360 390 363 393 
rect 360 393 363 396 
rect 360 396 363 399 
rect 360 399 363 402 
rect 360 402 363 405 
rect 360 405 363 408 
rect 360 408 363 411 
rect 360 411 363 414 
rect 360 414 363 417 
rect 360 417 363 420 
rect 360 420 363 423 
rect 360 423 363 426 
rect 360 426 363 429 
rect 360 429 363 432 
rect 360 432 363 435 
rect 360 435 363 438 
rect 360 438 363 441 
rect 360 441 363 444 
rect 360 444 363 447 
rect 360 447 363 450 
rect 360 450 363 453 
rect 360 453 363 456 
rect 360 456 363 459 
rect 360 459 363 462 
rect 360 462 363 465 
rect 360 465 363 468 
rect 360 468 363 471 
rect 360 471 363 474 
rect 360 474 363 477 
rect 360 477 363 480 
rect 360 480 363 483 
rect 360 483 363 486 
rect 360 486 363 489 
rect 360 489 363 492 
rect 360 492 363 495 
rect 360 495 363 498 
rect 360 498 363 501 
rect 360 501 363 504 
rect 360 504 363 507 
rect 360 507 363 510 
rect 363 0 366 3 
rect 363 3 366 6 
rect 363 6 366 9 
rect 363 9 366 12 
rect 363 12 366 15 
rect 363 15 366 18 
rect 363 18 366 21 
rect 363 21 366 24 
rect 363 24 366 27 
rect 363 27 366 30 
rect 363 30 366 33 
rect 363 33 366 36 
rect 363 36 366 39 
rect 363 39 366 42 
rect 363 42 366 45 
rect 363 45 366 48 
rect 363 48 366 51 
rect 363 51 366 54 
rect 363 54 366 57 
rect 363 57 366 60 
rect 363 60 366 63 
rect 363 63 366 66 
rect 363 66 366 69 
rect 363 69 366 72 
rect 363 72 366 75 
rect 363 75 366 78 
rect 363 78 366 81 
rect 363 81 366 84 
rect 363 84 366 87 
rect 363 87 366 90 
rect 363 90 366 93 
rect 363 93 366 96 
rect 363 96 366 99 
rect 363 99 366 102 
rect 363 102 366 105 
rect 363 105 366 108 
rect 363 108 366 111 
rect 363 111 366 114 
rect 363 114 366 117 
rect 363 117 366 120 
rect 363 120 366 123 
rect 363 123 366 126 
rect 363 126 366 129 
rect 363 129 366 132 
rect 363 132 366 135 
rect 363 135 366 138 
rect 363 138 366 141 
rect 363 141 366 144 
rect 363 144 366 147 
rect 363 147 366 150 
rect 363 150 366 153 
rect 363 153 366 156 
rect 363 156 366 159 
rect 363 159 366 162 
rect 363 162 366 165 
rect 363 165 366 168 
rect 363 168 366 171 
rect 363 171 366 174 
rect 363 174 366 177 
rect 363 177 366 180 
rect 363 180 366 183 
rect 363 183 366 186 
rect 363 186 366 189 
rect 363 189 366 192 
rect 363 192 366 195 
rect 363 195 366 198 
rect 363 198 366 201 
rect 363 201 366 204 
rect 363 204 366 207 
rect 363 207 366 210 
rect 363 210 366 213 
rect 363 213 366 216 
rect 363 216 366 219 
rect 363 219 366 222 
rect 363 222 366 225 
rect 363 225 366 228 
rect 363 228 366 231 
rect 363 231 366 234 
rect 363 234 366 237 
rect 363 237 366 240 
rect 363 240 366 243 
rect 363 243 366 246 
rect 363 246 366 249 
rect 363 249 366 252 
rect 363 252 366 255 
rect 363 255 366 258 
rect 363 258 366 261 
rect 363 261 366 264 
rect 363 264 366 267 
rect 363 267 366 270 
rect 363 270 366 273 
rect 363 273 366 276 
rect 363 276 366 279 
rect 363 279 366 282 
rect 363 282 366 285 
rect 363 285 366 288 
rect 363 288 366 291 
rect 363 291 366 294 
rect 363 294 366 297 
rect 363 297 366 300 
rect 363 300 366 303 
rect 363 303 366 306 
rect 363 306 366 309 
rect 363 309 366 312 
rect 363 312 366 315 
rect 363 315 366 318 
rect 363 318 366 321 
rect 363 321 366 324 
rect 363 324 366 327 
rect 363 327 366 330 
rect 363 330 366 333 
rect 363 333 366 336 
rect 363 336 366 339 
rect 363 339 366 342 
rect 363 342 366 345 
rect 363 345 366 348 
rect 363 348 366 351 
rect 363 351 366 354 
rect 363 354 366 357 
rect 363 357 366 360 
rect 363 360 366 363 
rect 363 363 366 366 
rect 363 366 366 369 
rect 363 369 366 372 
rect 363 372 366 375 
rect 363 375 366 378 
rect 363 378 366 381 
rect 363 381 366 384 
rect 363 384 366 387 
rect 363 387 366 390 
rect 363 390 366 393 
rect 363 393 366 396 
rect 363 396 366 399 
rect 363 399 366 402 
rect 363 402 366 405 
rect 363 405 366 408 
rect 363 408 366 411 
rect 363 411 366 414 
rect 363 414 366 417 
rect 363 417 366 420 
rect 363 420 366 423 
rect 363 423 366 426 
rect 363 426 366 429 
rect 363 429 366 432 
rect 363 432 366 435 
rect 363 435 366 438 
rect 363 438 366 441 
rect 363 441 366 444 
rect 363 444 366 447 
rect 363 447 366 450 
rect 363 450 366 453 
rect 363 453 366 456 
rect 363 456 366 459 
rect 363 459 366 462 
rect 363 462 366 465 
rect 363 465 366 468 
rect 363 468 366 471 
rect 363 471 366 474 
rect 363 474 366 477 
rect 363 477 366 480 
rect 363 480 366 483 
rect 363 483 366 486 
rect 363 486 366 489 
rect 363 489 366 492 
rect 363 492 366 495 
rect 363 495 366 498 
rect 363 498 366 501 
rect 363 501 366 504 
rect 363 504 366 507 
rect 363 507 366 510 
rect 366 0 369 3 
rect 366 3 369 6 
rect 366 6 369 9 
rect 366 9 369 12 
rect 366 12 369 15 
rect 366 15 369 18 
rect 366 18 369 21 
rect 366 21 369 24 
rect 366 24 369 27 
rect 366 27 369 30 
rect 366 30 369 33 
rect 366 33 369 36 
rect 366 36 369 39 
rect 366 39 369 42 
rect 366 42 369 45 
rect 366 45 369 48 
rect 366 48 369 51 
rect 366 51 369 54 
rect 366 54 369 57 
rect 366 57 369 60 
rect 366 60 369 63 
rect 366 63 369 66 
rect 366 66 369 69 
rect 366 69 369 72 
rect 366 72 369 75 
rect 366 75 369 78 
rect 366 78 369 81 
rect 366 81 369 84 
rect 366 84 369 87 
rect 366 87 369 90 
rect 366 90 369 93 
rect 366 93 369 96 
rect 366 96 369 99 
rect 366 99 369 102 
rect 366 102 369 105 
rect 366 105 369 108 
rect 366 108 369 111 
rect 366 111 369 114 
rect 366 114 369 117 
rect 366 117 369 120 
rect 366 120 369 123 
rect 366 123 369 126 
rect 366 126 369 129 
rect 366 129 369 132 
rect 366 132 369 135 
rect 366 135 369 138 
rect 366 138 369 141 
rect 366 141 369 144 
rect 366 144 369 147 
rect 366 147 369 150 
rect 366 150 369 153 
rect 366 153 369 156 
rect 366 156 369 159 
rect 366 159 369 162 
rect 366 162 369 165 
rect 366 165 369 168 
rect 366 168 369 171 
rect 366 171 369 174 
rect 366 174 369 177 
rect 366 177 369 180 
rect 366 180 369 183 
rect 366 183 369 186 
rect 366 186 369 189 
rect 366 189 369 192 
rect 366 192 369 195 
rect 366 195 369 198 
rect 366 198 369 201 
rect 366 201 369 204 
rect 366 204 369 207 
rect 366 207 369 210 
rect 366 210 369 213 
rect 366 213 369 216 
rect 366 216 369 219 
rect 366 219 369 222 
rect 366 222 369 225 
rect 366 225 369 228 
rect 366 228 369 231 
rect 366 231 369 234 
rect 366 234 369 237 
rect 366 237 369 240 
rect 366 240 369 243 
rect 366 243 369 246 
rect 366 246 369 249 
rect 366 249 369 252 
rect 366 252 369 255 
rect 366 255 369 258 
rect 366 258 369 261 
rect 366 261 369 264 
rect 366 264 369 267 
rect 366 267 369 270 
rect 366 270 369 273 
rect 366 273 369 276 
rect 366 276 369 279 
rect 366 279 369 282 
rect 366 282 369 285 
rect 366 285 369 288 
rect 366 288 369 291 
rect 366 291 369 294 
rect 366 294 369 297 
rect 366 297 369 300 
rect 366 300 369 303 
rect 366 303 369 306 
rect 366 306 369 309 
rect 366 309 369 312 
rect 366 312 369 315 
rect 366 315 369 318 
rect 366 318 369 321 
rect 366 321 369 324 
rect 366 324 369 327 
rect 366 327 369 330 
rect 366 330 369 333 
rect 366 333 369 336 
rect 366 336 369 339 
rect 366 339 369 342 
rect 366 342 369 345 
rect 366 345 369 348 
rect 366 348 369 351 
rect 366 351 369 354 
rect 366 354 369 357 
rect 366 357 369 360 
rect 366 360 369 363 
rect 366 363 369 366 
rect 366 366 369 369 
rect 366 369 369 372 
rect 366 372 369 375 
rect 366 375 369 378 
rect 366 378 369 381 
rect 366 381 369 384 
rect 366 384 369 387 
rect 366 387 369 390 
rect 366 390 369 393 
rect 366 393 369 396 
rect 366 396 369 399 
rect 366 399 369 402 
rect 366 402 369 405 
rect 366 405 369 408 
rect 366 408 369 411 
rect 366 411 369 414 
rect 366 414 369 417 
rect 366 417 369 420 
rect 366 420 369 423 
rect 366 423 369 426 
rect 366 426 369 429 
rect 366 429 369 432 
rect 366 432 369 435 
rect 366 435 369 438 
rect 366 438 369 441 
rect 366 441 369 444 
rect 366 444 369 447 
rect 366 447 369 450 
rect 366 450 369 453 
rect 366 453 369 456 
rect 366 456 369 459 
rect 366 459 369 462 
rect 366 462 369 465 
rect 366 465 369 468 
rect 366 468 369 471 
rect 366 471 369 474 
rect 366 474 369 477 
rect 366 477 369 480 
rect 366 480 369 483 
rect 366 483 369 486 
rect 366 486 369 489 
rect 366 489 369 492 
rect 366 492 369 495 
rect 366 495 369 498 
rect 366 498 369 501 
rect 366 501 369 504 
rect 366 504 369 507 
rect 366 507 369 510 
rect 369 0 372 3 
rect 369 3 372 6 
rect 369 6 372 9 
rect 369 9 372 12 
rect 369 12 372 15 
rect 369 15 372 18 
rect 369 18 372 21 
rect 369 21 372 24 
rect 369 24 372 27 
rect 369 27 372 30 
rect 369 30 372 33 
rect 369 33 372 36 
rect 369 36 372 39 
rect 369 39 372 42 
rect 369 42 372 45 
rect 369 45 372 48 
rect 369 48 372 51 
rect 369 51 372 54 
rect 369 54 372 57 
rect 369 57 372 60 
rect 369 60 372 63 
rect 369 63 372 66 
rect 369 66 372 69 
rect 369 69 372 72 
rect 369 72 372 75 
rect 369 75 372 78 
rect 369 78 372 81 
rect 369 81 372 84 
rect 369 84 372 87 
rect 369 87 372 90 
rect 369 90 372 93 
rect 369 93 372 96 
rect 369 96 372 99 
rect 369 99 372 102 
rect 369 102 372 105 
rect 369 105 372 108 
rect 369 108 372 111 
rect 369 111 372 114 
rect 369 114 372 117 
rect 369 117 372 120 
rect 369 120 372 123 
rect 369 123 372 126 
rect 369 126 372 129 
rect 369 129 372 132 
rect 369 132 372 135 
rect 369 135 372 138 
rect 369 138 372 141 
rect 369 141 372 144 
rect 369 144 372 147 
rect 369 147 372 150 
rect 369 150 372 153 
rect 369 153 372 156 
rect 369 156 372 159 
rect 369 159 372 162 
rect 369 162 372 165 
rect 369 165 372 168 
rect 369 168 372 171 
rect 369 171 372 174 
rect 369 174 372 177 
rect 369 177 372 180 
rect 369 180 372 183 
rect 369 183 372 186 
rect 369 186 372 189 
rect 369 189 372 192 
rect 369 192 372 195 
rect 369 195 372 198 
rect 369 198 372 201 
rect 369 201 372 204 
rect 369 204 372 207 
rect 369 207 372 210 
rect 369 210 372 213 
rect 369 213 372 216 
rect 369 216 372 219 
rect 369 219 372 222 
rect 369 222 372 225 
rect 369 225 372 228 
rect 369 228 372 231 
rect 369 231 372 234 
rect 369 234 372 237 
rect 369 237 372 240 
rect 369 240 372 243 
rect 369 243 372 246 
rect 369 246 372 249 
rect 369 249 372 252 
rect 369 252 372 255 
rect 369 255 372 258 
rect 369 258 372 261 
rect 369 261 372 264 
rect 369 264 372 267 
rect 369 267 372 270 
rect 369 270 372 273 
rect 369 273 372 276 
rect 369 276 372 279 
rect 369 279 372 282 
rect 369 282 372 285 
rect 369 285 372 288 
rect 369 288 372 291 
rect 369 291 372 294 
rect 369 294 372 297 
rect 369 297 372 300 
rect 369 300 372 303 
rect 369 303 372 306 
rect 369 306 372 309 
rect 369 309 372 312 
rect 369 312 372 315 
rect 369 315 372 318 
rect 369 318 372 321 
rect 369 321 372 324 
rect 369 324 372 327 
rect 369 327 372 330 
rect 369 330 372 333 
rect 369 333 372 336 
rect 369 336 372 339 
rect 369 339 372 342 
rect 369 342 372 345 
rect 369 345 372 348 
rect 369 348 372 351 
rect 369 351 372 354 
rect 369 354 372 357 
rect 369 357 372 360 
rect 369 360 372 363 
rect 369 363 372 366 
rect 369 366 372 369 
rect 369 369 372 372 
rect 369 372 372 375 
rect 369 375 372 378 
rect 369 378 372 381 
rect 369 381 372 384 
rect 369 384 372 387 
rect 369 387 372 390 
rect 369 390 372 393 
rect 369 393 372 396 
rect 369 396 372 399 
rect 369 399 372 402 
rect 369 402 372 405 
rect 369 405 372 408 
rect 369 408 372 411 
rect 369 411 372 414 
rect 369 414 372 417 
rect 369 417 372 420 
rect 369 420 372 423 
rect 369 423 372 426 
rect 369 426 372 429 
rect 369 429 372 432 
rect 369 432 372 435 
rect 369 435 372 438 
rect 369 438 372 441 
rect 369 441 372 444 
rect 369 444 372 447 
rect 369 447 372 450 
rect 369 450 372 453 
rect 369 453 372 456 
rect 369 456 372 459 
rect 369 459 372 462 
rect 369 462 372 465 
rect 369 465 372 468 
rect 369 468 372 471 
rect 369 471 372 474 
rect 369 474 372 477 
rect 369 477 372 480 
rect 369 480 372 483 
rect 369 483 372 486 
rect 369 486 372 489 
rect 369 489 372 492 
rect 369 492 372 495 
rect 369 495 372 498 
rect 369 498 372 501 
rect 369 501 372 504 
rect 369 504 372 507 
rect 369 507 372 510 
rect 372 0 375 3 
rect 372 3 375 6 
rect 372 6 375 9 
rect 372 9 375 12 
rect 372 12 375 15 
rect 372 15 375 18 
rect 372 18 375 21 
rect 372 21 375 24 
rect 372 24 375 27 
rect 372 27 375 30 
rect 372 30 375 33 
rect 372 33 375 36 
rect 372 36 375 39 
rect 372 39 375 42 
rect 372 42 375 45 
rect 372 45 375 48 
rect 372 48 375 51 
rect 372 51 375 54 
rect 372 54 375 57 
rect 372 57 375 60 
rect 372 60 375 63 
rect 372 63 375 66 
rect 372 66 375 69 
rect 372 69 375 72 
rect 372 72 375 75 
rect 372 75 375 78 
rect 372 78 375 81 
rect 372 81 375 84 
rect 372 84 375 87 
rect 372 87 375 90 
rect 372 90 375 93 
rect 372 93 375 96 
rect 372 96 375 99 
rect 372 99 375 102 
rect 372 102 375 105 
rect 372 105 375 108 
rect 372 108 375 111 
rect 372 111 375 114 
rect 372 114 375 117 
rect 372 117 375 120 
rect 372 120 375 123 
rect 372 123 375 126 
rect 372 126 375 129 
rect 372 129 375 132 
rect 372 132 375 135 
rect 372 135 375 138 
rect 372 138 375 141 
rect 372 141 375 144 
rect 372 144 375 147 
rect 372 147 375 150 
rect 372 150 375 153 
rect 372 153 375 156 
rect 372 156 375 159 
rect 372 159 375 162 
rect 372 162 375 165 
rect 372 165 375 168 
rect 372 168 375 171 
rect 372 171 375 174 
rect 372 174 375 177 
rect 372 177 375 180 
rect 372 180 375 183 
rect 372 183 375 186 
rect 372 186 375 189 
rect 372 189 375 192 
rect 372 192 375 195 
rect 372 195 375 198 
rect 372 198 375 201 
rect 372 201 375 204 
rect 372 204 375 207 
rect 372 207 375 210 
rect 372 210 375 213 
rect 372 213 375 216 
rect 372 216 375 219 
rect 372 219 375 222 
rect 372 222 375 225 
rect 372 225 375 228 
rect 372 228 375 231 
rect 372 231 375 234 
rect 372 234 375 237 
rect 372 237 375 240 
rect 372 240 375 243 
rect 372 243 375 246 
rect 372 246 375 249 
rect 372 249 375 252 
rect 372 252 375 255 
rect 372 255 375 258 
rect 372 258 375 261 
rect 372 261 375 264 
rect 372 264 375 267 
rect 372 267 375 270 
rect 372 270 375 273 
rect 372 273 375 276 
rect 372 276 375 279 
rect 372 279 375 282 
rect 372 282 375 285 
rect 372 285 375 288 
rect 372 288 375 291 
rect 372 291 375 294 
rect 372 294 375 297 
rect 372 297 375 300 
rect 372 300 375 303 
rect 372 303 375 306 
rect 372 306 375 309 
rect 372 309 375 312 
rect 372 312 375 315 
rect 372 315 375 318 
rect 372 318 375 321 
rect 372 321 375 324 
rect 372 324 375 327 
rect 372 327 375 330 
rect 372 330 375 333 
rect 372 333 375 336 
rect 372 336 375 339 
rect 372 339 375 342 
rect 372 342 375 345 
rect 372 345 375 348 
rect 372 348 375 351 
rect 372 351 375 354 
rect 372 354 375 357 
rect 372 357 375 360 
rect 372 360 375 363 
rect 372 363 375 366 
rect 372 366 375 369 
rect 372 369 375 372 
rect 372 372 375 375 
rect 372 375 375 378 
rect 372 378 375 381 
rect 372 381 375 384 
rect 372 384 375 387 
rect 372 387 375 390 
rect 372 390 375 393 
rect 372 393 375 396 
rect 372 396 375 399 
rect 372 399 375 402 
rect 372 402 375 405 
rect 372 405 375 408 
rect 372 408 375 411 
rect 372 411 375 414 
rect 372 414 375 417 
rect 372 417 375 420 
rect 372 420 375 423 
rect 372 423 375 426 
rect 372 426 375 429 
rect 372 429 375 432 
rect 372 432 375 435 
rect 372 435 375 438 
rect 372 438 375 441 
rect 372 441 375 444 
rect 372 444 375 447 
rect 372 447 375 450 
rect 372 450 375 453 
rect 372 453 375 456 
rect 372 456 375 459 
rect 372 459 375 462 
rect 372 462 375 465 
rect 372 465 375 468 
rect 372 468 375 471 
rect 372 471 375 474 
rect 372 474 375 477 
rect 372 477 375 480 
rect 372 480 375 483 
rect 372 483 375 486 
rect 372 486 375 489 
rect 372 489 375 492 
rect 372 492 375 495 
rect 372 495 375 498 
rect 372 498 375 501 
rect 372 501 375 504 
rect 372 504 375 507 
rect 372 507 375 510 
rect 375 0 378 3 
rect 375 3 378 6 
rect 375 6 378 9 
rect 375 9 378 12 
rect 375 12 378 15 
rect 375 15 378 18 
rect 375 18 378 21 
rect 375 21 378 24 
rect 375 24 378 27 
rect 375 27 378 30 
rect 375 30 378 33 
rect 375 33 378 36 
rect 375 36 378 39 
rect 375 39 378 42 
rect 375 42 378 45 
rect 375 45 378 48 
rect 375 48 378 51 
rect 375 51 378 54 
rect 375 54 378 57 
rect 375 57 378 60 
rect 375 60 378 63 
rect 375 63 378 66 
rect 375 66 378 69 
rect 375 69 378 72 
rect 375 72 378 75 
rect 375 75 378 78 
rect 375 78 378 81 
rect 375 81 378 84 
rect 375 84 378 87 
rect 375 87 378 90 
rect 375 90 378 93 
rect 375 93 378 96 
rect 375 96 378 99 
rect 375 99 378 102 
rect 375 102 378 105 
rect 375 105 378 108 
rect 375 108 378 111 
rect 375 111 378 114 
rect 375 114 378 117 
rect 375 117 378 120 
rect 375 120 378 123 
rect 375 123 378 126 
rect 375 126 378 129 
rect 375 129 378 132 
rect 375 132 378 135 
rect 375 135 378 138 
rect 375 138 378 141 
rect 375 141 378 144 
rect 375 144 378 147 
rect 375 147 378 150 
rect 375 150 378 153 
rect 375 153 378 156 
rect 375 156 378 159 
rect 375 159 378 162 
rect 375 162 378 165 
rect 375 165 378 168 
rect 375 168 378 171 
rect 375 171 378 174 
rect 375 174 378 177 
rect 375 177 378 180 
rect 375 180 378 183 
rect 375 183 378 186 
rect 375 186 378 189 
rect 375 189 378 192 
rect 375 192 378 195 
rect 375 195 378 198 
rect 375 198 378 201 
rect 375 201 378 204 
rect 375 204 378 207 
rect 375 207 378 210 
rect 375 210 378 213 
rect 375 213 378 216 
rect 375 216 378 219 
rect 375 219 378 222 
rect 375 222 378 225 
rect 375 225 378 228 
rect 375 228 378 231 
rect 375 231 378 234 
rect 375 234 378 237 
rect 375 237 378 240 
rect 375 240 378 243 
rect 375 243 378 246 
rect 375 246 378 249 
rect 375 249 378 252 
rect 375 252 378 255 
rect 375 255 378 258 
rect 375 258 378 261 
rect 375 261 378 264 
rect 375 264 378 267 
rect 375 267 378 270 
rect 375 270 378 273 
rect 375 273 378 276 
rect 375 276 378 279 
rect 375 279 378 282 
rect 375 282 378 285 
rect 375 285 378 288 
rect 375 288 378 291 
rect 375 291 378 294 
rect 375 294 378 297 
rect 375 297 378 300 
rect 375 300 378 303 
rect 375 303 378 306 
rect 375 306 378 309 
rect 375 309 378 312 
rect 375 312 378 315 
rect 375 315 378 318 
rect 375 318 378 321 
rect 375 321 378 324 
rect 375 324 378 327 
rect 375 327 378 330 
rect 375 330 378 333 
rect 375 333 378 336 
rect 375 336 378 339 
rect 375 339 378 342 
rect 375 342 378 345 
rect 375 345 378 348 
rect 375 348 378 351 
rect 375 351 378 354 
rect 375 354 378 357 
rect 375 357 378 360 
rect 375 360 378 363 
rect 375 363 378 366 
rect 375 366 378 369 
rect 375 369 378 372 
rect 375 372 378 375 
rect 375 375 378 378 
rect 375 378 378 381 
rect 375 381 378 384 
rect 375 384 378 387 
rect 375 387 378 390 
rect 375 390 378 393 
rect 375 393 378 396 
rect 375 396 378 399 
rect 375 399 378 402 
rect 375 402 378 405 
rect 375 405 378 408 
rect 375 408 378 411 
rect 375 411 378 414 
rect 375 414 378 417 
rect 375 417 378 420 
rect 375 420 378 423 
rect 375 423 378 426 
rect 375 426 378 429 
rect 375 429 378 432 
rect 375 432 378 435 
rect 375 435 378 438 
rect 375 438 378 441 
rect 375 441 378 444 
rect 375 444 378 447 
rect 375 447 378 450 
rect 375 450 378 453 
rect 375 453 378 456 
rect 375 456 378 459 
rect 375 459 378 462 
rect 375 462 378 465 
rect 375 465 378 468 
rect 375 468 378 471 
rect 375 471 378 474 
rect 375 474 378 477 
rect 375 477 378 480 
rect 375 480 378 483 
rect 375 483 378 486 
rect 375 486 378 489 
rect 375 489 378 492 
rect 375 492 378 495 
rect 375 495 378 498 
rect 375 498 378 501 
rect 375 501 378 504 
rect 375 504 378 507 
rect 375 507 378 510 
rect 378 0 381 3 
rect 378 3 381 6 
rect 378 6 381 9 
rect 378 9 381 12 
rect 378 12 381 15 
rect 378 15 381 18 
rect 378 18 381 21 
rect 378 21 381 24 
rect 378 24 381 27 
rect 378 27 381 30 
rect 378 30 381 33 
rect 378 33 381 36 
rect 378 36 381 39 
rect 378 39 381 42 
rect 378 42 381 45 
rect 378 45 381 48 
rect 378 48 381 51 
rect 378 51 381 54 
rect 378 54 381 57 
rect 378 57 381 60 
rect 378 60 381 63 
rect 378 63 381 66 
rect 378 66 381 69 
rect 378 69 381 72 
rect 378 72 381 75 
rect 378 75 381 78 
rect 378 78 381 81 
rect 378 81 381 84 
rect 378 84 381 87 
rect 378 87 381 90 
rect 378 90 381 93 
rect 378 93 381 96 
rect 378 96 381 99 
rect 378 99 381 102 
rect 378 102 381 105 
rect 378 105 381 108 
rect 378 108 381 111 
rect 378 111 381 114 
rect 378 114 381 117 
rect 378 117 381 120 
rect 378 120 381 123 
rect 378 123 381 126 
rect 378 126 381 129 
rect 378 129 381 132 
rect 378 132 381 135 
rect 378 135 381 138 
rect 378 138 381 141 
rect 378 141 381 144 
rect 378 144 381 147 
rect 378 147 381 150 
rect 378 150 381 153 
rect 378 153 381 156 
rect 378 156 381 159 
rect 378 159 381 162 
rect 378 162 381 165 
rect 378 165 381 168 
rect 378 168 381 171 
rect 378 171 381 174 
rect 378 174 381 177 
rect 378 177 381 180 
rect 378 180 381 183 
rect 378 183 381 186 
rect 378 186 381 189 
rect 378 189 381 192 
rect 378 192 381 195 
rect 378 195 381 198 
rect 378 198 381 201 
rect 378 201 381 204 
rect 378 204 381 207 
rect 378 207 381 210 
rect 378 210 381 213 
rect 378 213 381 216 
rect 378 216 381 219 
rect 378 219 381 222 
rect 378 222 381 225 
rect 378 225 381 228 
rect 378 228 381 231 
rect 378 231 381 234 
rect 378 234 381 237 
rect 378 237 381 240 
rect 378 240 381 243 
rect 378 243 381 246 
rect 378 246 381 249 
rect 378 249 381 252 
rect 378 252 381 255 
rect 378 255 381 258 
rect 378 258 381 261 
rect 378 261 381 264 
rect 378 264 381 267 
rect 378 267 381 270 
rect 378 270 381 273 
rect 378 273 381 276 
rect 378 276 381 279 
rect 378 279 381 282 
rect 378 282 381 285 
rect 378 285 381 288 
rect 378 288 381 291 
rect 378 291 381 294 
rect 378 294 381 297 
rect 378 297 381 300 
rect 378 300 381 303 
rect 378 303 381 306 
rect 378 306 381 309 
rect 378 309 381 312 
rect 378 312 381 315 
rect 378 315 381 318 
rect 378 318 381 321 
rect 378 321 381 324 
rect 378 324 381 327 
rect 378 327 381 330 
rect 378 330 381 333 
rect 378 333 381 336 
rect 378 336 381 339 
rect 378 339 381 342 
rect 378 342 381 345 
rect 378 345 381 348 
rect 378 348 381 351 
rect 378 351 381 354 
rect 378 354 381 357 
rect 378 357 381 360 
rect 378 360 381 363 
rect 378 363 381 366 
rect 378 366 381 369 
rect 378 369 381 372 
rect 378 372 381 375 
rect 378 375 381 378 
rect 378 378 381 381 
rect 378 381 381 384 
rect 378 384 381 387 
rect 378 387 381 390 
rect 378 390 381 393 
rect 378 393 381 396 
rect 378 396 381 399 
rect 378 399 381 402 
rect 378 402 381 405 
rect 378 405 381 408 
rect 378 408 381 411 
rect 378 411 381 414 
rect 378 414 381 417 
rect 378 417 381 420 
rect 378 420 381 423 
rect 378 423 381 426 
rect 378 426 381 429 
rect 378 429 381 432 
rect 378 432 381 435 
rect 378 435 381 438 
rect 378 438 381 441 
rect 378 441 381 444 
rect 378 444 381 447 
rect 378 447 381 450 
rect 378 450 381 453 
rect 378 453 381 456 
rect 378 456 381 459 
rect 378 459 381 462 
rect 378 462 381 465 
rect 378 465 381 468 
rect 378 468 381 471 
rect 378 471 381 474 
rect 378 474 381 477 
rect 378 477 381 480 
rect 378 480 381 483 
rect 378 483 381 486 
rect 378 486 381 489 
rect 378 489 381 492 
rect 378 492 381 495 
rect 378 495 381 498 
rect 378 498 381 501 
rect 378 501 381 504 
rect 378 504 381 507 
rect 378 507 381 510 
rect 381 0 384 3 
rect 381 3 384 6 
rect 381 6 384 9 
rect 381 9 384 12 
rect 381 12 384 15 
rect 381 15 384 18 
rect 381 18 384 21 
rect 381 21 384 24 
rect 381 24 384 27 
rect 381 27 384 30 
rect 381 30 384 33 
rect 381 33 384 36 
rect 381 36 384 39 
rect 381 39 384 42 
rect 381 42 384 45 
rect 381 45 384 48 
rect 381 48 384 51 
rect 381 51 384 54 
rect 381 54 384 57 
rect 381 57 384 60 
rect 381 60 384 63 
rect 381 63 384 66 
rect 381 66 384 69 
rect 381 69 384 72 
rect 381 72 384 75 
rect 381 75 384 78 
rect 381 78 384 81 
rect 381 81 384 84 
rect 381 84 384 87 
rect 381 87 384 90 
rect 381 90 384 93 
rect 381 93 384 96 
rect 381 96 384 99 
rect 381 99 384 102 
rect 381 102 384 105 
rect 381 105 384 108 
rect 381 108 384 111 
rect 381 111 384 114 
rect 381 114 384 117 
rect 381 117 384 120 
rect 381 120 384 123 
rect 381 123 384 126 
rect 381 126 384 129 
rect 381 129 384 132 
rect 381 132 384 135 
rect 381 135 384 138 
rect 381 138 384 141 
rect 381 141 384 144 
rect 381 144 384 147 
rect 381 147 384 150 
rect 381 150 384 153 
rect 381 153 384 156 
rect 381 156 384 159 
rect 381 159 384 162 
rect 381 162 384 165 
rect 381 165 384 168 
rect 381 168 384 171 
rect 381 171 384 174 
rect 381 174 384 177 
rect 381 177 384 180 
rect 381 180 384 183 
rect 381 183 384 186 
rect 381 186 384 189 
rect 381 189 384 192 
rect 381 192 384 195 
rect 381 195 384 198 
rect 381 198 384 201 
rect 381 201 384 204 
rect 381 204 384 207 
rect 381 207 384 210 
rect 381 210 384 213 
rect 381 213 384 216 
rect 381 216 384 219 
rect 381 219 384 222 
rect 381 222 384 225 
rect 381 225 384 228 
rect 381 228 384 231 
rect 381 231 384 234 
rect 381 234 384 237 
rect 381 237 384 240 
rect 381 240 384 243 
rect 381 243 384 246 
rect 381 246 384 249 
rect 381 249 384 252 
rect 381 252 384 255 
rect 381 255 384 258 
rect 381 258 384 261 
rect 381 261 384 264 
rect 381 264 384 267 
rect 381 267 384 270 
rect 381 270 384 273 
rect 381 273 384 276 
rect 381 276 384 279 
rect 381 279 384 282 
rect 381 282 384 285 
rect 381 285 384 288 
rect 381 288 384 291 
rect 381 291 384 294 
rect 381 294 384 297 
rect 381 297 384 300 
rect 381 300 384 303 
rect 381 303 384 306 
rect 381 306 384 309 
rect 381 309 384 312 
rect 381 312 384 315 
rect 381 315 384 318 
rect 381 318 384 321 
rect 381 321 384 324 
rect 381 324 384 327 
rect 381 327 384 330 
rect 381 330 384 333 
rect 381 333 384 336 
rect 381 336 384 339 
rect 381 339 384 342 
rect 381 342 384 345 
rect 381 345 384 348 
rect 381 348 384 351 
rect 381 351 384 354 
rect 381 354 384 357 
rect 381 357 384 360 
rect 381 360 384 363 
rect 381 363 384 366 
rect 381 366 384 369 
rect 381 369 384 372 
rect 381 372 384 375 
rect 381 375 384 378 
rect 381 378 384 381 
rect 381 381 384 384 
rect 381 384 384 387 
rect 381 387 384 390 
rect 381 390 384 393 
rect 381 393 384 396 
rect 381 396 384 399 
rect 381 399 384 402 
rect 381 402 384 405 
rect 381 405 384 408 
rect 381 408 384 411 
rect 381 411 384 414 
rect 381 414 384 417 
rect 381 417 384 420 
rect 381 420 384 423 
rect 381 423 384 426 
rect 381 426 384 429 
rect 381 429 384 432 
rect 381 432 384 435 
rect 381 435 384 438 
rect 381 438 384 441 
rect 381 441 384 444 
rect 381 444 384 447 
rect 381 447 384 450 
rect 381 450 384 453 
rect 381 453 384 456 
rect 381 456 384 459 
rect 381 459 384 462 
rect 381 462 384 465 
rect 381 465 384 468 
rect 381 468 384 471 
rect 381 471 384 474 
rect 381 474 384 477 
rect 381 477 384 480 
rect 381 480 384 483 
rect 381 483 384 486 
rect 381 486 384 489 
rect 381 489 384 492 
rect 381 492 384 495 
rect 381 495 384 498 
rect 381 498 384 501 
rect 381 501 384 504 
rect 381 504 384 507 
rect 381 507 384 510 
rect 384 0 387 3 
rect 384 3 387 6 
rect 384 6 387 9 
rect 384 9 387 12 
rect 384 12 387 15 
rect 384 15 387 18 
rect 384 18 387 21 
rect 384 21 387 24 
rect 384 24 387 27 
rect 384 27 387 30 
rect 384 30 387 33 
rect 384 33 387 36 
rect 384 36 387 39 
rect 384 39 387 42 
rect 384 42 387 45 
rect 384 45 387 48 
rect 384 48 387 51 
rect 384 51 387 54 
rect 384 54 387 57 
rect 384 57 387 60 
rect 384 60 387 63 
rect 384 63 387 66 
rect 384 66 387 69 
rect 384 69 387 72 
rect 384 72 387 75 
rect 384 75 387 78 
rect 384 78 387 81 
rect 384 81 387 84 
rect 384 84 387 87 
rect 384 87 387 90 
rect 384 90 387 93 
rect 384 93 387 96 
rect 384 96 387 99 
rect 384 99 387 102 
rect 384 102 387 105 
rect 384 105 387 108 
rect 384 108 387 111 
rect 384 111 387 114 
rect 384 114 387 117 
rect 384 117 387 120 
rect 384 120 387 123 
rect 384 123 387 126 
rect 384 126 387 129 
rect 384 129 387 132 
rect 384 132 387 135 
rect 384 135 387 138 
rect 384 138 387 141 
rect 384 141 387 144 
rect 384 144 387 147 
rect 384 147 387 150 
rect 384 150 387 153 
rect 384 153 387 156 
rect 384 156 387 159 
rect 384 159 387 162 
rect 384 162 387 165 
rect 384 165 387 168 
rect 384 168 387 171 
rect 384 171 387 174 
rect 384 174 387 177 
rect 384 177 387 180 
rect 384 180 387 183 
rect 384 183 387 186 
rect 384 186 387 189 
rect 384 189 387 192 
rect 384 192 387 195 
rect 384 195 387 198 
rect 384 198 387 201 
rect 384 201 387 204 
rect 384 204 387 207 
rect 384 207 387 210 
rect 384 210 387 213 
rect 384 213 387 216 
rect 384 216 387 219 
rect 384 219 387 222 
rect 384 222 387 225 
rect 384 225 387 228 
rect 384 228 387 231 
rect 384 231 387 234 
rect 384 234 387 237 
rect 384 237 387 240 
rect 384 240 387 243 
rect 384 243 387 246 
rect 384 246 387 249 
rect 384 249 387 252 
rect 384 252 387 255 
rect 384 255 387 258 
rect 384 258 387 261 
rect 384 261 387 264 
rect 384 264 387 267 
rect 384 267 387 270 
rect 384 270 387 273 
rect 384 273 387 276 
rect 384 276 387 279 
rect 384 279 387 282 
rect 384 282 387 285 
rect 384 285 387 288 
rect 384 288 387 291 
rect 384 291 387 294 
rect 384 294 387 297 
rect 384 297 387 300 
rect 384 300 387 303 
rect 384 303 387 306 
rect 384 306 387 309 
rect 384 309 387 312 
rect 384 312 387 315 
rect 384 315 387 318 
rect 384 318 387 321 
rect 384 321 387 324 
rect 384 324 387 327 
rect 384 327 387 330 
rect 384 330 387 333 
rect 384 333 387 336 
rect 384 336 387 339 
rect 384 339 387 342 
rect 384 342 387 345 
rect 384 345 387 348 
rect 384 348 387 351 
rect 384 351 387 354 
rect 384 354 387 357 
rect 384 357 387 360 
rect 384 360 387 363 
rect 384 363 387 366 
rect 384 366 387 369 
rect 384 369 387 372 
rect 384 372 387 375 
rect 384 375 387 378 
rect 384 378 387 381 
rect 384 381 387 384 
rect 384 384 387 387 
rect 384 387 387 390 
rect 384 390 387 393 
rect 384 393 387 396 
rect 384 396 387 399 
rect 384 399 387 402 
rect 384 402 387 405 
rect 384 405 387 408 
rect 384 408 387 411 
rect 384 411 387 414 
rect 384 414 387 417 
rect 384 417 387 420 
rect 384 420 387 423 
rect 384 423 387 426 
rect 384 426 387 429 
rect 384 429 387 432 
rect 384 432 387 435 
rect 384 435 387 438 
rect 384 438 387 441 
rect 384 441 387 444 
rect 384 444 387 447 
rect 384 447 387 450 
rect 384 450 387 453 
rect 384 453 387 456 
rect 384 456 387 459 
rect 384 459 387 462 
rect 384 462 387 465 
rect 384 465 387 468 
rect 384 468 387 471 
rect 384 471 387 474 
rect 384 474 387 477 
rect 384 477 387 480 
rect 384 480 387 483 
rect 384 483 387 486 
rect 384 486 387 489 
rect 384 489 387 492 
rect 384 492 387 495 
rect 384 495 387 498 
rect 384 498 387 501 
rect 384 501 387 504 
rect 384 504 387 507 
rect 384 507 387 510 
rect 387 0 390 3 
rect 387 3 390 6 
rect 387 6 390 9 
rect 387 9 390 12 
rect 387 12 390 15 
rect 387 15 390 18 
rect 387 18 390 21 
rect 387 21 390 24 
rect 387 24 390 27 
rect 387 27 390 30 
rect 387 30 390 33 
rect 387 33 390 36 
rect 387 36 390 39 
rect 387 39 390 42 
rect 387 42 390 45 
rect 387 45 390 48 
rect 387 48 390 51 
rect 387 51 390 54 
rect 387 54 390 57 
rect 387 57 390 60 
rect 387 60 390 63 
rect 387 63 390 66 
rect 387 66 390 69 
rect 387 69 390 72 
rect 387 72 390 75 
rect 387 75 390 78 
rect 387 78 390 81 
rect 387 81 390 84 
rect 387 84 390 87 
rect 387 87 390 90 
rect 387 90 390 93 
rect 387 93 390 96 
rect 387 96 390 99 
rect 387 99 390 102 
rect 387 102 390 105 
rect 387 105 390 108 
rect 387 108 390 111 
rect 387 111 390 114 
rect 387 114 390 117 
rect 387 117 390 120 
rect 387 120 390 123 
rect 387 123 390 126 
rect 387 126 390 129 
rect 387 129 390 132 
rect 387 132 390 135 
rect 387 135 390 138 
rect 387 138 390 141 
rect 387 141 390 144 
rect 387 144 390 147 
rect 387 147 390 150 
rect 387 150 390 153 
rect 387 153 390 156 
rect 387 156 390 159 
rect 387 159 390 162 
rect 387 162 390 165 
rect 387 165 390 168 
rect 387 168 390 171 
rect 387 171 390 174 
rect 387 174 390 177 
rect 387 177 390 180 
rect 387 180 390 183 
rect 387 183 390 186 
rect 387 186 390 189 
rect 387 189 390 192 
rect 387 192 390 195 
rect 387 195 390 198 
rect 387 198 390 201 
rect 387 201 390 204 
rect 387 204 390 207 
rect 387 207 390 210 
rect 387 210 390 213 
rect 387 213 390 216 
rect 387 216 390 219 
rect 387 219 390 222 
rect 387 222 390 225 
rect 387 225 390 228 
rect 387 228 390 231 
rect 387 231 390 234 
rect 387 234 390 237 
rect 387 237 390 240 
rect 387 240 390 243 
rect 387 243 390 246 
rect 387 246 390 249 
rect 387 249 390 252 
rect 387 252 390 255 
rect 387 255 390 258 
rect 387 258 390 261 
rect 387 261 390 264 
rect 387 264 390 267 
rect 387 267 390 270 
rect 387 270 390 273 
rect 387 273 390 276 
rect 387 276 390 279 
rect 387 279 390 282 
rect 387 282 390 285 
rect 387 285 390 288 
rect 387 288 390 291 
rect 387 291 390 294 
rect 387 294 390 297 
rect 387 297 390 300 
rect 387 300 390 303 
rect 387 303 390 306 
rect 387 306 390 309 
rect 387 309 390 312 
rect 387 312 390 315 
rect 387 315 390 318 
rect 387 318 390 321 
rect 387 321 390 324 
rect 387 324 390 327 
rect 387 327 390 330 
rect 387 330 390 333 
rect 387 333 390 336 
rect 387 336 390 339 
rect 387 339 390 342 
rect 387 342 390 345 
rect 387 345 390 348 
rect 387 348 390 351 
rect 387 351 390 354 
rect 387 354 390 357 
rect 387 357 390 360 
rect 387 360 390 363 
rect 387 363 390 366 
rect 387 366 390 369 
rect 387 369 390 372 
rect 387 372 390 375 
rect 387 375 390 378 
rect 387 378 390 381 
rect 387 381 390 384 
rect 387 384 390 387 
rect 387 387 390 390 
rect 387 390 390 393 
rect 387 393 390 396 
rect 387 396 390 399 
rect 387 399 390 402 
rect 387 402 390 405 
rect 387 405 390 408 
rect 387 408 390 411 
rect 387 411 390 414 
rect 387 414 390 417 
rect 387 417 390 420 
rect 387 420 390 423 
rect 387 423 390 426 
rect 387 426 390 429 
rect 387 429 390 432 
rect 387 432 390 435 
rect 387 435 390 438 
rect 387 438 390 441 
rect 387 441 390 444 
rect 387 444 390 447 
rect 387 447 390 450 
rect 387 450 390 453 
rect 387 453 390 456 
rect 387 456 390 459 
rect 387 459 390 462 
rect 387 462 390 465 
rect 387 465 390 468 
rect 387 468 390 471 
rect 387 471 390 474 
rect 387 474 390 477 
rect 387 477 390 480 
rect 387 480 390 483 
rect 387 483 390 486 
rect 387 486 390 489 
rect 387 489 390 492 
rect 387 492 390 495 
rect 387 495 390 498 
rect 387 498 390 501 
rect 387 501 390 504 
rect 387 504 390 507 
rect 387 507 390 510 
rect 390 0 393 3 
rect 390 3 393 6 
rect 390 6 393 9 
rect 390 9 393 12 
rect 390 12 393 15 
rect 390 15 393 18 
rect 390 18 393 21 
rect 390 21 393 24 
rect 390 24 393 27 
rect 390 27 393 30 
rect 390 30 393 33 
rect 390 33 393 36 
rect 390 36 393 39 
rect 390 39 393 42 
rect 390 42 393 45 
rect 390 45 393 48 
rect 390 48 393 51 
rect 390 51 393 54 
rect 390 54 393 57 
rect 390 57 393 60 
rect 390 60 393 63 
rect 390 63 393 66 
rect 390 66 393 69 
rect 390 69 393 72 
rect 390 72 393 75 
rect 390 75 393 78 
rect 390 78 393 81 
rect 390 81 393 84 
rect 390 84 393 87 
rect 390 87 393 90 
rect 390 90 393 93 
rect 390 93 393 96 
rect 390 96 393 99 
rect 390 99 393 102 
rect 390 102 393 105 
rect 390 105 393 108 
rect 390 108 393 111 
rect 390 111 393 114 
rect 390 114 393 117 
rect 390 117 393 120 
rect 390 120 393 123 
rect 390 123 393 126 
rect 390 126 393 129 
rect 390 129 393 132 
rect 390 132 393 135 
rect 390 135 393 138 
rect 390 138 393 141 
rect 390 141 393 144 
rect 390 144 393 147 
rect 390 147 393 150 
rect 390 150 393 153 
rect 390 153 393 156 
rect 390 156 393 159 
rect 390 159 393 162 
rect 390 162 393 165 
rect 390 165 393 168 
rect 390 168 393 171 
rect 390 171 393 174 
rect 390 174 393 177 
rect 390 177 393 180 
rect 390 180 393 183 
rect 390 183 393 186 
rect 390 186 393 189 
rect 390 189 393 192 
rect 390 192 393 195 
rect 390 195 393 198 
rect 390 198 393 201 
rect 390 201 393 204 
rect 390 204 393 207 
rect 390 207 393 210 
rect 390 210 393 213 
rect 390 213 393 216 
rect 390 216 393 219 
rect 390 219 393 222 
rect 390 222 393 225 
rect 390 225 393 228 
rect 390 228 393 231 
rect 390 231 393 234 
rect 390 234 393 237 
rect 390 237 393 240 
rect 390 240 393 243 
rect 390 243 393 246 
rect 390 246 393 249 
rect 390 249 393 252 
rect 390 252 393 255 
rect 390 255 393 258 
rect 390 258 393 261 
rect 390 261 393 264 
rect 390 264 393 267 
rect 390 267 393 270 
rect 390 270 393 273 
rect 390 273 393 276 
rect 390 276 393 279 
rect 390 279 393 282 
rect 390 282 393 285 
rect 390 285 393 288 
rect 390 288 393 291 
rect 390 291 393 294 
rect 390 294 393 297 
rect 390 297 393 300 
rect 390 300 393 303 
rect 390 303 393 306 
rect 390 306 393 309 
rect 390 309 393 312 
rect 390 312 393 315 
rect 390 315 393 318 
rect 390 318 393 321 
rect 390 321 393 324 
rect 390 324 393 327 
rect 390 327 393 330 
rect 390 330 393 333 
rect 390 333 393 336 
rect 390 336 393 339 
rect 390 339 393 342 
rect 390 342 393 345 
rect 390 345 393 348 
rect 390 348 393 351 
rect 390 351 393 354 
rect 390 354 393 357 
rect 390 357 393 360 
rect 390 360 393 363 
rect 390 363 393 366 
rect 390 366 393 369 
rect 390 369 393 372 
rect 390 372 393 375 
rect 390 375 393 378 
rect 390 378 393 381 
rect 390 381 393 384 
rect 390 384 393 387 
rect 390 387 393 390 
rect 390 390 393 393 
rect 390 393 393 396 
rect 390 396 393 399 
rect 390 399 393 402 
rect 390 402 393 405 
rect 390 405 393 408 
rect 390 408 393 411 
rect 390 411 393 414 
rect 390 414 393 417 
rect 390 417 393 420 
rect 390 420 393 423 
rect 390 423 393 426 
rect 390 426 393 429 
rect 390 429 393 432 
rect 390 432 393 435 
rect 390 435 393 438 
rect 390 438 393 441 
rect 390 441 393 444 
rect 390 444 393 447 
rect 390 447 393 450 
rect 390 450 393 453 
rect 390 453 393 456 
rect 390 456 393 459 
rect 390 459 393 462 
rect 390 462 393 465 
rect 390 465 393 468 
rect 390 468 393 471 
rect 390 471 393 474 
rect 390 474 393 477 
rect 390 477 393 480 
rect 390 480 393 483 
rect 390 483 393 486 
rect 390 486 393 489 
rect 390 489 393 492 
rect 390 492 393 495 
rect 390 495 393 498 
rect 390 498 393 501 
rect 390 501 393 504 
rect 390 504 393 507 
rect 390 507 393 510 
rect 393 0 396 3 
rect 393 3 396 6 
rect 393 6 396 9 
rect 393 9 396 12 
rect 393 12 396 15 
rect 393 15 396 18 
rect 393 18 396 21 
rect 393 21 396 24 
rect 393 24 396 27 
rect 393 27 396 30 
rect 393 30 396 33 
rect 393 33 396 36 
rect 393 36 396 39 
rect 393 39 396 42 
rect 393 42 396 45 
rect 393 45 396 48 
rect 393 48 396 51 
rect 393 51 396 54 
rect 393 54 396 57 
rect 393 57 396 60 
rect 393 60 396 63 
rect 393 63 396 66 
rect 393 66 396 69 
rect 393 69 396 72 
rect 393 72 396 75 
rect 393 75 396 78 
rect 393 78 396 81 
rect 393 81 396 84 
rect 393 84 396 87 
rect 393 87 396 90 
rect 393 90 396 93 
rect 393 93 396 96 
rect 393 96 396 99 
rect 393 99 396 102 
rect 393 102 396 105 
rect 393 105 396 108 
rect 393 108 396 111 
rect 393 111 396 114 
rect 393 114 396 117 
rect 393 117 396 120 
rect 393 120 396 123 
rect 393 123 396 126 
rect 393 126 396 129 
rect 393 129 396 132 
rect 393 132 396 135 
rect 393 135 396 138 
rect 393 138 396 141 
rect 393 141 396 144 
rect 393 144 396 147 
rect 393 147 396 150 
rect 393 150 396 153 
rect 393 153 396 156 
rect 393 156 396 159 
rect 393 159 396 162 
rect 393 162 396 165 
rect 393 165 396 168 
rect 393 168 396 171 
rect 393 171 396 174 
rect 393 174 396 177 
rect 393 177 396 180 
rect 393 180 396 183 
rect 393 183 396 186 
rect 393 186 396 189 
rect 393 189 396 192 
rect 393 192 396 195 
rect 393 195 396 198 
rect 393 198 396 201 
rect 393 201 396 204 
rect 393 204 396 207 
rect 393 207 396 210 
rect 393 210 396 213 
rect 393 213 396 216 
rect 393 216 396 219 
rect 393 219 396 222 
rect 393 222 396 225 
rect 393 225 396 228 
rect 393 228 396 231 
rect 393 231 396 234 
rect 393 234 396 237 
rect 393 237 396 240 
rect 393 240 396 243 
rect 393 243 396 246 
rect 393 246 396 249 
rect 393 249 396 252 
rect 393 252 396 255 
rect 393 255 396 258 
rect 393 258 396 261 
rect 393 261 396 264 
rect 393 264 396 267 
rect 393 267 396 270 
rect 393 270 396 273 
rect 393 273 396 276 
rect 393 276 396 279 
rect 393 279 396 282 
rect 393 282 396 285 
rect 393 285 396 288 
rect 393 288 396 291 
rect 393 291 396 294 
rect 393 294 396 297 
rect 393 297 396 300 
rect 393 300 396 303 
rect 393 303 396 306 
rect 393 306 396 309 
rect 393 309 396 312 
rect 393 312 396 315 
rect 393 315 396 318 
rect 393 318 396 321 
rect 393 321 396 324 
rect 393 324 396 327 
rect 393 327 396 330 
rect 393 330 396 333 
rect 393 333 396 336 
rect 393 336 396 339 
rect 393 339 396 342 
rect 393 342 396 345 
rect 393 345 396 348 
rect 393 348 396 351 
rect 393 351 396 354 
rect 393 354 396 357 
rect 393 357 396 360 
rect 393 360 396 363 
rect 393 363 396 366 
rect 393 366 396 369 
rect 393 369 396 372 
rect 393 372 396 375 
rect 393 375 396 378 
rect 393 378 396 381 
rect 393 381 396 384 
rect 393 384 396 387 
rect 393 387 396 390 
rect 393 390 396 393 
rect 393 393 396 396 
rect 393 396 396 399 
rect 393 399 396 402 
rect 393 402 396 405 
rect 393 405 396 408 
rect 393 408 396 411 
rect 393 411 396 414 
rect 393 414 396 417 
rect 393 417 396 420 
rect 393 420 396 423 
rect 393 423 396 426 
rect 393 426 396 429 
rect 393 429 396 432 
rect 393 432 396 435 
rect 393 435 396 438 
rect 393 438 396 441 
rect 393 441 396 444 
rect 393 444 396 447 
rect 393 447 396 450 
rect 393 450 396 453 
rect 393 453 396 456 
rect 393 456 396 459 
rect 393 459 396 462 
rect 393 462 396 465 
rect 393 465 396 468 
rect 393 468 396 471 
rect 393 471 396 474 
rect 393 474 396 477 
rect 393 477 396 480 
rect 393 480 396 483 
rect 393 483 396 486 
rect 393 486 396 489 
rect 393 489 396 492 
rect 393 492 396 495 
rect 393 495 396 498 
rect 393 498 396 501 
rect 393 501 396 504 
rect 393 504 396 507 
rect 393 507 396 510 
rect 396 0 399 3 
rect 396 3 399 6 
rect 396 6 399 9 
rect 396 9 399 12 
rect 396 12 399 15 
rect 396 15 399 18 
rect 396 18 399 21 
rect 396 21 399 24 
rect 396 24 399 27 
rect 396 27 399 30 
rect 396 30 399 33 
rect 396 33 399 36 
rect 396 36 399 39 
rect 396 39 399 42 
rect 396 42 399 45 
rect 396 45 399 48 
rect 396 48 399 51 
rect 396 51 399 54 
rect 396 54 399 57 
rect 396 57 399 60 
rect 396 60 399 63 
rect 396 63 399 66 
rect 396 66 399 69 
rect 396 69 399 72 
rect 396 72 399 75 
rect 396 75 399 78 
rect 396 78 399 81 
rect 396 81 399 84 
rect 396 84 399 87 
rect 396 87 399 90 
rect 396 90 399 93 
rect 396 93 399 96 
rect 396 96 399 99 
rect 396 99 399 102 
rect 396 102 399 105 
rect 396 105 399 108 
rect 396 108 399 111 
rect 396 111 399 114 
rect 396 114 399 117 
rect 396 117 399 120 
rect 396 120 399 123 
rect 396 123 399 126 
rect 396 126 399 129 
rect 396 129 399 132 
rect 396 132 399 135 
rect 396 135 399 138 
rect 396 138 399 141 
rect 396 141 399 144 
rect 396 144 399 147 
rect 396 147 399 150 
rect 396 150 399 153 
rect 396 153 399 156 
rect 396 156 399 159 
rect 396 159 399 162 
rect 396 162 399 165 
rect 396 165 399 168 
rect 396 168 399 171 
rect 396 171 399 174 
rect 396 174 399 177 
rect 396 177 399 180 
rect 396 180 399 183 
rect 396 183 399 186 
rect 396 186 399 189 
rect 396 189 399 192 
rect 396 192 399 195 
rect 396 195 399 198 
rect 396 198 399 201 
rect 396 201 399 204 
rect 396 204 399 207 
rect 396 207 399 210 
rect 396 210 399 213 
rect 396 213 399 216 
rect 396 216 399 219 
rect 396 219 399 222 
rect 396 222 399 225 
rect 396 225 399 228 
rect 396 228 399 231 
rect 396 231 399 234 
rect 396 234 399 237 
rect 396 237 399 240 
rect 396 240 399 243 
rect 396 243 399 246 
rect 396 246 399 249 
rect 396 249 399 252 
rect 396 252 399 255 
rect 396 255 399 258 
rect 396 258 399 261 
rect 396 261 399 264 
rect 396 264 399 267 
rect 396 267 399 270 
rect 396 270 399 273 
rect 396 273 399 276 
rect 396 276 399 279 
rect 396 279 399 282 
rect 396 282 399 285 
rect 396 285 399 288 
rect 396 288 399 291 
rect 396 291 399 294 
rect 396 294 399 297 
rect 396 297 399 300 
rect 396 300 399 303 
rect 396 303 399 306 
rect 396 306 399 309 
rect 396 309 399 312 
rect 396 312 399 315 
rect 396 315 399 318 
rect 396 318 399 321 
rect 396 321 399 324 
rect 396 324 399 327 
rect 396 327 399 330 
rect 396 330 399 333 
rect 396 333 399 336 
rect 396 336 399 339 
rect 396 339 399 342 
rect 396 342 399 345 
rect 396 345 399 348 
rect 396 348 399 351 
rect 396 351 399 354 
rect 396 354 399 357 
rect 396 357 399 360 
rect 396 360 399 363 
rect 396 363 399 366 
rect 396 366 399 369 
rect 396 369 399 372 
rect 396 372 399 375 
rect 396 375 399 378 
rect 396 378 399 381 
rect 396 381 399 384 
rect 396 384 399 387 
rect 396 387 399 390 
rect 396 390 399 393 
rect 396 393 399 396 
rect 396 396 399 399 
rect 396 399 399 402 
rect 396 402 399 405 
rect 396 405 399 408 
rect 396 408 399 411 
rect 396 411 399 414 
rect 396 414 399 417 
rect 396 417 399 420 
rect 396 420 399 423 
rect 396 423 399 426 
rect 396 426 399 429 
rect 396 429 399 432 
rect 396 432 399 435 
rect 396 435 399 438 
rect 396 438 399 441 
rect 396 441 399 444 
rect 396 444 399 447 
rect 396 447 399 450 
rect 396 450 399 453 
rect 396 453 399 456 
rect 396 456 399 459 
rect 396 459 399 462 
rect 396 462 399 465 
rect 396 465 399 468 
rect 396 468 399 471 
rect 396 471 399 474 
rect 396 474 399 477 
rect 396 477 399 480 
rect 396 480 399 483 
rect 396 483 399 486 
rect 396 486 399 489 
rect 396 489 399 492 
rect 396 492 399 495 
rect 396 495 399 498 
rect 396 498 399 501 
rect 396 501 399 504 
rect 396 504 399 507 
rect 396 507 399 510 
rect 399 0 402 3 
rect 399 3 402 6 
rect 399 6 402 9 
rect 399 9 402 12 
rect 399 12 402 15 
rect 399 15 402 18 
rect 399 18 402 21 
rect 399 21 402 24 
rect 399 24 402 27 
rect 399 27 402 30 
rect 399 30 402 33 
rect 399 33 402 36 
rect 399 36 402 39 
rect 399 39 402 42 
rect 399 42 402 45 
rect 399 45 402 48 
rect 399 48 402 51 
rect 399 51 402 54 
rect 399 54 402 57 
rect 399 57 402 60 
rect 399 60 402 63 
rect 399 63 402 66 
rect 399 66 402 69 
rect 399 69 402 72 
rect 399 72 402 75 
rect 399 75 402 78 
rect 399 78 402 81 
rect 399 81 402 84 
rect 399 84 402 87 
rect 399 87 402 90 
rect 399 90 402 93 
rect 399 93 402 96 
rect 399 96 402 99 
rect 399 99 402 102 
rect 399 102 402 105 
rect 399 105 402 108 
rect 399 108 402 111 
rect 399 111 402 114 
rect 399 114 402 117 
rect 399 117 402 120 
rect 399 120 402 123 
rect 399 123 402 126 
rect 399 126 402 129 
rect 399 129 402 132 
rect 399 132 402 135 
rect 399 135 402 138 
rect 399 138 402 141 
rect 399 141 402 144 
rect 399 144 402 147 
rect 399 147 402 150 
rect 399 150 402 153 
rect 399 153 402 156 
rect 399 156 402 159 
rect 399 159 402 162 
rect 399 162 402 165 
rect 399 165 402 168 
rect 399 168 402 171 
rect 399 171 402 174 
rect 399 174 402 177 
rect 399 177 402 180 
rect 399 180 402 183 
rect 399 183 402 186 
rect 399 186 402 189 
rect 399 189 402 192 
rect 399 192 402 195 
rect 399 195 402 198 
rect 399 198 402 201 
rect 399 201 402 204 
rect 399 204 402 207 
rect 399 207 402 210 
rect 399 210 402 213 
rect 399 213 402 216 
rect 399 216 402 219 
rect 399 219 402 222 
rect 399 222 402 225 
rect 399 225 402 228 
rect 399 228 402 231 
rect 399 231 402 234 
rect 399 234 402 237 
rect 399 237 402 240 
rect 399 240 402 243 
rect 399 243 402 246 
rect 399 246 402 249 
rect 399 249 402 252 
rect 399 252 402 255 
rect 399 255 402 258 
rect 399 258 402 261 
rect 399 261 402 264 
rect 399 264 402 267 
rect 399 267 402 270 
rect 399 270 402 273 
rect 399 273 402 276 
rect 399 276 402 279 
rect 399 279 402 282 
rect 399 282 402 285 
rect 399 285 402 288 
rect 399 288 402 291 
rect 399 291 402 294 
rect 399 294 402 297 
rect 399 297 402 300 
rect 399 300 402 303 
rect 399 303 402 306 
rect 399 306 402 309 
rect 399 309 402 312 
rect 399 312 402 315 
rect 399 315 402 318 
rect 399 318 402 321 
rect 399 321 402 324 
rect 399 324 402 327 
rect 399 327 402 330 
rect 399 330 402 333 
rect 399 333 402 336 
rect 399 336 402 339 
rect 399 339 402 342 
rect 399 342 402 345 
rect 399 345 402 348 
rect 399 348 402 351 
rect 399 351 402 354 
rect 399 354 402 357 
rect 399 357 402 360 
rect 399 360 402 363 
rect 399 363 402 366 
rect 399 366 402 369 
rect 399 369 402 372 
rect 399 372 402 375 
rect 399 375 402 378 
rect 399 378 402 381 
rect 399 381 402 384 
rect 399 384 402 387 
rect 399 387 402 390 
rect 399 390 402 393 
rect 399 393 402 396 
rect 399 396 402 399 
rect 399 399 402 402 
rect 399 402 402 405 
rect 399 405 402 408 
rect 399 408 402 411 
rect 399 411 402 414 
rect 399 414 402 417 
rect 399 417 402 420 
rect 399 420 402 423 
rect 399 423 402 426 
rect 399 426 402 429 
rect 399 429 402 432 
rect 399 432 402 435 
rect 399 435 402 438 
rect 399 438 402 441 
rect 399 441 402 444 
rect 399 444 402 447 
rect 399 447 402 450 
rect 399 450 402 453 
rect 399 453 402 456 
rect 399 456 402 459 
rect 399 459 402 462 
rect 399 462 402 465 
rect 399 465 402 468 
rect 399 468 402 471 
rect 399 471 402 474 
rect 399 474 402 477 
rect 399 477 402 480 
rect 399 480 402 483 
rect 399 483 402 486 
rect 399 486 402 489 
rect 399 489 402 492 
rect 399 492 402 495 
rect 399 495 402 498 
rect 399 498 402 501 
rect 399 501 402 504 
rect 399 504 402 507 
rect 399 507 402 510 
rect 402 0 405 3 
rect 402 3 405 6 
rect 402 6 405 9 
rect 402 9 405 12 
rect 402 12 405 15 
rect 402 15 405 18 
rect 402 18 405 21 
rect 402 21 405 24 
rect 402 24 405 27 
rect 402 27 405 30 
rect 402 30 405 33 
rect 402 33 405 36 
rect 402 36 405 39 
rect 402 39 405 42 
rect 402 42 405 45 
rect 402 45 405 48 
rect 402 48 405 51 
rect 402 51 405 54 
rect 402 54 405 57 
rect 402 57 405 60 
rect 402 60 405 63 
rect 402 63 405 66 
rect 402 66 405 69 
rect 402 69 405 72 
rect 402 72 405 75 
rect 402 75 405 78 
rect 402 78 405 81 
rect 402 81 405 84 
rect 402 84 405 87 
rect 402 87 405 90 
rect 402 90 405 93 
rect 402 93 405 96 
rect 402 96 405 99 
rect 402 99 405 102 
rect 402 102 405 105 
rect 402 105 405 108 
rect 402 108 405 111 
rect 402 111 405 114 
rect 402 114 405 117 
rect 402 117 405 120 
rect 402 120 405 123 
rect 402 123 405 126 
rect 402 126 405 129 
rect 402 129 405 132 
rect 402 132 405 135 
rect 402 135 405 138 
rect 402 138 405 141 
rect 402 141 405 144 
rect 402 144 405 147 
rect 402 147 405 150 
rect 402 150 405 153 
rect 402 153 405 156 
rect 402 156 405 159 
rect 402 159 405 162 
rect 402 162 405 165 
rect 402 165 405 168 
rect 402 168 405 171 
rect 402 171 405 174 
rect 402 174 405 177 
rect 402 177 405 180 
rect 402 180 405 183 
rect 402 183 405 186 
rect 402 186 405 189 
rect 402 189 405 192 
rect 402 192 405 195 
rect 402 195 405 198 
rect 402 198 405 201 
rect 402 201 405 204 
rect 402 204 405 207 
rect 402 207 405 210 
rect 402 210 405 213 
rect 402 213 405 216 
rect 402 216 405 219 
rect 402 219 405 222 
rect 402 222 405 225 
rect 402 225 405 228 
rect 402 228 405 231 
rect 402 231 405 234 
rect 402 234 405 237 
rect 402 237 405 240 
rect 402 240 405 243 
rect 402 243 405 246 
rect 402 246 405 249 
rect 402 249 405 252 
rect 402 252 405 255 
rect 402 255 405 258 
rect 402 258 405 261 
rect 402 261 405 264 
rect 402 264 405 267 
rect 402 267 405 270 
rect 402 270 405 273 
rect 402 273 405 276 
rect 402 276 405 279 
rect 402 279 405 282 
rect 402 282 405 285 
rect 402 285 405 288 
rect 402 288 405 291 
rect 402 291 405 294 
rect 402 294 405 297 
rect 402 297 405 300 
rect 402 300 405 303 
rect 402 303 405 306 
rect 402 306 405 309 
rect 402 309 405 312 
rect 402 312 405 315 
rect 402 315 405 318 
rect 402 318 405 321 
rect 402 321 405 324 
rect 402 324 405 327 
rect 402 327 405 330 
rect 402 330 405 333 
rect 402 333 405 336 
rect 402 336 405 339 
rect 402 339 405 342 
rect 402 342 405 345 
rect 402 345 405 348 
rect 402 348 405 351 
rect 402 351 405 354 
rect 402 354 405 357 
rect 402 357 405 360 
rect 402 360 405 363 
rect 402 363 405 366 
rect 402 366 405 369 
rect 402 369 405 372 
rect 402 372 405 375 
rect 402 375 405 378 
rect 402 378 405 381 
rect 402 381 405 384 
rect 402 384 405 387 
rect 402 387 405 390 
rect 402 390 405 393 
rect 402 393 405 396 
rect 402 396 405 399 
rect 402 399 405 402 
rect 402 402 405 405 
rect 402 405 405 408 
rect 402 408 405 411 
rect 402 411 405 414 
rect 402 414 405 417 
rect 402 417 405 420 
rect 402 420 405 423 
rect 402 423 405 426 
rect 402 426 405 429 
rect 402 429 405 432 
rect 402 432 405 435 
rect 402 435 405 438 
rect 402 438 405 441 
rect 402 441 405 444 
rect 402 444 405 447 
rect 402 447 405 450 
rect 402 450 405 453 
rect 402 453 405 456 
rect 402 456 405 459 
rect 402 459 405 462 
rect 402 462 405 465 
rect 402 465 405 468 
rect 402 468 405 471 
rect 402 471 405 474 
rect 402 474 405 477 
rect 402 477 405 480 
rect 402 480 405 483 
rect 402 483 405 486 
rect 402 486 405 489 
rect 402 489 405 492 
rect 402 492 405 495 
rect 402 495 405 498 
rect 402 498 405 501 
rect 402 501 405 504 
rect 402 504 405 507 
rect 402 507 405 510 
rect 405 0 408 3 
rect 405 3 408 6 
rect 405 6 408 9 
rect 405 9 408 12 
rect 405 12 408 15 
rect 405 15 408 18 
rect 405 18 408 21 
rect 405 21 408 24 
rect 405 24 408 27 
rect 405 27 408 30 
rect 405 30 408 33 
rect 405 33 408 36 
rect 405 36 408 39 
rect 405 39 408 42 
rect 405 42 408 45 
rect 405 45 408 48 
rect 405 48 408 51 
rect 405 51 408 54 
rect 405 54 408 57 
rect 405 57 408 60 
rect 405 60 408 63 
rect 405 63 408 66 
rect 405 66 408 69 
rect 405 69 408 72 
rect 405 72 408 75 
rect 405 75 408 78 
rect 405 78 408 81 
rect 405 81 408 84 
rect 405 84 408 87 
rect 405 87 408 90 
rect 405 90 408 93 
rect 405 93 408 96 
rect 405 96 408 99 
rect 405 99 408 102 
rect 405 102 408 105 
rect 405 105 408 108 
rect 405 108 408 111 
rect 405 111 408 114 
rect 405 114 408 117 
rect 405 117 408 120 
rect 405 120 408 123 
rect 405 123 408 126 
rect 405 126 408 129 
rect 405 129 408 132 
rect 405 132 408 135 
rect 405 135 408 138 
rect 405 138 408 141 
rect 405 141 408 144 
rect 405 144 408 147 
rect 405 147 408 150 
rect 405 150 408 153 
rect 405 153 408 156 
rect 405 156 408 159 
rect 405 159 408 162 
rect 405 162 408 165 
rect 405 165 408 168 
rect 405 168 408 171 
rect 405 171 408 174 
rect 405 174 408 177 
rect 405 177 408 180 
rect 405 180 408 183 
rect 405 183 408 186 
rect 405 186 408 189 
rect 405 189 408 192 
rect 405 192 408 195 
rect 405 195 408 198 
rect 405 198 408 201 
rect 405 201 408 204 
rect 405 204 408 207 
rect 405 207 408 210 
rect 405 210 408 213 
rect 405 213 408 216 
rect 405 216 408 219 
rect 405 219 408 222 
rect 405 222 408 225 
rect 405 225 408 228 
rect 405 228 408 231 
rect 405 231 408 234 
rect 405 234 408 237 
rect 405 237 408 240 
rect 405 240 408 243 
rect 405 243 408 246 
rect 405 246 408 249 
rect 405 249 408 252 
rect 405 252 408 255 
rect 405 255 408 258 
rect 405 258 408 261 
rect 405 261 408 264 
rect 405 264 408 267 
rect 405 267 408 270 
rect 405 270 408 273 
rect 405 273 408 276 
rect 405 276 408 279 
rect 405 279 408 282 
rect 405 282 408 285 
rect 405 285 408 288 
rect 405 288 408 291 
rect 405 291 408 294 
rect 405 294 408 297 
rect 405 297 408 300 
rect 405 300 408 303 
rect 405 303 408 306 
rect 405 306 408 309 
rect 405 309 408 312 
rect 405 312 408 315 
rect 405 315 408 318 
rect 405 318 408 321 
rect 405 321 408 324 
rect 405 324 408 327 
rect 405 327 408 330 
rect 405 330 408 333 
rect 405 333 408 336 
rect 405 336 408 339 
rect 405 339 408 342 
rect 405 342 408 345 
rect 405 345 408 348 
rect 405 348 408 351 
rect 405 351 408 354 
rect 405 354 408 357 
rect 405 357 408 360 
rect 405 360 408 363 
rect 405 363 408 366 
rect 405 366 408 369 
rect 405 369 408 372 
rect 405 372 408 375 
rect 405 375 408 378 
rect 405 378 408 381 
rect 405 381 408 384 
rect 405 384 408 387 
rect 405 387 408 390 
rect 405 390 408 393 
rect 405 393 408 396 
rect 405 396 408 399 
rect 405 399 408 402 
rect 405 402 408 405 
rect 405 405 408 408 
rect 405 408 408 411 
rect 405 411 408 414 
rect 405 414 408 417 
rect 405 417 408 420 
rect 405 420 408 423 
rect 405 423 408 426 
rect 405 426 408 429 
rect 405 429 408 432 
rect 405 432 408 435 
rect 405 435 408 438 
rect 405 438 408 441 
rect 405 441 408 444 
rect 405 444 408 447 
rect 405 447 408 450 
rect 405 450 408 453 
rect 405 453 408 456 
rect 405 456 408 459 
rect 405 459 408 462 
rect 405 462 408 465 
rect 405 465 408 468 
rect 405 468 408 471 
rect 405 471 408 474 
rect 405 474 408 477 
rect 405 477 408 480 
rect 405 480 408 483 
rect 405 483 408 486 
rect 405 486 408 489 
rect 405 489 408 492 
rect 405 492 408 495 
rect 405 495 408 498 
rect 405 498 408 501 
rect 405 501 408 504 
rect 405 504 408 507 
rect 405 507 408 510 
rect 408 0 411 3 
rect 408 3 411 6 
rect 408 6 411 9 
rect 408 9 411 12 
rect 408 12 411 15 
rect 408 15 411 18 
rect 408 18 411 21 
rect 408 21 411 24 
rect 408 24 411 27 
rect 408 27 411 30 
rect 408 30 411 33 
rect 408 33 411 36 
rect 408 36 411 39 
rect 408 39 411 42 
rect 408 42 411 45 
rect 408 45 411 48 
rect 408 48 411 51 
rect 408 51 411 54 
rect 408 54 411 57 
rect 408 57 411 60 
rect 408 60 411 63 
rect 408 63 411 66 
rect 408 66 411 69 
rect 408 69 411 72 
rect 408 72 411 75 
rect 408 75 411 78 
rect 408 78 411 81 
rect 408 81 411 84 
rect 408 84 411 87 
rect 408 87 411 90 
rect 408 90 411 93 
rect 408 93 411 96 
rect 408 96 411 99 
rect 408 99 411 102 
rect 408 102 411 105 
rect 408 105 411 108 
rect 408 108 411 111 
rect 408 111 411 114 
rect 408 114 411 117 
rect 408 117 411 120 
rect 408 120 411 123 
rect 408 123 411 126 
rect 408 126 411 129 
rect 408 129 411 132 
rect 408 132 411 135 
rect 408 135 411 138 
rect 408 138 411 141 
rect 408 141 411 144 
rect 408 144 411 147 
rect 408 147 411 150 
rect 408 150 411 153 
rect 408 153 411 156 
rect 408 156 411 159 
rect 408 159 411 162 
rect 408 162 411 165 
rect 408 165 411 168 
rect 408 168 411 171 
rect 408 171 411 174 
rect 408 174 411 177 
rect 408 177 411 180 
rect 408 180 411 183 
rect 408 183 411 186 
rect 408 186 411 189 
rect 408 189 411 192 
rect 408 192 411 195 
rect 408 195 411 198 
rect 408 198 411 201 
rect 408 201 411 204 
rect 408 204 411 207 
rect 408 207 411 210 
rect 408 210 411 213 
rect 408 213 411 216 
rect 408 216 411 219 
rect 408 219 411 222 
rect 408 222 411 225 
rect 408 225 411 228 
rect 408 228 411 231 
rect 408 231 411 234 
rect 408 234 411 237 
rect 408 237 411 240 
rect 408 240 411 243 
rect 408 243 411 246 
rect 408 246 411 249 
rect 408 249 411 252 
rect 408 252 411 255 
rect 408 255 411 258 
rect 408 258 411 261 
rect 408 261 411 264 
rect 408 264 411 267 
rect 408 267 411 270 
rect 408 270 411 273 
rect 408 273 411 276 
rect 408 276 411 279 
rect 408 279 411 282 
rect 408 282 411 285 
rect 408 285 411 288 
rect 408 288 411 291 
rect 408 291 411 294 
rect 408 294 411 297 
rect 408 297 411 300 
rect 408 300 411 303 
rect 408 303 411 306 
rect 408 306 411 309 
rect 408 309 411 312 
rect 408 312 411 315 
rect 408 315 411 318 
rect 408 318 411 321 
rect 408 321 411 324 
rect 408 324 411 327 
rect 408 327 411 330 
rect 408 330 411 333 
rect 408 333 411 336 
rect 408 336 411 339 
rect 408 339 411 342 
rect 408 342 411 345 
rect 408 345 411 348 
rect 408 348 411 351 
rect 408 351 411 354 
rect 408 354 411 357 
rect 408 357 411 360 
rect 408 360 411 363 
rect 408 363 411 366 
rect 408 366 411 369 
rect 408 369 411 372 
rect 408 372 411 375 
rect 408 375 411 378 
rect 408 378 411 381 
rect 408 381 411 384 
rect 408 384 411 387 
rect 408 387 411 390 
rect 408 390 411 393 
rect 408 393 411 396 
rect 408 396 411 399 
rect 408 399 411 402 
rect 408 402 411 405 
rect 408 405 411 408 
rect 408 408 411 411 
rect 408 411 411 414 
rect 408 414 411 417 
rect 408 417 411 420 
rect 408 420 411 423 
rect 408 423 411 426 
rect 408 426 411 429 
rect 408 429 411 432 
rect 408 432 411 435 
rect 408 435 411 438 
rect 408 438 411 441 
rect 408 441 411 444 
rect 408 444 411 447 
rect 408 447 411 450 
rect 408 450 411 453 
rect 408 453 411 456 
rect 408 456 411 459 
rect 408 459 411 462 
rect 408 462 411 465 
rect 408 465 411 468 
rect 408 468 411 471 
rect 408 471 411 474 
rect 408 474 411 477 
rect 408 477 411 480 
rect 408 480 411 483 
rect 408 483 411 486 
rect 408 486 411 489 
rect 408 489 411 492 
rect 408 492 411 495 
rect 408 495 411 498 
rect 408 498 411 501 
rect 408 501 411 504 
rect 408 504 411 507 
rect 408 507 411 510 
rect 411 0 414 3 
rect 411 3 414 6 
rect 411 6 414 9 
rect 411 9 414 12 
rect 411 12 414 15 
rect 411 15 414 18 
rect 411 18 414 21 
rect 411 21 414 24 
rect 411 24 414 27 
rect 411 27 414 30 
rect 411 30 414 33 
rect 411 33 414 36 
rect 411 36 414 39 
rect 411 39 414 42 
rect 411 42 414 45 
rect 411 45 414 48 
rect 411 48 414 51 
rect 411 51 414 54 
rect 411 54 414 57 
rect 411 57 414 60 
rect 411 60 414 63 
rect 411 63 414 66 
rect 411 66 414 69 
rect 411 69 414 72 
rect 411 72 414 75 
rect 411 75 414 78 
rect 411 78 414 81 
rect 411 81 414 84 
rect 411 84 414 87 
rect 411 87 414 90 
rect 411 90 414 93 
rect 411 93 414 96 
rect 411 96 414 99 
rect 411 99 414 102 
rect 411 102 414 105 
rect 411 105 414 108 
rect 411 108 414 111 
rect 411 111 414 114 
rect 411 114 414 117 
rect 411 117 414 120 
rect 411 120 414 123 
rect 411 123 414 126 
rect 411 126 414 129 
rect 411 129 414 132 
rect 411 132 414 135 
rect 411 135 414 138 
rect 411 138 414 141 
rect 411 141 414 144 
rect 411 144 414 147 
rect 411 147 414 150 
rect 411 150 414 153 
rect 411 153 414 156 
rect 411 156 414 159 
rect 411 159 414 162 
rect 411 162 414 165 
rect 411 165 414 168 
rect 411 168 414 171 
rect 411 171 414 174 
rect 411 174 414 177 
rect 411 177 414 180 
rect 411 180 414 183 
rect 411 183 414 186 
rect 411 186 414 189 
rect 411 189 414 192 
rect 411 192 414 195 
rect 411 195 414 198 
rect 411 198 414 201 
rect 411 201 414 204 
rect 411 204 414 207 
rect 411 207 414 210 
rect 411 210 414 213 
rect 411 213 414 216 
rect 411 216 414 219 
rect 411 219 414 222 
rect 411 222 414 225 
rect 411 225 414 228 
rect 411 228 414 231 
rect 411 231 414 234 
rect 411 234 414 237 
rect 411 237 414 240 
rect 411 240 414 243 
rect 411 243 414 246 
rect 411 246 414 249 
rect 411 249 414 252 
rect 411 252 414 255 
rect 411 255 414 258 
rect 411 258 414 261 
rect 411 261 414 264 
rect 411 264 414 267 
rect 411 267 414 270 
rect 411 270 414 273 
rect 411 273 414 276 
rect 411 276 414 279 
rect 411 279 414 282 
rect 411 282 414 285 
rect 411 285 414 288 
rect 411 288 414 291 
rect 411 291 414 294 
rect 411 294 414 297 
rect 411 297 414 300 
rect 411 300 414 303 
rect 411 303 414 306 
rect 411 306 414 309 
rect 411 309 414 312 
rect 411 312 414 315 
rect 411 315 414 318 
rect 411 318 414 321 
rect 411 321 414 324 
rect 411 324 414 327 
rect 411 327 414 330 
rect 411 330 414 333 
rect 411 333 414 336 
rect 411 336 414 339 
rect 411 339 414 342 
rect 411 342 414 345 
rect 411 345 414 348 
rect 411 348 414 351 
rect 411 351 414 354 
rect 411 354 414 357 
rect 411 357 414 360 
rect 411 360 414 363 
rect 411 363 414 366 
rect 411 366 414 369 
rect 411 369 414 372 
rect 411 372 414 375 
rect 411 375 414 378 
rect 411 378 414 381 
rect 411 381 414 384 
rect 411 384 414 387 
rect 411 387 414 390 
rect 411 390 414 393 
rect 411 393 414 396 
rect 411 396 414 399 
rect 411 399 414 402 
rect 411 402 414 405 
rect 411 405 414 408 
rect 411 408 414 411 
rect 411 411 414 414 
rect 411 414 414 417 
rect 411 417 414 420 
rect 411 420 414 423 
rect 411 423 414 426 
rect 411 426 414 429 
rect 411 429 414 432 
rect 411 432 414 435 
rect 411 435 414 438 
rect 411 438 414 441 
rect 411 441 414 444 
rect 411 444 414 447 
rect 411 447 414 450 
rect 411 450 414 453 
rect 411 453 414 456 
rect 411 456 414 459 
rect 411 459 414 462 
rect 411 462 414 465 
rect 411 465 414 468 
rect 411 468 414 471 
rect 411 471 414 474 
rect 411 474 414 477 
rect 411 477 414 480 
rect 411 480 414 483 
rect 411 483 414 486 
rect 411 486 414 489 
rect 411 489 414 492 
rect 411 492 414 495 
rect 411 495 414 498 
rect 411 498 414 501 
rect 411 501 414 504 
rect 411 504 414 507 
rect 411 507 414 510 
rect 414 0 417 3 
rect 414 3 417 6 
rect 414 6 417 9 
rect 414 9 417 12 
rect 414 12 417 15 
rect 414 15 417 18 
rect 414 18 417 21 
rect 414 21 417 24 
rect 414 24 417 27 
rect 414 27 417 30 
rect 414 30 417 33 
rect 414 33 417 36 
rect 414 36 417 39 
rect 414 39 417 42 
rect 414 42 417 45 
rect 414 45 417 48 
rect 414 48 417 51 
rect 414 51 417 54 
rect 414 54 417 57 
rect 414 57 417 60 
rect 414 60 417 63 
rect 414 63 417 66 
rect 414 66 417 69 
rect 414 69 417 72 
rect 414 72 417 75 
rect 414 75 417 78 
rect 414 78 417 81 
rect 414 81 417 84 
rect 414 84 417 87 
rect 414 87 417 90 
rect 414 90 417 93 
rect 414 93 417 96 
rect 414 96 417 99 
rect 414 99 417 102 
rect 414 102 417 105 
rect 414 105 417 108 
rect 414 108 417 111 
rect 414 111 417 114 
rect 414 114 417 117 
rect 414 117 417 120 
rect 414 120 417 123 
rect 414 123 417 126 
rect 414 126 417 129 
rect 414 129 417 132 
rect 414 132 417 135 
rect 414 135 417 138 
rect 414 138 417 141 
rect 414 141 417 144 
rect 414 144 417 147 
rect 414 147 417 150 
rect 414 150 417 153 
rect 414 153 417 156 
rect 414 156 417 159 
rect 414 159 417 162 
rect 414 162 417 165 
rect 414 165 417 168 
rect 414 168 417 171 
rect 414 171 417 174 
rect 414 174 417 177 
rect 414 177 417 180 
rect 414 180 417 183 
rect 414 183 417 186 
rect 414 186 417 189 
rect 414 189 417 192 
rect 414 192 417 195 
rect 414 195 417 198 
rect 414 198 417 201 
rect 414 201 417 204 
rect 414 204 417 207 
rect 414 207 417 210 
rect 414 210 417 213 
rect 414 213 417 216 
rect 414 216 417 219 
rect 414 219 417 222 
rect 414 222 417 225 
rect 414 225 417 228 
rect 414 228 417 231 
rect 414 231 417 234 
rect 414 234 417 237 
rect 414 237 417 240 
rect 414 240 417 243 
rect 414 243 417 246 
rect 414 246 417 249 
rect 414 249 417 252 
rect 414 252 417 255 
rect 414 255 417 258 
rect 414 258 417 261 
rect 414 261 417 264 
rect 414 264 417 267 
rect 414 267 417 270 
rect 414 270 417 273 
rect 414 273 417 276 
rect 414 276 417 279 
rect 414 279 417 282 
rect 414 282 417 285 
rect 414 285 417 288 
rect 414 288 417 291 
rect 414 291 417 294 
rect 414 294 417 297 
rect 414 297 417 300 
rect 414 300 417 303 
rect 414 303 417 306 
rect 414 306 417 309 
rect 414 309 417 312 
rect 414 312 417 315 
rect 414 315 417 318 
rect 414 318 417 321 
rect 414 321 417 324 
rect 414 324 417 327 
rect 414 327 417 330 
rect 414 330 417 333 
rect 414 333 417 336 
rect 414 336 417 339 
rect 414 339 417 342 
rect 414 342 417 345 
rect 414 345 417 348 
rect 414 348 417 351 
rect 414 351 417 354 
rect 414 354 417 357 
rect 414 357 417 360 
rect 414 360 417 363 
rect 414 363 417 366 
rect 414 366 417 369 
rect 414 369 417 372 
rect 414 372 417 375 
rect 414 375 417 378 
rect 414 378 417 381 
rect 414 381 417 384 
rect 414 384 417 387 
rect 414 387 417 390 
rect 414 390 417 393 
rect 414 393 417 396 
rect 414 396 417 399 
rect 414 399 417 402 
rect 414 402 417 405 
rect 414 405 417 408 
rect 414 408 417 411 
rect 414 411 417 414 
rect 414 414 417 417 
rect 414 417 417 420 
rect 414 420 417 423 
rect 414 423 417 426 
rect 414 426 417 429 
rect 414 429 417 432 
rect 414 432 417 435 
rect 414 435 417 438 
rect 414 438 417 441 
rect 414 441 417 444 
rect 414 444 417 447 
rect 414 447 417 450 
rect 414 450 417 453 
rect 414 453 417 456 
rect 414 456 417 459 
rect 414 459 417 462 
rect 414 462 417 465 
rect 414 465 417 468 
rect 414 468 417 471 
rect 414 471 417 474 
rect 414 474 417 477 
rect 414 477 417 480 
rect 414 480 417 483 
rect 414 483 417 486 
rect 414 486 417 489 
rect 414 489 417 492 
rect 414 492 417 495 
rect 414 495 417 498 
rect 414 498 417 501 
rect 414 501 417 504 
rect 414 504 417 507 
rect 414 507 417 510 
rect 417 0 420 3 
rect 417 3 420 6 
rect 417 6 420 9 
rect 417 9 420 12 
rect 417 12 420 15 
rect 417 15 420 18 
rect 417 18 420 21 
rect 417 21 420 24 
rect 417 24 420 27 
rect 417 27 420 30 
rect 417 30 420 33 
rect 417 33 420 36 
rect 417 36 420 39 
rect 417 39 420 42 
rect 417 42 420 45 
rect 417 45 420 48 
rect 417 48 420 51 
rect 417 51 420 54 
rect 417 54 420 57 
rect 417 57 420 60 
rect 417 60 420 63 
rect 417 63 420 66 
rect 417 66 420 69 
rect 417 69 420 72 
rect 417 72 420 75 
rect 417 75 420 78 
rect 417 78 420 81 
rect 417 81 420 84 
rect 417 84 420 87 
rect 417 87 420 90 
rect 417 90 420 93 
rect 417 93 420 96 
rect 417 96 420 99 
rect 417 99 420 102 
rect 417 102 420 105 
rect 417 105 420 108 
rect 417 108 420 111 
rect 417 111 420 114 
rect 417 114 420 117 
rect 417 117 420 120 
rect 417 120 420 123 
rect 417 123 420 126 
rect 417 126 420 129 
rect 417 129 420 132 
rect 417 132 420 135 
rect 417 135 420 138 
rect 417 138 420 141 
rect 417 141 420 144 
rect 417 144 420 147 
rect 417 147 420 150 
rect 417 150 420 153 
rect 417 153 420 156 
rect 417 156 420 159 
rect 417 159 420 162 
rect 417 162 420 165 
rect 417 165 420 168 
rect 417 168 420 171 
rect 417 171 420 174 
rect 417 174 420 177 
rect 417 177 420 180 
rect 417 180 420 183 
rect 417 183 420 186 
rect 417 186 420 189 
rect 417 189 420 192 
rect 417 192 420 195 
rect 417 195 420 198 
rect 417 198 420 201 
rect 417 201 420 204 
rect 417 204 420 207 
rect 417 207 420 210 
rect 417 210 420 213 
rect 417 213 420 216 
rect 417 216 420 219 
rect 417 219 420 222 
rect 417 222 420 225 
rect 417 225 420 228 
rect 417 228 420 231 
rect 417 231 420 234 
rect 417 234 420 237 
rect 417 237 420 240 
rect 417 240 420 243 
rect 417 243 420 246 
rect 417 246 420 249 
rect 417 249 420 252 
rect 417 252 420 255 
rect 417 255 420 258 
rect 417 258 420 261 
rect 417 261 420 264 
rect 417 264 420 267 
rect 417 267 420 270 
rect 417 270 420 273 
rect 417 273 420 276 
rect 417 276 420 279 
rect 417 279 420 282 
rect 417 282 420 285 
rect 417 285 420 288 
rect 417 288 420 291 
rect 417 291 420 294 
rect 417 294 420 297 
rect 417 297 420 300 
rect 417 300 420 303 
rect 417 303 420 306 
rect 417 306 420 309 
rect 417 309 420 312 
rect 417 312 420 315 
rect 417 315 420 318 
rect 417 318 420 321 
rect 417 321 420 324 
rect 417 324 420 327 
rect 417 327 420 330 
rect 417 330 420 333 
rect 417 333 420 336 
rect 417 336 420 339 
rect 417 339 420 342 
rect 417 342 420 345 
rect 417 345 420 348 
rect 417 348 420 351 
rect 417 351 420 354 
rect 417 354 420 357 
rect 417 357 420 360 
rect 417 360 420 363 
rect 417 363 420 366 
rect 417 366 420 369 
rect 417 369 420 372 
rect 417 372 420 375 
rect 417 375 420 378 
rect 417 378 420 381 
rect 417 381 420 384 
rect 417 384 420 387 
rect 417 387 420 390 
rect 417 390 420 393 
rect 417 393 420 396 
rect 417 396 420 399 
rect 417 399 420 402 
rect 417 402 420 405 
rect 417 405 420 408 
rect 417 408 420 411 
rect 417 411 420 414 
rect 417 414 420 417 
rect 417 417 420 420 
rect 417 420 420 423 
rect 417 423 420 426 
rect 417 426 420 429 
rect 417 429 420 432 
rect 417 432 420 435 
rect 417 435 420 438 
rect 417 438 420 441 
rect 417 441 420 444 
rect 417 444 420 447 
rect 417 447 420 450 
rect 417 450 420 453 
rect 417 453 420 456 
rect 417 456 420 459 
rect 417 459 420 462 
rect 417 462 420 465 
rect 417 465 420 468 
rect 417 468 420 471 
rect 417 471 420 474 
rect 417 474 420 477 
rect 417 477 420 480 
rect 417 480 420 483 
rect 417 483 420 486 
rect 417 486 420 489 
rect 417 489 420 492 
rect 417 492 420 495 
rect 417 495 420 498 
rect 417 498 420 501 
rect 417 501 420 504 
rect 417 504 420 507 
rect 417 507 420 510 
rect 420 0 423 3 
rect 420 3 423 6 
rect 420 6 423 9 
rect 420 9 423 12 
rect 420 12 423 15 
rect 420 15 423 18 
rect 420 18 423 21 
rect 420 21 423 24 
rect 420 24 423 27 
rect 420 27 423 30 
rect 420 30 423 33 
rect 420 33 423 36 
rect 420 36 423 39 
rect 420 39 423 42 
rect 420 42 423 45 
rect 420 45 423 48 
rect 420 48 423 51 
rect 420 51 423 54 
rect 420 54 423 57 
rect 420 57 423 60 
rect 420 60 423 63 
rect 420 63 423 66 
rect 420 66 423 69 
rect 420 69 423 72 
rect 420 72 423 75 
rect 420 75 423 78 
rect 420 78 423 81 
rect 420 81 423 84 
rect 420 84 423 87 
rect 420 87 423 90 
rect 420 90 423 93 
rect 420 93 423 96 
rect 420 96 423 99 
rect 420 99 423 102 
rect 420 102 423 105 
rect 420 105 423 108 
rect 420 108 423 111 
rect 420 111 423 114 
rect 420 114 423 117 
rect 420 117 423 120 
rect 420 120 423 123 
rect 420 123 423 126 
rect 420 126 423 129 
rect 420 129 423 132 
rect 420 132 423 135 
rect 420 135 423 138 
rect 420 138 423 141 
rect 420 141 423 144 
rect 420 144 423 147 
rect 420 147 423 150 
rect 420 150 423 153 
rect 420 153 423 156 
rect 420 156 423 159 
rect 420 159 423 162 
rect 420 162 423 165 
rect 420 165 423 168 
rect 420 168 423 171 
rect 420 171 423 174 
rect 420 174 423 177 
rect 420 177 423 180 
rect 420 180 423 183 
rect 420 183 423 186 
rect 420 186 423 189 
rect 420 189 423 192 
rect 420 192 423 195 
rect 420 195 423 198 
rect 420 198 423 201 
rect 420 201 423 204 
rect 420 204 423 207 
rect 420 207 423 210 
rect 420 210 423 213 
rect 420 213 423 216 
rect 420 216 423 219 
rect 420 219 423 222 
rect 420 222 423 225 
rect 420 225 423 228 
rect 420 228 423 231 
rect 420 231 423 234 
rect 420 234 423 237 
rect 420 237 423 240 
rect 420 240 423 243 
rect 420 243 423 246 
rect 420 246 423 249 
rect 420 249 423 252 
rect 420 252 423 255 
rect 420 255 423 258 
rect 420 258 423 261 
rect 420 261 423 264 
rect 420 264 423 267 
rect 420 267 423 270 
rect 420 270 423 273 
rect 420 273 423 276 
rect 420 276 423 279 
rect 420 279 423 282 
rect 420 282 423 285 
rect 420 285 423 288 
rect 420 288 423 291 
rect 420 291 423 294 
rect 420 294 423 297 
rect 420 297 423 300 
rect 420 300 423 303 
rect 420 303 423 306 
rect 420 306 423 309 
rect 420 309 423 312 
rect 420 312 423 315 
rect 420 315 423 318 
rect 420 318 423 321 
rect 420 321 423 324 
rect 420 324 423 327 
rect 420 327 423 330 
rect 420 330 423 333 
rect 420 333 423 336 
rect 420 336 423 339 
rect 420 339 423 342 
rect 420 342 423 345 
rect 420 345 423 348 
rect 420 348 423 351 
rect 420 351 423 354 
rect 420 354 423 357 
rect 420 357 423 360 
rect 420 360 423 363 
rect 420 363 423 366 
rect 420 366 423 369 
rect 420 369 423 372 
rect 420 372 423 375 
rect 420 375 423 378 
rect 420 378 423 381 
rect 420 381 423 384 
rect 420 384 423 387 
rect 420 387 423 390 
rect 420 390 423 393 
rect 420 393 423 396 
rect 420 396 423 399 
rect 420 399 423 402 
rect 420 402 423 405 
rect 420 405 423 408 
rect 420 408 423 411 
rect 420 411 423 414 
rect 420 414 423 417 
rect 420 417 423 420 
rect 420 420 423 423 
rect 420 423 423 426 
rect 420 426 423 429 
rect 420 429 423 432 
rect 420 432 423 435 
rect 420 435 423 438 
rect 420 438 423 441 
rect 420 441 423 444 
rect 420 444 423 447 
rect 420 447 423 450 
rect 420 450 423 453 
rect 420 453 423 456 
rect 420 456 423 459 
rect 420 459 423 462 
rect 420 462 423 465 
rect 420 465 423 468 
rect 420 468 423 471 
rect 420 471 423 474 
rect 420 474 423 477 
rect 420 477 423 480 
rect 420 480 423 483 
rect 420 483 423 486 
rect 420 486 423 489 
rect 420 489 423 492 
rect 420 492 423 495 
rect 420 495 423 498 
rect 420 498 423 501 
rect 420 501 423 504 
rect 420 504 423 507 
rect 420 507 423 510 
rect 423 0 426 3 
rect 423 3 426 6 
rect 423 6 426 9 
rect 423 9 426 12 
rect 423 12 426 15 
rect 423 15 426 18 
rect 423 18 426 21 
rect 423 21 426 24 
rect 423 24 426 27 
rect 423 27 426 30 
rect 423 30 426 33 
rect 423 33 426 36 
rect 423 36 426 39 
rect 423 39 426 42 
rect 423 42 426 45 
rect 423 45 426 48 
rect 423 48 426 51 
rect 423 51 426 54 
rect 423 54 426 57 
rect 423 57 426 60 
rect 423 60 426 63 
rect 423 63 426 66 
rect 423 66 426 69 
rect 423 69 426 72 
rect 423 72 426 75 
rect 423 75 426 78 
rect 423 78 426 81 
rect 423 81 426 84 
rect 423 84 426 87 
rect 423 87 426 90 
rect 423 90 426 93 
rect 423 93 426 96 
rect 423 96 426 99 
rect 423 99 426 102 
rect 423 102 426 105 
rect 423 105 426 108 
rect 423 108 426 111 
rect 423 111 426 114 
rect 423 114 426 117 
rect 423 117 426 120 
rect 423 120 426 123 
rect 423 123 426 126 
rect 423 126 426 129 
rect 423 129 426 132 
rect 423 132 426 135 
rect 423 135 426 138 
rect 423 138 426 141 
rect 423 141 426 144 
rect 423 144 426 147 
rect 423 147 426 150 
rect 423 150 426 153 
rect 423 153 426 156 
rect 423 156 426 159 
rect 423 159 426 162 
rect 423 162 426 165 
rect 423 165 426 168 
rect 423 168 426 171 
rect 423 171 426 174 
rect 423 174 426 177 
rect 423 177 426 180 
rect 423 180 426 183 
rect 423 183 426 186 
rect 423 186 426 189 
rect 423 189 426 192 
rect 423 192 426 195 
rect 423 195 426 198 
rect 423 198 426 201 
rect 423 201 426 204 
rect 423 204 426 207 
rect 423 207 426 210 
rect 423 210 426 213 
rect 423 213 426 216 
rect 423 216 426 219 
rect 423 219 426 222 
rect 423 222 426 225 
rect 423 225 426 228 
rect 423 228 426 231 
rect 423 231 426 234 
rect 423 234 426 237 
rect 423 237 426 240 
rect 423 240 426 243 
rect 423 243 426 246 
rect 423 246 426 249 
rect 423 249 426 252 
rect 423 252 426 255 
rect 423 255 426 258 
rect 423 258 426 261 
rect 423 261 426 264 
rect 423 264 426 267 
rect 423 267 426 270 
rect 423 270 426 273 
rect 423 273 426 276 
rect 423 276 426 279 
rect 423 279 426 282 
rect 423 282 426 285 
rect 423 285 426 288 
rect 423 288 426 291 
rect 423 291 426 294 
rect 423 294 426 297 
rect 423 297 426 300 
rect 423 300 426 303 
rect 423 303 426 306 
rect 423 306 426 309 
rect 423 309 426 312 
rect 423 312 426 315 
rect 423 315 426 318 
rect 423 318 426 321 
rect 423 321 426 324 
rect 423 324 426 327 
rect 423 327 426 330 
rect 423 330 426 333 
rect 423 333 426 336 
rect 423 336 426 339 
rect 423 339 426 342 
rect 423 342 426 345 
rect 423 345 426 348 
rect 423 348 426 351 
rect 423 351 426 354 
rect 423 354 426 357 
rect 423 357 426 360 
rect 423 360 426 363 
rect 423 363 426 366 
rect 423 366 426 369 
rect 423 369 426 372 
rect 423 372 426 375 
rect 423 375 426 378 
rect 423 378 426 381 
rect 423 381 426 384 
rect 423 384 426 387 
rect 423 387 426 390 
rect 423 390 426 393 
rect 423 393 426 396 
rect 423 396 426 399 
rect 423 399 426 402 
rect 423 402 426 405 
rect 423 405 426 408 
rect 423 408 426 411 
rect 423 411 426 414 
rect 423 414 426 417 
rect 423 417 426 420 
rect 423 420 426 423 
rect 423 423 426 426 
rect 423 426 426 429 
rect 423 429 426 432 
rect 423 432 426 435 
rect 423 435 426 438 
rect 423 438 426 441 
rect 423 441 426 444 
rect 423 444 426 447 
rect 423 447 426 450 
rect 423 450 426 453 
rect 423 453 426 456 
rect 423 456 426 459 
rect 423 459 426 462 
rect 423 462 426 465 
rect 423 465 426 468 
rect 423 468 426 471 
rect 423 471 426 474 
rect 423 474 426 477 
rect 423 477 426 480 
rect 423 480 426 483 
rect 423 483 426 486 
rect 423 486 426 489 
rect 423 489 426 492 
rect 423 492 426 495 
rect 423 495 426 498 
rect 423 498 426 501 
rect 423 501 426 504 
rect 423 504 426 507 
rect 423 507 426 510 
rect 426 0 429 3 
rect 426 3 429 6 
rect 426 6 429 9 
rect 426 9 429 12 
rect 426 12 429 15 
rect 426 15 429 18 
rect 426 18 429 21 
rect 426 21 429 24 
rect 426 24 429 27 
rect 426 27 429 30 
rect 426 30 429 33 
rect 426 33 429 36 
rect 426 36 429 39 
rect 426 39 429 42 
rect 426 42 429 45 
rect 426 45 429 48 
rect 426 48 429 51 
rect 426 51 429 54 
rect 426 54 429 57 
rect 426 57 429 60 
rect 426 60 429 63 
rect 426 63 429 66 
rect 426 66 429 69 
rect 426 69 429 72 
rect 426 72 429 75 
rect 426 75 429 78 
rect 426 78 429 81 
rect 426 81 429 84 
rect 426 84 429 87 
rect 426 87 429 90 
rect 426 90 429 93 
rect 426 93 429 96 
rect 426 96 429 99 
rect 426 99 429 102 
rect 426 102 429 105 
rect 426 105 429 108 
rect 426 108 429 111 
rect 426 111 429 114 
rect 426 114 429 117 
rect 426 117 429 120 
rect 426 120 429 123 
rect 426 123 429 126 
rect 426 126 429 129 
rect 426 129 429 132 
rect 426 132 429 135 
rect 426 135 429 138 
rect 426 138 429 141 
rect 426 141 429 144 
rect 426 144 429 147 
rect 426 147 429 150 
rect 426 150 429 153 
rect 426 153 429 156 
rect 426 156 429 159 
rect 426 159 429 162 
rect 426 162 429 165 
rect 426 165 429 168 
rect 426 168 429 171 
rect 426 171 429 174 
rect 426 174 429 177 
rect 426 177 429 180 
rect 426 180 429 183 
rect 426 183 429 186 
rect 426 186 429 189 
rect 426 189 429 192 
rect 426 192 429 195 
rect 426 195 429 198 
rect 426 198 429 201 
rect 426 201 429 204 
rect 426 204 429 207 
rect 426 207 429 210 
rect 426 210 429 213 
rect 426 213 429 216 
rect 426 216 429 219 
rect 426 219 429 222 
rect 426 222 429 225 
rect 426 225 429 228 
rect 426 228 429 231 
rect 426 231 429 234 
rect 426 234 429 237 
rect 426 237 429 240 
rect 426 240 429 243 
rect 426 243 429 246 
rect 426 246 429 249 
rect 426 249 429 252 
rect 426 252 429 255 
rect 426 255 429 258 
rect 426 258 429 261 
rect 426 261 429 264 
rect 426 264 429 267 
rect 426 267 429 270 
rect 426 270 429 273 
rect 426 273 429 276 
rect 426 276 429 279 
rect 426 279 429 282 
rect 426 282 429 285 
rect 426 285 429 288 
rect 426 288 429 291 
rect 426 291 429 294 
rect 426 294 429 297 
rect 426 297 429 300 
rect 426 300 429 303 
rect 426 303 429 306 
rect 426 306 429 309 
rect 426 309 429 312 
rect 426 312 429 315 
rect 426 315 429 318 
rect 426 318 429 321 
rect 426 321 429 324 
rect 426 324 429 327 
rect 426 327 429 330 
rect 426 330 429 333 
rect 426 333 429 336 
rect 426 336 429 339 
rect 426 339 429 342 
rect 426 342 429 345 
rect 426 345 429 348 
rect 426 348 429 351 
rect 426 351 429 354 
rect 426 354 429 357 
rect 426 357 429 360 
rect 426 360 429 363 
rect 426 363 429 366 
rect 426 366 429 369 
rect 426 369 429 372 
rect 426 372 429 375 
rect 426 375 429 378 
rect 426 378 429 381 
rect 426 381 429 384 
rect 426 384 429 387 
rect 426 387 429 390 
rect 426 390 429 393 
rect 426 393 429 396 
rect 426 396 429 399 
rect 426 399 429 402 
rect 426 402 429 405 
rect 426 405 429 408 
rect 426 408 429 411 
rect 426 411 429 414 
rect 426 414 429 417 
rect 426 417 429 420 
rect 426 420 429 423 
rect 426 423 429 426 
rect 426 426 429 429 
rect 426 429 429 432 
rect 426 432 429 435 
rect 426 435 429 438 
rect 426 438 429 441 
rect 426 441 429 444 
rect 426 444 429 447 
rect 426 447 429 450 
rect 426 450 429 453 
rect 426 453 429 456 
rect 426 456 429 459 
rect 426 459 429 462 
rect 426 462 429 465 
rect 426 465 429 468 
rect 426 468 429 471 
rect 426 471 429 474 
rect 426 474 429 477 
rect 426 477 429 480 
rect 426 480 429 483 
rect 426 483 429 486 
rect 426 486 429 489 
rect 426 489 429 492 
rect 426 492 429 495 
rect 426 495 429 498 
rect 426 498 429 501 
rect 426 501 429 504 
rect 426 504 429 507 
rect 426 507 429 510 
rect 429 0 432 3 
rect 429 3 432 6 
rect 429 6 432 9 
rect 429 9 432 12 
rect 429 12 432 15 
rect 429 15 432 18 
rect 429 18 432 21 
rect 429 21 432 24 
rect 429 24 432 27 
rect 429 27 432 30 
rect 429 30 432 33 
rect 429 33 432 36 
rect 429 36 432 39 
rect 429 39 432 42 
rect 429 42 432 45 
rect 429 45 432 48 
rect 429 48 432 51 
rect 429 51 432 54 
rect 429 54 432 57 
rect 429 57 432 60 
rect 429 60 432 63 
rect 429 63 432 66 
rect 429 66 432 69 
rect 429 69 432 72 
rect 429 72 432 75 
rect 429 75 432 78 
rect 429 78 432 81 
rect 429 81 432 84 
rect 429 84 432 87 
rect 429 87 432 90 
rect 429 90 432 93 
rect 429 93 432 96 
rect 429 96 432 99 
rect 429 99 432 102 
rect 429 102 432 105 
rect 429 105 432 108 
rect 429 108 432 111 
rect 429 111 432 114 
rect 429 114 432 117 
rect 429 117 432 120 
rect 429 120 432 123 
rect 429 123 432 126 
rect 429 126 432 129 
rect 429 129 432 132 
rect 429 132 432 135 
rect 429 135 432 138 
rect 429 138 432 141 
rect 429 141 432 144 
rect 429 144 432 147 
rect 429 147 432 150 
rect 429 150 432 153 
rect 429 153 432 156 
rect 429 156 432 159 
rect 429 159 432 162 
rect 429 162 432 165 
rect 429 165 432 168 
rect 429 168 432 171 
rect 429 171 432 174 
rect 429 174 432 177 
rect 429 177 432 180 
rect 429 180 432 183 
rect 429 183 432 186 
rect 429 186 432 189 
rect 429 189 432 192 
rect 429 192 432 195 
rect 429 195 432 198 
rect 429 198 432 201 
rect 429 201 432 204 
rect 429 204 432 207 
rect 429 207 432 210 
rect 429 210 432 213 
rect 429 213 432 216 
rect 429 216 432 219 
rect 429 219 432 222 
rect 429 222 432 225 
rect 429 225 432 228 
rect 429 228 432 231 
rect 429 231 432 234 
rect 429 234 432 237 
rect 429 237 432 240 
rect 429 240 432 243 
rect 429 243 432 246 
rect 429 246 432 249 
rect 429 249 432 252 
rect 429 252 432 255 
rect 429 255 432 258 
rect 429 258 432 261 
rect 429 261 432 264 
rect 429 264 432 267 
rect 429 267 432 270 
rect 429 270 432 273 
rect 429 273 432 276 
rect 429 276 432 279 
rect 429 279 432 282 
rect 429 282 432 285 
rect 429 285 432 288 
rect 429 288 432 291 
rect 429 291 432 294 
rect 429 294 432 297 
rect 429 297 432 300 
rect 429 300 432 303 
rect 429 303 432 306 
rect 429 306 432 309 
rect 429 309 432 312 
rect 429 312 432 315 
rect 429 315 432 318 
rect 429 318 432 321 
rect 429 321 432 324 
rect 429 324 432 327 
rect 429 327 432 330 
rect 429 330 432 333 
rect 429 333 432 336 
rect 429 336 432 339 
rect 429 339 432 342 
rect 429 342 432 345 
rect 429 345 432 348 
rect 429 348 432 351 
rect 429 351 432 354 
rect 429 354 432 357 
rect 429 357 432 360 
rect 429 360 432 363 
rect 429 363 432 366 
rect 429 366 432 369 
rect 429 369 432 372 
rect 429 372 432 375 
rect 429 375 432 378 
rect 429 378 432 381 
rect 429 381 432 384 
rect 429 384 432 387 
rect 429 387 432 390 
rect 429 390 432 393 
rect 429 393 432 396 
rect 429 396 432 399 
rect 429 399 432 402 
rect 429 402 432 405 
rect 429 405 432 408 
rect 429 408 432 411 
rect 429 411 432 414 
rect 429 414 432 417 
rect 429 417 432 420 
rect 429 420 432 423 
rect 429 423 432 426 
rect 429 426 432 429 
rect 429 429 432 432 
rect 429 432 432 435 
rect 429 435 432 438 
rect 429 438 432 441 
rect 429 441 432 444 
rect 429 444 432 447 
rect 429 447 432 450 
rect 429 450 432 453 
rect 429 453 432 456 
rect 429 456 432 459 
rect 429 459 432 462 
rect 429 462 432 465 
rect 429 465 432 468 
rect 429 468 432 471 
rect 429 471 432 474 
rect 429 474 432 477 
rect 429 477 432 480 
rect 429 480 432 483 
rect 429 483 432 486 
rect 429 486 432 489 
rect 429 489 432 492 
rect 429 492 432 495 
rect 429 495 432 498 
rect 429 498 432 501 
rect 429 501 432 504 
rect 429 504 432 507 
rect 429 507 432 510 
rect 432 0 435 3 
rect 432 3 435 6 
rect 432 6 435 9 
rect 432 9 435 12 
rect 432 12 435 15 
rect 432 15 435 18 
rect 432 18 435 21 
rect 432 21 435 24 
rect 432 24 435 27 
rect 432 27 435 30 
rect 432 30 435 33 
rect 432 33 435 36 
rect 432 36 435 39 
rect 432 39 435 42 
rect 432 42 435 45 
rect 432 45 435 48 
rect 432 48 435 51 
rect 432 51 435 54 
rect 432 54 435 57 
rect 432 57 435 60 
rect 432 60 435 63 
rect 432 63 435 66 
rect 432 66 435 69 
rect 432 69 435 72 
rect 432 72 435 75 
rect 432 75 435 78 
rect 432 78 435 81 
rect 432 81 435 84 
rect 432 84 435 87 
rect 432 87 435 90 
rect 432 90 435 93 
rect 432 93 435 96 
rect 432 96 435 99 
rect 432 99 435 102 
rect 432 102 435 105 
rect 432 105 435 108 
rect 432 108 435 111 
rect 432 111 435 114 
rect 432 114 435 117 
rect 432 117 435 120 
rect 432 120 435 123 
rect 432 123 435 126 
rect 432 126 435 129 
rect 432 129 435 132 
rect 432 132 435 135 
rect 432 135 435 138 
rect 432 138 435 141 
rect 432 141 435 144 
rect 432 144 435 147 
rect 432 147 435 150 
rect 432 150 435 153 
rect 432 153 435 156 
rect 432 156 435 159 
rect 432 159 435 162 
rect 432 162 435 165 
rect 432 165 435 168 
rect 432 168 435 171 
rect 432 171 435 174 
rect 432 174 435 177 
rect 432 177 435 180 
rect 432 180 435 183 
rect 432 183 435 186 
rect 432 186 435 189 
rect 432 189 435 192 
rect 432 192 435 195 
rect 432 195 435 198 
rect 432 198 435 201 
rect 432 201 435 204 
rect 432 204 435 207 
rect 432 207 435 210 
rect 432 210 435 213 
rect 432 213 435 216 
rect 432 216 435 219 
rect 432 219 435 222 
rect 432 222 435 225 
rect 432 225 435 228 
rect 432 228 435 231 
rect 432 231 435 234 
rect 432 234 435 237 
rect 432 237 435 240 
rect 432 240 435 243 
rect 432 243 435 246 
rect 432 246 435 249 
rect 432 249 435 252 
rect 432 252 435 255 
rect 432 255 435 258 
rect 432 258 435 261 
rect 432 261 435 264 
rect 432 264 435 267 
rect 432 267 435 270 
rect 432 270 435 273 
rect 432 273 435 276 
rect 432 276 435 279 
rect 432 279 435 282 
rect 432 282 435 285 
rect 432 285 435 288 
rect 432 288 435 291 
rect 432 291 435 294 
rect 432 294 435 297 
rect 432 297 435 300 
rect 432 300 435 303 
rect 432 303 435 306 
rect 432 306 435 309 
rect 432 309 435 312 
rect 432 312 435 315 
rect 432 315 435 318 
rect 432 318 435 321 
rect 432 321 435 324 
rect 432 324 435 327 
rect 432 327 435 330 
rect 432 330 435 333 
rect 432 333 435 336 
rect 432 336 435 339 
rect 432 339 435 342 
rect 432 342 435 345 
rect 432 345 435 348 
rect 432 348 435 351 
rect 432 351 435 354 
rect 432 354 435 357 
rect 432 357 435 360 
rect 432 360 435 363 
rect 432 363 435 366 
rect 432 366 435 369 
rect 432 369 435 372 
rect 432 372 435 375 
rect 432 375 435 378 
rect 432 378 435 381 
rect 432 381 435 384 
rect 432 384 435 387 
rect 432 387 435 390 
rect 432 390 435 393 
rect 432 393 435 396 
rect 432 396 435 399 
rect 432 399 435 402 
rect 432 402 435 405 
rect 432 405 435 408 
rect 432 408 435 411 
rect 432 411 435 414 
rect 432 414 435 417 
rect 432 417 435 420 
rect 432 420 435 423 
rect 432 423 435 426 
rect 432 426 435 429 
rect 432 429 435 432 
rect 432 432 435 435 
rect 432 435 435 438 
rect 432 438 435 441 
rect 432 441 435 444 
rect 432 444 435 447 
rect 432 447 435 450 
rect 432 450 435 453 
rect 432 453 435 456 
rect 432 456 435 459 
rect 432 459 435 462 
rect 432 462 435 465 
rect 432 465 435 468 
rect 432 468 435 471 
rect 432 471 435 474 
rect 432 474 435 477 
rect 432 477 435 480 
rect 432 480 435 483 
rect 432 483 435 486 
rect 432 486 435 489 
rect 432 489 435 492 
rect 432 492 435 495 
rect 432 495 435 498 
rect 432 498 435 501 
rect 432 501 435 504 
rect 432 504 435 507 
rect 432 507 435 510 
rect 435 0 438 3 
rect 435 3 438 6 
rect 435 6 438 9 
rect 435 9 438 12 
rect 435 12 438 15 
rect 435 15 438 18 
rect 435 18 438 21 
rect 435 21 438 24 
rect 435 24 438 27 
rect 435 27 438 30 
rect 435 30 438 33 
rect 435 33 438 36 
rect 435 36 438 39 
rect 435 39 438 42 
rect 435 42 438 45 
rect 435 45 438 48 
rect 435 48 438 51 
rect 435 51 438 54 
rect 435 54 438 57 
rect 435 57 438 60 
rect 435 60 438 63 
rect 435 63 438 66 
rect 435 66 438 69 
rect 435 69 438 72 
rect 435 72 438 75 
rect 435 75 438 78 
rect 435 78 438 81 
rect 435 81 438 84 
rect 435 84 438 87 
rect 435 87 438 90 
rect 435 90 438 93 
rect 435 93 438 96 
rect 435 96 438 99 
rect 435 99 438 102 
rect 435 102 438 105 
rect 435 105 438 108 
rect 435 108 438 111 
rect 435 111 438 114 
rect 435 114 438 117 
rect 435 117 438 120 
rect 435 120 438 123 
rect 435 123 438 126 
rect 435 126 438 129 
rect 435 129 438 132 
rect 435 132 438 135 
rect 435 135 438 138 
rect 435 138 438 141 
rect 435 141 438 144 
rect 435 144 438 147 
rect 435 147 438 150 
rect 435 150 438 153 
rect 435 153 438 156 
rect 435 156 438 159 
rect 435 159 438 162 
rect 435 162 438 165 
rect 435 165 438 168 
rect 435 168 438 171 
rect 435 171 438 174 
rect 435 174 438 177 
rect 435 177 438 180 
rect 435 180 438 183 
rect 435 183 438 186 
rect 435 186 438 189 
rect 435 189 438 192 
rect 435 192 438 195 
rect 435 195 438 198 
rect 435 198 438 201 
rect 435 201 438 204 
rect 435 204 438 207 
rect 435 207 438 210 
rect 435 210 438 213 
rect 435 213 438 216 
rect 435 216 438 219 
rect 435 219 438 222 
rect 435 222 438 225 
rect 435 225 438 228 
rect 435 228 438 231 
rect 435 231 438 234 
rect 435 234 438 237 
rect 435 237 438 240 
rect 435 240 438 243 
rect 435 243 438 246 
rect 435 246 438 249 
rect 435 249 438 252 
rect 435 252 438 255 
rect 435 255 438 258 
rect 435 258 438 261 
rect 435 261 438 264 
rect 435 264 438 267 
rect 435 267 438 270 
rect 435 270 438 273 
rect 435 273 438 276 
rect 435 276 438 279 
rect 435 279 438 282 
rect 435 282 438 285 
rect 435 285 438 288 
rect 435 288 438 291 
rect 435 291 438 294 
rect 435 294 438 297 
rect 435 297 438 300 
rect 435 300 438 303 
rect 435 303 438 306 
rect 435 306 438 309 
rect 435 309 438 312 
rect 435 312 438 315 
rect 435 315 438 318 
rect 435 318 438 321 
rect 435 321 438 324 
rect 435 324 438 327 
rect 435 327 438 330 
rect 435 330 438 333 
rect 435 333 438 336 
rect 435 336 438 339 
rect 435 339 438 342 
rect 435 342 438 345 
rect 435 345 438 348 
rect 435 348 438 351 
rect 435 351 438 354 
rect 435 354 438 357 
rect 435 357 438 360 
rect 435 360 438 363 
rect 435 363 438 366 
rect 435 366 438 369 
rect 435 369 438 372 
rect 435 372 438 375 
rect 435 375 438 378 
rect 435 378 438 381 
rect 435 381 438 384 
rect 435 384 438 387 
rect 435 387 438 390 
rect 435 390 438 393 
rect 435 393 438 396 
rect 435 396 438 399 
rect 435 399 438 402 
rect 435 402 438 405 
rect 435 405 438 408 
rect 435 408 438 411 
rect 435 411 438 414 
rect 435 414 438 417 
rect 435 417 438 420 
rect 435 420 438 423 
rect 435 423 438 426 
rect 435 426 438 429 
rect 435 429 438 432 
rect 435 432 438 435 
rect 435 435 438 438 
rect 435 438 438 441 
rect 435 441 438 444 
rect 435 444 438 447 
rect 435 447 438 450 
rect 435 450 438 453 
rect 435 453 438 456 
rect 435 456 438 459 
rect 435 459 438 462 
rect 435 462 438 465 
rect 435 465 438 468 
rect 435 468 438 471 
rect 435 471 438 474 
rect 435 474 438 477 
rect 435 477 438 480 
rect 435 480 438 483 
rect 435 483 438 486 
rect 435 486 438 489 
rect 435 489 438 492 
rect 435 492 438 495 
rect 435 495 438 498 
rect 435 498 438 501 
rect 435 501 438 504 
rect 435 504 438 507 
rect 435 507 438 510 
rect 438 0 441 3 
rect 438 3 441 6 
rect 438 6 441 9 
rect 438 9 441 12 
rect 438 12 441 15 
rect 438 15 441 18 
rect 438 18 441 21 
rect 438 21 441 24 
rect 438 24 441 27 
rect 438 27 441 30 
rect 438 30 441 33 
rect 438 33 441 36 
rect 438 36 441 39 
rect 438 39 441 42 
rect 438 42 441 45 
rect 438 45 441 48 
rect 438 48 441 51 
rect 438 51 441 54 
rect 438 54 441 57 
rect 438 57 441 60 
rect 438 60 441 63 
rect 438 63 441 66 
rect 438 66 441 69 
rect 438 69 441 72 
rect 438 72 441 75 
rect 438 75 441 78 
rect 438 78 441 81 
rect 438 81 441 84 
rect 438 84 441 87 
rect 438 87 441 90 
rect 438 90 441 93 
rect 438 93 441 96 
rect 438 96 441 99 
rect 438 99 441 102 
rect 438 102 441 105 
rect 438 105 441 108 
rect 438 108 441 111 
rect 438 111 441 114 
rect 438 114 441 117 
rect 438 117 441 120 
rect 438 120 441 123 
rect 438 123 441 126 
rect 438 126 441 129 
rect 438 129 441 132 
rect 438 132 441 135 
rect 438 135 441 138 
rect 438 138 441 141 
rect 438 141 441 144 
rect 438 144 441 147 
rect 438 147 441 150 
rect 438 150 441 153 
rect 438 153 441 156 
rect 438 156 441 159 
rect 438 159 441 162 
rect 438 162 441 165 
rect 438 165 441 168 
rect 438 168 441 171 
rect 438 171 441 174 
rect 438 174 441 177 
rect 438 177 441 180 
rect 438 180 441 183 
rect 438 183 441 186 
rect 438 186 441 189 
rect 438 189 441 192 
rect 438 192 441 195 
rect 438 195 441 198 
rect 438 198 441 201 
rect 438 201 441 204 
rect 438 204 441 207 
rect 438 207 441 210 
rect 438 210 441 213 
rect 438 213 441 216 
rect 438 216 441 219 
rect 438 219 441 222 
rect 438 222 441 225 
rect 438 225 441 228 
rect 438 228 441 231 
rect 438 231 441 234 
rect 438 234 441 237 
rect 438 237 441 240 
rect 438 240 441 243 
rect 438 243 441 246 
rect 438 246 441 249 
rect 438 249 441 252 
rect 438 252 441 255 
rect 438 255 441 258 
rect 438 258 441 261 
rect 438 261 441 264 
rect 438 264 441 267 
rect 438 267 441 270 
rect 438 270 441 273 
rect 438 273 441 276 
rect 438 276 441 279 
rect 438 279 441 282 
rect 438 282 441 285 
rect 438 285 441 288 
rect 438 288 441 291 
rect 438 291 441 294 
rect 438 294 441 297 
rect 438 297 441 300 
rect 438 300 441 303 
rect 438 303 441 306 
rect 438 306 441 309 
rect 438 309 441 312 
rect 438 312 441 315 
rect 438 315 441 318 
rect 438 318 441 321 
rect 438 321 441 324 
rect 438 324 441 327 
rect 438 327 441 330 
rect 438 330 441 333 
rect 438 333 441 336 
rect 438 336 441 339 
rect 438 339 441 342 
rect 438 342 441 345 
rect 438 345 441 348 
rect 438 348 441 351 
rect 438 351 441 354 
rect 438 354 441 357 
rect 438 357 441 360 
rect 438 360 441 363 
rect 438 363 441 366 
rect 438 366 441 369 
rect 438 369 441 372 
rect 438 372 441 375 
rect 438 375 441 378 
rect 438 378 441 381 
rect 438 381 441 384 
rect 438 384 441 387 
rect 438 387 441 390 
rect 438 390 441 393 
rect 438 393 441 396 
rect 438 396 441 399 
rect 438 399 441 402 
rect 438 402 441 405 
rect 438 405 441 408 
rect 438 408 441 411 
rect 438 411 441 414 
rect 438 414 441 417 
rect 438 417 441 420 
rect 438 420 441 423 
rect 438 423 441 426 
rect 438 426 441 429 
rect 438 429 441 432 
rect 438 432 441 435 
rect 438 435 441 438 
rect 438 438 441 441 
rect 438 441 441 444 
rect 438 444 441 447 
rect 438 447 441 450 
rect 438 450 441 453 
rect 438 453 441 456 
rect 438 456 441 459 
rect 438 459 441 462 
rect 438 462 441 465 
rect 438 465 441 468 
rect 438 468 441 471 
rect 438 471 441 474 
rect 438 474 441 477 
rect 438 477 441 480 
rect 438 480 441 483 
rect 438 483 441 486 
rect 438 486 441 489 
rect 438 489 441 492 
rect 438 492 441 495 
rect 438 495 441 498 
rect 438 498 441 501 
rect 438 501 441 504 
rect 438 504 441 507 
rect 438 507 441 510 
rect 441 0 444 3 
rect 441 3 444 6 
rect 441 6 444 9 
rect 441 9 444 12 
rect 441 12 444 15 
rect 441 15 444 18 
rect 441 18 444 21 
rect 441 21 444 24 
rect 441 24 444 27 
rect 441 27 444 30 
rect 441 30 444 33 
rect 441 33 444 36 
rect 441 36 444 39 
rect 441 39 444 42 
rect 441 42 444 45 
rect 441 45 444 48 
rect 441 48 444 51 
rect 441 51 444 54 
rect 441 54 444 57 
rect 441 57 444 60 
rect 441 60 444 63 
rect 441 63 444 66 
rect 441 66 444 69 
rect 441 69 444 72 
rect 441 72 444 75 
rect 441 75 444 78 
rect 441 78 444 81 
rect 441 81 444 84 
rect 441 84 444 87 
rect 441 87 444 90 
rect 441 90 444 93 
rect 441 93 444 96 
rect 441 96 444 99 
rect 441 99 444 102 
rect 441 102 444 105 
rect 441 105 444 108 
rect 441 108 444 111 
rect 441 111 444 114 
rect 441 114 444 117 
rect 441 117 444 120 
rect 441 120 444 123 
rect 441 123 444 126 
rect 441 126 444 129 
rect 441 129 444 132 
rect 441 132 444 135 
rect 441 135 444 138 
rect 441 138 444 141 
rect 441 141 444 144 
rect 441 144 444 147 
rect 441 147 444 150 
rect 441 150 444 153 
rect 441 153 444 156 
rect 441 156 444 159 
rect 441 159 444 162 
rect 441 162 444 165 
rect 441 165 444 168 
rect 441 168 444 171 
rect 441 171 444 174 
rect 441 174 444 177 
rect 441 177 444 180 
rect 441 180 444 183 
rect 441 183 444 186 
rect 441 186 444 189 
rect 441 189 444 192 
rect 441 192 444 195 
rect 441 195 444 198 
rect 441 198 444 201 
rect 441 201 444 204 
rect 441 204 444 207 
rect 441 207 444 210 
rect 441 210 444 213 
rect 441 213 444 216 
rect 441 216 444 219 
rect 441 219 444 222 
rect 441 222 444 225 
rect 441 225 444 228 
rect 441 228 444 231 
rect 441 231 444 234 
rect 441 234 444 237 
rect 441 237 444 240 
rect 441 240 444 243 
rect 441 243 444 246 
rect 441 246 444 249 
rect 441 249 444 252 
rect 441 252 444 255 
rect 441 255 444 258 
rect 441 258 444 261 
rect 441 261 444 264 
rect 441 264 444 267 
rect 441 267 444 270 
rect 441 270 444 273 
rect 441 273 444 276 
rect 441 276 444 279 
rect 441 279 444 282 
rect 441 282 444 285 
rect 441 285 444 288 
rect 441 288 444 291 
rect 441 291 444 294 
rect 441 294 444 297 
rect 441 297 444 300 
rect 441 300 444 303 
rect 441 303 444 306 
rect 441 306 444 309 
rect 441 309 444 312 
rect 441 312 444 315 
rect 441 315 444 318 
rect 441 318 444 321 
rect 441 321 444 324 
rect 441 324 444 327 
rect 441 327 444 330 
rect 441 330 444 333 
rect 441 333 444 336 
rect 441 336 444 339 
rect 441 339 444 342 
rect 441 342 444 345 
rect 441 345 444 348 
rect 441 348 444 351 
rect 441 351 444 354 
rect 441 354 444 357 
rect 441 357 444 360 
rect 441 360 444 363 
rect 441 363 444 366 
rect 441 366 444 369 
rect 441 369 444 372 
rect 441 372 444 375 
rect 441 375 444 378 
rect 441 378 444 381 
rect 441 381 444 384 
rect 441 384 444 387 
rect 441 387 444 390 
rect 441 390 444 393 
rect 441 393 444 396 
rect 441 396 444 399 
rect 441 399 444 402 
rect 441 402 444 405 
rect 441 405 444 408 
rect 441 408 444 411 
rect 441 411 444 414 
rect 441 414 444 417 
rect 441 417 444 420 
rect 441 420 444 423 
rect 441 423 444 426 
rect 441 426 444 429 
rect 441 429 444 432 
rect 441 432 444 435 
rect 441 435 444 438 
rect 441 438 444 441 
rect 441 441 444 444 
rect 441 444 444 447 
rect 441 447 444 450 
rect 441 450 444 453 
rect 441 453 444 456 
rect 441 456 444 459 
rect 441 459 444 462 
rect 441 462 444 465 
rect 441 465 444 468 
rect 441 468 444 471 
rect 441 471 444 474 
rect 441 474 444 477 
rect 441 477 444 480 
rect 441 480 444 483 
rect 441 483 444 486 
rect 441 486 444 489 
rect 441 489 444 492 
rect 441 492 444 495 
rect 441 495 444 498 
rect 441 498 444 501 
rect 441 501 444 504 
rect 441 504 444 507 
rect 441 507 444 510 
rect 444 0 447 3 
rect 444 3 447 6 
rect 444 6 447 9 
rect 444 9 447 12 
rect 444 12 447 15 
rect 444 15 447 18 
rect 444 18 447 21 
rect 444 21 447 24 
rect 444 24 447 27 
rect 444 27 447 30 
rect 444 30 447 33 
rect 444 33 447 36 
rect 444 36 447 39 
rect 444 39 447 42 
rect 444 42 447 45 
rect 444 45 447 48 
rect 444 48 447 51 
rect 444 51 447 54 
rect 444 54 447 57 
rect 444 57 447 60 
rect 444 60 447 63 
rect 444 63 447 66 
rect 444 66 447 69 
rect 444 69 447 72 
rect 444 72 447 75 
rect 444 75 447 78 
rect 444 78 447 81 
rect 444 81 447 84 
rect 444 84 447 87 
rect 444 87 447 90 
rect 444 90 447 93 
rect 444 93 447 96 
rect 444 96 447 99 
rect 444 99 447 102 
rect 444 102 447 105 
rect 444 105 447 108 
rect 444 108 447 111 
rect 444 111 447 114 
rect 444 114 447 117 
rect 444 117 447 120 
rect 444 120 447 123 
rect 444 123 447 126 
rect 444 126 447 129 
rect 444 129 447 132 
rect 444 132 447 135 
rect 444 135 447 138 
rect 444 138 447 141 
rect 444 141 447 144 
rect 444 144 447 147 
rect 444 147 447 150 
rect 444 150 447 153 
rect 444 153 447 156 
rect 444 156 447 159 
rect 444 159 447 162 
rect 444 162 447 165 
rect 444 165 447 168 
rect 444 168 447 171 
rect 444 171 447 174 
rect 444 174 447 177 
rect 444 177 447 180 
rect 444 180 447 183 
rect 444 183 447 186 
rect 444 186 447 189 
rect 444 189 447 192 
rect 444 192 447 195 
rect 444 195 447 198 
rect 444 198 447 201 
rect 444 201 447 204 
rect 444 204 447 207 
rect 444 207 447 210 
rect 444 210 447 213 
rect 444 213 447 216 
rect 444 216 447 219 
rect 444 219 447 222 
rect 444 222 447 225 
rect 444 225 447 228 
rect 444 228 447 231 
rect 444 231 447 234 
rect 444 234 447 237 
rect 444 237 447 240 
rect 444 240 447 243 
rect 444 243 447 246 
rect 444 246 447 249 
rect 444 249 447 252 
rect 444 252 447 255 
rect 444 255 447 258 
rect 444 258 447 261 
rect 444 261 447 264 
rect 444 264 447 267 
rect 444 267 447 270 
rect 444 270 447 273 
rect 444 273 447 276 
rect 444 276 447 279 
rect 444 279 447 282 
rect 444 282 447 285 
rect 444 285 447 288 
rect 444 288 447 291 
rect 444 291 447 294 
rect 444 294 447 297 
rect 444 297 447 300 
rect 444 300 447 303 
rect 444 303 447 306 
rect 444 306 447 309 
rect 444 309 447 312 
rect 444 312 447 315 
rect 444 315 447 318 
rect 444 318 447 321 
rect 444 321 447 324 
rect 444 324 447 327 
rect 444 327 447 330 
rect 444 330 447 333 
rect 444 333 447 336 
rect 444 336 447 339 
rect 444 339 447 342 
rect 444 342 447 345 
rect 444 345 447 348 
rect 444 348 447 351 
rect 444 351 447 354 
rect 444 354 447 357 
rect 444 357 447 360 
rect 444 360 447 363 
rect 444 363 447 366 
rect 444 366 447 369 
rect 444 369 447 372 
rect 444 372 447 375 
rect 444 375 447 378 
rect 444 378 447 381 
rect 444 381 447 384 
rect 444 384 447 387 
rect 444 387 447 390 
rect 444 390 447 393 
rect 444 393 447 396 
rect 444 396 447 399 
rect 444 399 447 402 
rect 444 402 447 405 
rect 444 405 447 408 
rect 444 408 447 411 
rect 444 411 447 414 
rect 444 414 447 417 
rect 444 417 447 420 
rect 444 420 447 423 
rect 444 423 447 426 
rect 444 426 447 429 
rect 444 429 447 432 
rect 444 432 447 435 
rect 444 435 447 438 
rect 444 438 447 441 
rect 444 441 447 444 
rect 444 444 447 447 
rect 444 447 447 450 
rect 444 450 447 453 
rect 444 453 447 456 
rect 444 456 447 459 
rect 444 459 447 462 
rect 444 462 447 465 
rect 444 465 447 468 
rect 444 468 447 471 
rect 444 471 447 474 
rect 444 474 447 477 
rect 444 477 447 480 
rect 444 480 447 483 
rect 444 483 447 486 
rect 444 486 447 489 
rect 444 489 447 492 
rect 444 492 447 495 
rect 444 495 447 498 
rect 444 498 447 501 
rect 444 501 447 504 
rect 444 504 447 507 
rect 444 507 447 510 
rect 447 0 450 3 
rect 447 3 450 6 
rect 447 6 450 9 
rect 447 9 450 12 
rect 447 12 450 15 
rect 447 15 450 18 
rect 447 18 450 21 
rect 447 21 450 24 
rect 447 24 450 27 
rect 447 27 450 30 
rect 447 30 450 33 
rect 447 33 450 36 
rect 447 36 450 39 
rect 447 39 450 42 
rect 447 42 450 45 
rect 447 45 450 48 
rect 447 48 450 51 
rect 447 51 450 54 
rect 447 54 450 57 
rect 447 57 450 60 
rect 447 60 450 63 
rect 447 63 450 66 
rect 447 66 450 69 
rect 447 69 450 72 
rect 447 72 450 75 
rect 447 75 450 78 
rect 447 78 450 81 
rect 447 81 450 84 
rect 447 84 450 87 
rect 447 87 450 90 
rect 447 90 450 93 
rect 447 93 450 96 
rect 447 96 450 99 
rect 447 99 450 102 
rect 447 102 450 105 
rect 447 105 450 108 
rect 447 108 450 111 
rect 447 111 450 114 
rect 447 114 450 117 
rect 447 117 450 120 
rect 447 120 450 123 
rect 447 123 450 126 
rect 447 126 450 129 
rect 447 129 450 132 
rect 447 132 450 135 
rect 447 135 450 138 
rect 447 138 450 141 
rect 447 141 450 144 
rect 447 144 450 147 
rect 447 147 450 150 
rect 447 150 450 153 
rect 447 153 450 156 
rect 447 156 450 159 
rect 447 159 450 162 
rect 447 162 450 165 
rect 447 165 450 168 
rect 447 168 450 171 
rect 447 171 450 174 
rect 447 174 450 177 
rect 447 177 450 180 
rect 447 180 450 183 
rect 447 183 450 186 
rect 447 186 450 189 
rect 447 189 450 192 
rect 447 192 450 195 
rect 447 195 450 198 
rect 447 198 450 201 
rect 447 201 450 204 
rect 447 204 450 207 
rect 447 207 450 210 
rect 447 210 450 213 
rect 447 213 450 216 
rect 447 216 450 219 
rect 447 219 450 222 
rect 447 222 450 225 
rect 447 225 450 228 
rect 447 228 450 231 
rect 447 231 450 234 
rect 447 234 450 237 
rect 447 237 450 240 
rect 447 240 450 243 
rect 447 243 450 246 
rect 447 246 450 249 
rect 447 249 450 252 
rect 447 252 450 255 
rect 447 255 450 258 
rect 447 258 450 261 
rect 447 261 450 264 
rect 447 264 450 267 
rect 447 267 450 270 
rect 447 270 450 273 
rect 447 273 450 276 
rect 447 276 450 279 
rect 447 279 450 282 
rect 447 282 450 285 
rect 447 285 450 288 
rect 447 288 450 291 
rect 447 291 450 294 
rect 447 294 450 297 
rect 447 297 450 300 
rect 447 300 450 303 
rect 447 303 450 306 
rect 447 306 450 309 
rect 447 309 450 312 
rect 447 312 450 315 
rect 447 315 450 318 
rect 447 318 450 321 
rect 447 321 450 324 
rect 447 324 450 327 
rect 447 327 450 330 
rect 447 330 450 333 
rect 447 333 450 336 
rect 447 336 450 339 
rect 447 339 450 342 
rect 447 342 450 345 
rect 447 345 450 348 
rect 447 348 450 351 
rect 447 351 450 354 
rect 447 354 450 357 
rect 447 357 450 360 
rect 447 360 450 363 
rect 447 363 450 366 
rect 447 366 450 369 
rect 447 369 450 372 
rect 447 372 450 375 
rect 447 375 450 378 
rect 447 378 450 381 
rect 447 381 450 384 
rect 447 384 450 387 
rect 447 387 450 390 
rect 447 390 450 393 
rect 447 393 450 396 
rect 447 396 450 399 
rect 447 399 450 402 
rect 447 402 450 405 
rect 447 405 450 408 
rect 447 408 450 411 
rect 447 411 450 414 
rect 447 414 450 417 
rect 447 417 450 420 
rect 447 420 450 423 
rect 447 423 450 426 
rect 447 426 450 429 
rect 447 429 450 432 
rect 447 432 450 435 
rect 447 435 450 438 
rect 447 438 450 441 
rect 447 441 450 444 
rect 447 444 450 447 
rect 447 447 450 450 
rect 447 450 450 453 
rect 447 453 450 456 
rect 447 456 450 459 
rect 447 459 450 462 
rect 447 462 450 465 
rect 447 465 450 468 
rect 447 468 450 471 
rect 447 471 450 474 
rect 447 474 450 477 
rect 447 477 450 480 
rect 447 480 450 483 
rect 447 483 450 486 
rect 447 486 450 489 
rect 447 489 450 492 
rect 447 492 450 495 
rect 447 495 450 498 
rect 447 498 450 501 
rect 447 501 450 504 
rect 447 504 450 507 
rect 447 507 450 510 
rect 450 0 453 3 
rect 450 3 453 6 
rect 450 6 453 9 
rect 450 9 453 12 
rect 450 12 453 15 
rect 450 15 453 18 
rect 450 18 453 21 
rect 450 21 453 24 
rect 450 24 453 27 
rect 450 27 453 30 
rect 450 30 453 33 
rect 450 33 453 36 
rect 450 36 453 39 
rect 450 39 453 42 
rect 450 42 453 45 
rect 450 45 453 48 
rect 450 48 453 51 
rect 450 51 453 54 
rect 450 54 453 57 
rect 450 57 453 60 
rect 450 60 453 63 
rect 450 63 453 66 
rect 450 66 453 69 
rect 450 69 453 72 
rect 450 72 453 75 
rect 450 75 453 78 
rect 450 78 453 81 
rect 450 81 453 84 
rect 450 84 453 87 
rect 450 87 453 90 
rect 450 90 453 93 
rect 450 93 453 96 
rect 450 96 453 99 
rect 450 99 453 102 
rect 450 102 453 105 
rect 450 105 453 108 
rect 450 108 453 111 
rect 450 111 453 114 
rect 450 114 453 117 
rect 450 117 453 120 
rect 450 120 453 123 
rect 450 123 453 126 
rect 450 126 453 129 
rect 450 129 453 132 
rect 450 132 453 135 
rect 450 135 453 138 
rect 450 138 453 141 
rect 450 141 453 144 
rect 450 144 453 147 
rect 450 147 453 150 
rect 450 150 453 153 
rect 450 153 453 156 
rect 450 156 453 159 
rect 450 159 453 162 
rect 450 162 453 165 
rect 450 165 453 168 
rect 450 168 453 171 
rect 450 171 453 174 
rect 450 174 453 177 
rect 450 177 453 180 
rect 450 180 453 183 
rect 450 183 453 186 
rect 450 186 453 189 
rect 450 189 453 192 
rect 450 192 453 195 
rect 450 195 453 198 
rect 450 198 453 201 
rect 450 201 453 204 
rect 450 204 453 207 
rect 450 207 453 210 
rect 450 210 453 213 
rect 450 213 453 216 
rect 450 216 453 219 
rect 450 219 453 222 
rect 450 222 453 225 
rect 450 225 453 228 
rect 450 228 453 231 
rect 450 231 453 234 
rect 450 234 453 237 
rect 450 237 453 240 
rect 450 240 453 243 
rect 450 243 453 246 
rect 450 246 453 249 
rect 450 249 453 252 
rect 450 252 453 255 
rect 450 255 453 258 
rect 450 258 453 261 
rect 450 261 453 264 
rect 450 264 453 267 
rect 450 267 453 270 
rect 450 270 453 273 
rect 450 273 453 276 
rect 450 276 453 279 
rect 450 279 453 282 
rect 450 282 453 285 
rect 450 285 453 288 
rect 450 288 453 291 
rect 450 291 453 294 
rect 450 294 453 297 
rect 450 297 453 300 
rect 450 300 453 303 
rect 450 303 453 306 
rect 450 306 453 309 
rect 450 309 453 312 
rect 450 312 453 315 
rect 450 315 453 318 
rect 450 318 453 321 
rect 450 321 453 324 
rect 450 324 453 327 
rect 450 327 453 330 
rect 450 330 453 333 
rect 450 333 453 336 
rect 450 336 453 339 
rect 450 339 453 342 
rect 450 342 453 345 
rect 450 345 453 348 
rect 450 348 453 351 
rect 450 351 453 354 
rect 450 354 453 357 
rect 450 357 453 360 
rect 450 360 453 363 
rect 450 363 453 366 
rect 450 366 453 369 
rect 450 369 453 372 
rect 450 372 453 375 
rect 450 375 453 378 
rect 450 378 453 381 
rect 450 381 453 384 
rect 450 384 453 387 
rect 450 387 453 390 
rect 450 390 453 393 
rect 450 393 453 396 
rect 450 396 453 399 
rect 450 399 453 402 
rect 450 402 453 405 
rect 450 405 453 408 
rect 450 408 453 411 
rect 450 411 453 414 
rect 450 414 453 417 
rect 450 417 453 420 
rect 450 420 453 423 
rect 450 423 453 426 
rect 450 426 453 429 
rect 450 429 453 432 
rect 450 432 453 435 
rect 450 435 453 438 
rect 450 438 453 441 
rect 450 441 453 444 
rect 450 444 453 447 
rect 450 447 453 450 
rect 450 450 453 453 
rect 450 453 453 456 
rect 450 456 453 459 
rect 450 459 453 462 
rect 450 462 453 465 
rect 450 465 453 468 
rect 450 468 453 471 
rect 450 471 453 474 
rect 450 474 453 477 
rect 450 477 453 480 
rect 450 480 453 483 
rect 450 483 453 486 
rect 450 486 453 489 
rect 450 489 453 492 
rect 450 492 453 495 
rect 450 495 453 498 
rect 450 498 453 501 
rect 450 501 453 504 
rect 450 504 453 507 
rect 450 507 453 510 
rect 453 0 456 3 
rect 453 3 456 6 
rect 453 6 456 9 
rect 453 9 456 12 
rect 453 12 456 15 
rect 453 15 456 18 
rect 453 18 456 21 
rect 453 21 456 24 
rect 453 24 456 27 
rect 453 27 456 30 
rect 453 30 456 33 
rect 453 33 456 36 
rect 453 36 456 39 
rect 453 39 456 42 
rect 453 42 456 45 
rect 453 45 456 48 
rect 453 48 456 51 
rect 453 51 456 54 
rect 453 54 456 57 
rect 453 57 456 60 
rect 453 60 456 63 
rect 453 63 456 66 
rect 453 66 456 69 
rect 453 69 456 72 
rect 453 72 456 75 
rect 453 75 456 78 
rect 453 78 456 81 
rect 453 81 456 84 
rect 453 84 456 87 
rect 453 87 456 90 
rect 453 90 456 93 
rect 453 93 456 96 
rect 453 96 456 99 
rect 453 99 456 102 
rect 453 102 456 105 
rect 453 105 456 108 
rect 453 108 456 111 
rect 453 111 456 114 
rect 453 114 456 117 
rect 453 117 456 120 
rect 453 120 456 123 
rect 453 123 456 126 
rect 453 126 456 129 
rect 453 129 456 132 
rect 453 132 456 135 
rect 453 135 456 138 
rect 453 138 456 141 
rect 453 141 456 144 
rect 453 144 456 147 
rect 453 147 456 150 
rect 453 150 456 153 
rect 453 153 456 156 
rect 453 156 456 159 
rect 453 159 456 162 
rect 453 162 456 165 
rect 453 165 456 168 
rect 453 168 456 171 
rect 453 171 456 174 
rect 453 174 456 177 
rect 453 177 456 180 
rect 453 180 456 183 
rect 453 183 456 186 
rect 453 186 456 189 
rect 453 189 456 192 
rect 453 192 456 195 
rect 453 195 456 198 
rect 453 198 456 201 
rect 453 201 456 204 
rect 453 204 456 207 
rect 453 207 456 210 
rect 453 210 456 213 
rect 453 213 456 216 
rect 453 216 456 219 
rect 453 219 456 222 
rect 453 222 456 225 
rect 453 225 456 228 
rect 453 228 456 231 
rect 453 231 456 234 
rect 453 234 456 237 
rect 453 237 456 240 
rect 453 240 456 243 
rect 453 243 456 246 
rect 453 246 456 249 
rect 453 249 456 252 
rect 453 252 456 255 
rect 453 255 456 258 
rect 453 258 456 261 
rect 453 261 456 264 
rect 453 264 456 267 
rect 453 267 456 270 
rect 453 270 456 273 
rect 453 273 456 276 
rect 453 276 456 279 
rect 453 279 456 282 
rect 453 282 456 285 
rect 453 285 456 288 
rect 453 288 456 291 
rect 453 291 456 294 
rect 453 294 456 297 
rect 453 297 456 300 
rect 453 300 456 303 
rect 453 303 456 306 
rect 453 306 456 309 
rect 453 309 456 312 
rect 453 312 456 315 
rect 453 315 456 318 
rect 453 318 456 321 
rect 453 321 456 324 
rect 453 324 456 327 
rect 453 327 456 330 
rect 453 330 456 333 
rect 453 333 456 336 
rect 453 336 456 339 
rect 453 339 456 342 
rect 453 342 456 345 
rect 453 345 456 348 
rect 453 348 456 351 
rect 453 351 456 354 
rect 453 354 456 357 
rect 453 357 456 360 
rect 453 360 456 363 
rect 453 363 456 366 
rect 453 366 456 369 
rect 453 369 456 372 
rect 453 372 456 375 
rect 453 375 456 378 
rect 453 378 456 381 
rect 453 381 456 384 
rect 453 384 456 387 
rect 453 387 456 390 
rect 453 390 456 393 
rect 453 393 456 396 
rect 453 396 456 399 
rect 453 399 456 402 
rect 453 402 456 405 
rect 453 405 456 408 
rect 453 408 456 411 
rect 453 411 456 414 
rect 453 414 456 417 
rect 453 417 456 420 
rect 453 420 456 423 
rect 453 423 456 426 
rect 453 426 456 429 
rect 453 429 456 432 
rect 453 432 456 435 
rect 453 435 456 438 
rect 453 438 456 441 
rect 453 441 456 444 
rect 453 444 456 447 
rect 453 447 456 450 
rect 453 450 456 453 
rect 453 453 456 456 
rect 453 456 456 459 
rect 453 459 456 462 
rect 453 462 456 465 
rect 453 465 456 468 
rect 453 468 456 471 
rect 453 471 456 474 
rect 453 474 456 477 
rect 453 477 456 480 
rect 453 480 456 483 
rect 453 483 456 486 
rect 453 486 456 489 
rect 453 489 456 492 
rect 453 492 456 495 
rect 453 495 456 498 
rect 453 498 456 501 
rect 453 501 456 504 
rect 453 504 456 507 
rect 453 507 456 510 
rect 456 0 459 3 
rect 456 3 459 6 
rect 456 6 459 9 
rect 456 9 459 12 
rect 456 12 459 15 
rect 456 15 459 18 
rect 456 18 459 21 
rect 456 21 459 24 
rect 456 24 459 27 
rect 456 27 459 30 
rect 456 30 459 33 
rect 456 33 459 36 
rect 456 36 459 39 
rect 456 39 459 42 
rect 456 42 459 45 
rect 456 45 459 48 
rect 456 48 459 51 
rect 456 51 459 54 
rect 456 54 459 57 
rect 456 57 459 60 
rect 456 60 459 63 
rect 456 63 459 66 
rect 456 66 459 69 
rect 456 69 459 72 
rect 456 72 459 75 
rect 456 75 459 78 
rect 456 78 459 81 
rect 456 81 459 84 
rect 456 84 459 87 
rect 456 87 459 90 
rect 456 90 459 93 
rect 456 93 459 96 
rect 456 96 459 99 
rect 456 99 459 102 
rect 456 102 459 105 
rect 456 105 459 108 
rect 456 108 459 111 
rect 456 111 459 114 
rect 456 114 459 117 
rect 456 117 459 120 
rect 456 120 459 123 
rect 456 123 459 126 
rect 456 126 459 129 
rect 456 129 459 132 
rect 456 132 459 135 
rect 456 135 459 138 
rect 456 138 459 141 
rect 456 141 459 144 
rect 456 144 459 147 
rect 456 147 459 150 
rect 456 150 459 153 
rect 456 153 459 156 
rect 456 156 459 159 
rect 456 159 459 162 
rect 456 162 459 165 
rect 456 165 459 168 
rect 456 168 459 171 
rect 456 171 459 174 
rect 456 174 459 177 
rect 456 177 459 180 
rect 456 180 459 183 
rect 456 183 459 186 
rect 456 186 459 189 
rect 456 189 459 192 
rect 456 192 459 195 
rect 456 195 459 198 
rect 456 198 459 201 
rect 456 201 459 204 
rect 456 204 459 207 
rect 456 207 459 210 
rect 456 210 459 213 
rect 456 213 459 216 
rect 456 216 459 219 
rect 456 219 459 222 
rect 456 222 459 225 
rect 456 225 459 228 
rect 456 228 459 231 
rect 456 231 459 234 
rect 456 234 459 237 
rect 456 237 459 240 
rect 456 240 459 243 
rect 456 243 459 246 
rect 456 246 459 249 
rect 456 249 459 252 
rect 456 252 459 255 
rect 456 255 459 258 
rect 456 258 459 261 
rect 456 261 459 264 
rect 456 264 459 267 
rect 456 267 459 270 
rect 456 270 459 273 
rect 456 273 459 276 
rect 456 276 459 279 
rect 456 279 459 282 
rect 456 282 459 285 
rect 456 285 459 288 
rect 456 288 459 291 
rect 456 291 459 294 
rect 456 294 459 297 
rect 456 297 459 300 
rect 456 300 459 303 
rect 456 303 459 306 
rect 456 306 459 309 
rect 456 309 459 312 
rect 456 312 459 315 
rect 456 315 459 318 
rect 456 318 459 321 
rect 456 321 459 324 
rect 456 324 459 327 
rect 456 327 459 330 
rect 456 330 459 333 
rect 456 333 459 336 
rect 456 336 459 339 
rect 456 339 459 342 
rect 456 342 459 345 
rect 456 345 459 348 
rect 456 348 459 351 
rect 456 351 459 354 
rect 456 354 459 357 
rect 456 357 459 360 
rect 456 360 459 363 
rect 456 363 459 366 
rect 456 366 459 369 
rect 456 369 459 372 
rect 456 372 459 375 
rect 456 375 459 378 
rect 456 378 459 381 
rect 456 381 459 384 
rect 456 384 459 387 
rect 456 387 459 390 
rect 456 390 459 393 
rect 456 393 459 396 
rect 456 396 459 399 
rect 456 399 459 402 
rect 456 402 459 405 
rect 456 405 459 408 
rect 456 408 459 411 
rect 456 411 459 414 
rect 456 414 459 417 
rect 456 417 459 420 
rect 456 420 459 423 
rect 456 423 459 426 
rect 456 426 459 429 
rect 456 429 459 432 
rect 456 432 459 435 
rect 456 435 459 438 
rect 456 438 459 441 
rect 456 441 459 444 
rect 456 444 459 447 
rect 456 447 459 450 
rect 456 450 459 453 
rect 456 453 459 456 
rect 456 456 459 459 
rect 456 459 459 462 
rect 456 462 459 465 
rect 456 465 459 468 
rect 456 468 459 471 
rect 456 471 459 474 
rect 456 474 459 477 
rect 456 477 459 480 
rect 456 480 459 483 
rect 456 483 459 486 
rect 456 486 459 489 
rect 456 489 459 492 
rect 456 492 459 495 
rect 456 495 459 498 
rect 456 498 459 501 
rect 456 501 459 504 
rect 456 504 459 507 
rect 456 507 459 510 
rect 459 0 462 3 
rect 459 3 462 6 
rect 459 6 462 9 
rect 459 9 462 12 
rect 459 12 462 15 
rect 459 15 462 18 
rect 459 18 462 21 
rect 459 21 462 24 
rect 459 24 462 27 
rect 459 27 462 30 
rect 459 30 462 33 
rect 459 33 462 36 
rect 459 36 462 39 
rect 459 39 462 42 
rect 459 42 462 45 
rect 459 45 462 48 
rect 459 48 462 51 
rect 459 51 462 54 
rect 459 54 462 57 
rect 459 57 462 60 
rect 459 60 462 63 
rect 459 63 462 66 
rect 459 66 462 69 
rect 459 69 462 72 
rect 459 72 462 75 
rect 459 75 462 78 
rect 459 78 462 81 
rect 459 81 462 84 
rect 459 84 462 87 
rect 459 87 462 90 
rect 459 90 462 93 
rect 459 93 462 96 
rect 459 96 462 99 
rect 459 99 462 102 
rect 459 102 462 105 
rect 459 105 462 108 
rect 459 108 462 111 
rect 459 111 462 114 
rect 459 114 462 117 
rect 459 117 462 120 
rect 459 120 462 123 
rect 459 123 462 126 
rect 459 126 462 129 
rect 459 129 462 132 
rect 459 132 462 135 
rect 459 135 462 138 
rect 459 138 462 141 
rect 459 141 462 144 
rect 459 144 462 147 
rect 459 147 462 150 
rect 459 150 462 153 
rect 459 153 462 156 
rect 459 156 462 159 
rect 459 159 462 162 
rect 459 162 462 165 
rect 459 165 462 168 
rect 459 168 462 171 
rect 459 171 462 174 
rect 459 174 462 177 
rect 459 177 462 180 
rect 459 180 462 183 
rect 459 183 462 186 
rect 459 186 462 189 
rect 459 189 462 192 
rect 459 192 462 195 
rect 459 195 462 198 
rect 459 198 462 201 
rect 459 201 462 204 
rect 459 204 462 207 
rect 459 207 462 210 
rect 459 210 462 213 
rect 459 213 462 216 
rect 459 216 462 219 
rect 459 219 462 222 
rect 459 222 462 225 
rect 459 225 462 228 
rect 459 228 462 231 
rect 459 231 462 234 
rect 459 234 462 237 
rect 459 237 462 240 
rect 459 240 462 243 
rect 459 243 462 246 
rect 459 246 462 249 
rect 459 249 462 252 
rect 459 252 462 255 
rect 459 255 462 258 
rect 459 258 462 261 
rect 459 261 462 264 
rect 459 264 462 267 
rect 459 267 462 270 
rect 459 270 462 273 
rect 459 273 462 276 
rect 459 276 462 279 
rect 459 279 462 282 
rect 459 282 462 285 
rect 459 285 462 288 
rect 459 288 462 291 
rect 459 291 462 294 
rect 459 294 462 297 
rect 459 297 462 300 
rect 459 300 462 303 
rect 459 303 462 306 
rect 459 306 462 309 
rect 459 309 462 312 
rect 459 312 462 315 
rect 459 315 462 318 
rect 459 318 462 321 
rect 459 321 462 324 
rect 459 324 462 327 
rect 459 327 462 330 
rect 459 330 462 333 
rect 459 333 462 336 
rect 459 336 462 339 
rect 459 339 462 342 
rect 459 342 462 345 
rect 459 345 462 348 
rect 459 348 462 351 
rect 459 351 462 354 
rect 459 354 462 357 
rect 459 357 462 360 
rect 459 360 462 363 
rect 459 363 462 366 
rect 459 366 462 369 
rect 459 369 462 372 
rect 459 372 462 375 
rect 459 375 462 378 
rect 459 378 462 381 
rect 459 381 462 384 
rect 459 384 462 387 
rect 459 387 462 390 
rect 459 390 462 393 
rect 459 393 462 396 
rect 459 396 462 399 
rect 459 399 462 402 
rect 459 402 462 405 
rect 459 405 462 408 
rect 459 408 462 411 
rect 459 411 462 414 
rect 459 414 462 417 
rect 459 417 462 420 
rect 459 420 462 423 
rect 459 423 462 426 
rect 459 426 462 429 
rect 459 429 462 432 
rect 459 432 462 435 
rect 459 435 462 438 
rect 459 438 462 441 
rect 459 441 462 444 
rect 459 444 462 447 
rect 459 447 462 450 
rect 459 450 462 453 
rect 459 453 462 456 
rect 459 456 462 459 
rect 459 459 462 462 
rect 459 462 462 465 
rect 459 465 462 468 
rect 459 468 462 471 
rect 459 471 462 474 
rect 459 474 462 477 
rect 459 477 462 480 
rect 459 480 462 483 
rect 459 483 462 486 
rect 459 486 462 489 
rect 459 489 462 492 
rect 459 492 462 495 
rect 459 495 462 498 
rect 459 498 462 501 
rect 459 501 462 504 
rect 459 504 462 507 
rect 459 507 462 510 
rect 462 0 465 3 
rect 462 3 465 6 
rect 462 6 465 9 
rect 462 9 465 12 
rect 462 12 465 15 
rect 462 15 465 18 
rect 462 18 465 21 
rect 462 21 465 24 
rect 462 24 465 27 
rect 462 27 465 30 
rect 462 30 465 33 
rect 462 33 465 36 
rect 462 36 465 39 
rect 462 39 465 42 
rect 462 42 465 45 
rect 462 45 465 48 
rect 462 48 465 51 
rect 462 51 465 54 
rect 462 54 465 57 
rect 462 57 465 60 
rect 462 60 465 63 
rect 462 63 465 66 
rect 462 66 465 69 
rect 462 69 465 72 
rect 462 72 465 75 
rect 462 75 465 78 
rect 462 78 465 81 
rect 462 81 465 84 
rect 462 84 465 87 
rect 462 87 465 90 
rect 462 90 465 93 
rect 462 93 465 96 
rect 462 96 465 99 
rect 462 99 465 102 
rect 462 102 465 105 
rect 462 105 465 108 
rect 462 108 465 111 
rect 462 111 465 114 
rect 462 114 465 117 
rect 462 117 465 120 
rect 462 120 465 123 
rect 462 123 465 126 
rect 462 126 465 129 
rect 462 129 465 132 
rect 462 132 465 135 
rect 462 135 465 138 
rect 462 138 465 141 
rect 462 141 465 144 
rect 462 144 465 147 
rect 462 147 465 150 
rect 462 150 465 153 
rect 462 153 465 156 
rect 462 156 465 159 
rect 462 159 465 162 
rect 462 162 465 165 
rect 462 165 465 168 
rect 462 168 465 171 
rect 462 171 465 174 
rect 462 174 465 177 
rect 462 177 465 180 
rect 462 180 465 183 
rect 462 183 465 186 
rect 462 186 465 189 
rect 462 189 465 192 
rect 462 192 465 195 
rect 462 195 465 198 
rect 462 198 465 201 
rect 462 201 465 204 
rect 462 204 465 207 
rect 462 207 465 210 
rect 462 210 465 213 
rect 462 213 465 216 
rect 462 216 465 219 
rect 462 219 465 222 
rect 462 222 465 225 
rect 462 225 465 228 
rect 462 228 465 231 
rect 462 231 465 234 
rect 462 234 465 237 
rect 462 237 465 240 
rect 462 240 465 243 
rect 462 243 465 246 
rect 462 246 465 249 
rect 462 249 465 252 
rect 462 252 465 255 
rect 462 255 465 258 
rect 462 258 465 261 
rect 462 261 465 264 
rect 462 264 465 267 
rect 462 267 465 270 
rect 462 270 465 273 
rect 462 273 465 276 
rect 462 276 465 279 
rect 462 279 465 282 
rect 462 282 465 285 
rect 462 285 465 288 
rect 462 288 465 291 
rect 462 291 465 294 
rect 462 294 465 297 
rect 462 297 465 300 
rect 462 300 465 303 
rect 462 303 465 306 
rect 462 306 465 309 
rect 462 309 465 312 
rect 462 312 465 315 
rect 462 315 465 318 
rect 462 318 465 321 
rect 462 321 465 324 
rect 462 324 465 327 
rect 462 327 465 330 
rect 462 330 465 333 
rect 462 333 465 336 
rect 462 336 465 339 
rect 462 339 465 342 
rect 462 342 465 345 
rect 462 345 465 348 
rect 462 348 465 351 
rect 462 351 465 354 
rect 462 354 465 357 
rect 462 357 465 360 
rect 462 360 465 363 
rect 462 363 465 366 
rect 462 366 465 369 
rect 462 369 465 372 
rect 462 372 465 375 
rect 462 375 465 378 
rect 462 378 465 381 
rect 462 381 465 384 
rect 462 384 465 387 
rect 462 387 465 390 
rect 462 390 465 393 
rect 462 393 465 396 
rect 462 396 465 399 
rect 462 399 465 402 
rect 462 402 465 405 
rect 462 405 465 408 
rect 462 408 465 411 
rect 462 411 465 414 
rect 462 414 465 417 
rect 462 417 465 420 
rect 462 420 465 423 
rect 462 423 465 426 
rect 462 426 465 429 
rect 462 429 465 432 
rect 462 432 465 435 
rect 462 435 465 438 
rect 462 438 465 441 
rect 462 441 465 444 
rect 462 444 465 447 
rect 462 447 465 450 
rect 462 450 465 453 
rect 462 453 465 456 
rect 462 456 465 459 
rect 462 459 465 462 
rect 462 462 465 465 
rect 462 465 465 468 
rect 462 468 465 471 
rect 462 471 465 474 
rect 462 474 465 477 
rect 462 477 465 480 
rect 462 480 465 483 
rect 462 483 465 486 
rect 462 486 465 489 
rect 462 489 465 492 
rect 462 492 465 495 
rect 462 495 465 498 
rect 462 498 465 501 
rect 462 501 465 504 
rect 462 504 465 507 
rect 462 507 465 510 
rect 465 0 468 3 
rect 465 3 468 6 
rect 465 6 468 9 
rect 465 9 468 12 
rect 465 12 468 15 
rect 465 15 468 18 
rect 465 18 468 21 
rect 465 21 468 24 
rect 465 24 468 27 
rect 465 27 468 30 
rect 465 30 468 33 
rect 465 33 468 36 
rect 465 36 468 39 
rect 465 39 468 42 
rect 465 42 468 45 
rect 465 45 468 48 
rect 465 48 468 51 
rect 465 51 468 54 
rect 465 54 468 57 
rect 465 57 468 60 
rect 465 60 468 63 
rect 465 63 468 66 
rect 465 66 468 69 
rect 465 69 468 72 
rect 465 72 468 75 
rect 465 75 468 78 
rect 465 78 468 81 
rect 465 81 468 84 
rect 465 84 468 87 
rect 465 87 468 90 
rect 465 90 468 93 
rect 465 93 468 96 
rect 465 96 468 99 
rect 465 99 468 102 
rect 465 102 468 105 
rect 465 105 468 108 
rect 465 108 468 111 
rect 465 111 468 114 
rect 465 114 468 117 
rect 465 117 468 120 
rect 465 120 468 123 
rect 465 123 468 126 
rect 465 126 468 129 
rect 465 129 468 132 
rect 465 132 468 135 
rect 465 135 468 138 
rect 465 138 468 141 
rect 465 141 468 144 
rect 465 144 468 147 
rect 465 147 468 150 
rect 465 150 468 153 
rect 465 153 468 156 
rect 465 156 468 159 
rect 465 159 468 162 
rect 465 162 468 165 
rect 465 165 468 168 
rect 465 168 468 171 
rect 465 171 468 174 
rect 465 174 468 177 
rect 465 177 468 180 
rect 465 180 468 183 
rect 465 183 468 186 
rect 465 186 468 189 
rect 465 189 468 192 
rect 465 192 468 195 
rect 465 195 468 198 
rect 465 198 468 201 
rect 465 201 468 204 
rect 465 204 468 207 
rect 465 207 468 210 
rect 465 210 468 213 
rect 465 213 468 216 
rect 465 216 468 219 
rect 465 219 468 222 
rect 465 222 468 225 
rect 465 225 468 228 
rect 465 228 468 231 
rect 465 231 468 234 
rect 465 234 468 237 
rect 465 237 468 240 
rect 465 240 468 243 
rect 465 243 468 246 
rect 465 246 468 249 
rect 465 249 468 252 
rect 465 252 468 255 
rect 465 255 468 258 
rect 465 258 468 261 
rect 465 261 468 264 
rect 465 264 468 267 
rect 465 267 468 270 
rect 465 270 468 273 
rect 465 273 468 276 
rect 465 276 468 279 
rect 465 279 468 282 
rect 465 282 468 285 
rect 465 285 468 288 
rect 465 288 468 291 
rect 465 291 468 294 
rect 465 294 468 297 
rect 465 297 468 300 
rect 465 300 468 303 
rect 465 303 468 306 
rect 465 306 468 309 
rect 465 309 468 312 
rect 465 312 468 315 
rect 465 315 468 318 
rect 465 318 468 321 
rect 465 321 468 324 
rect 465 324 468 327 
rect 465 327 468 330 
rect 465 330 468 333 
rect 465 333 468 336 
rect 465 336 468 339 
rect 465 339 468 342 
rect 465 342 468 345 
rect 465 345 468 348 
rect 465 348 468 351 
rect 465 351 468 354 
rect 465 354 468 357 
rect 465 357 468 360 
rect 465 360 468 363 
rect 465 363 468 366 
rect 465 366 468 369 
rect 465 369 468 372 
rect 465 372 468 375 
rect 465 375 468 378 
rect 465 378 468 381 
rect 465 381 468 384 
rect 465 384 468 387 
rect 465 387 468 390 
rect 465 390 468 393 
rect 465 393 468 396 
rect 465 396 468 399 
rect 465 399 468 402 
rect 465 402 468 405 
rect 465 405 468 408 
rect 465 408 468 411 
rect 465 411 468 414 
rect 465 414 468 417 
rect 465 417 468 420 
rect 465 420 468 423 
rect 465 423 468 426 
rect 465 426 468 429 
rect 465 429 468 432 
rect 465 432 468 435 
rect 465 435 468 438 
rect 465 438 468 441 
rect 465 441 468 444 
rect 465 444 468 447 
rect 465 447 468 450 
rect 465 450 468 453 
rect 465 453 468 456 
rect 465 456 468 459 
rect 465 459 468 462 
rect 465 462 468 465 
rect 465 465 468 468 
rect 465 468 468 471 
rect 465 471 468 474 
rect 465 474 468 477 
rect 465 477 468 480 
rect 465 480 468 483 
rect 465 483 468 486 
rect 465 486 468 489 
rect 465 489 468 492 
rect 465 492 468 495 
rect 465 495 468 498 
rect 465 498 468 501 
rect 465 501 468 504 
rect 465 504 468 507 
rect 465 507 468 510 
rect 468 0 471 3 
rect 468 3 471 6 
rect 468 6 471 9 
rect 468 9 471 12 
rect 468 12 471 15 
rect 468 15 471 18 
rect 468 18 471 21 
rect 468 21 471 24 
rect 468 24 471 27 
rect 468 27 471 30 
rect 468 30 471 33 
rect 468 33 471 36 
rect 468 36 471 39 
rect 468 39 471 42 
rect 468 42 471 45 
rect 468 45 471 48 
rect 468 48 471 51 
rect 468 51 471 54 
rect 468 54 471 57 
rect 468 57 471 60 
rect 468 60 471 63 
rect 468 63 471 66 
rect 468 66 471 69 
rect 468 69 471 72 
rect 468 72 471 75 
rect 468 75 471 78 
rect 468 78 471 81 
rect 468 81 471 84 
rect 468 84 471 87 
rect 468 87 471 90 
rect 468 90 471 93 
rect 468 93 471 96 
rect 468 96 471 99 
rect 468 99 471 102 
rect 468 102 471 105 
rect 468 105 471 108 
rect 468 108 471 111 
rect 468 111 471 114 
rect 468 114 471 117 
rect 468 117 471 120 
rect 468 120 471 123 
rect 468 123 471 126 
rect 468 126 471 129 
rect 468 129 471 132 
rect 468 132 471 135 
rect 468 135 471 138 
rect 468 138 471 141 
rect 468 141 471 144 
rect 468 144 471 147 
rect 468 147 471 150 
rect 468 150 471 153 
rect 468 153 471 156 
rect 468 156 471 159 
rect 468 159 471 162 
rect 468 162 471 165 
rect 468 165 471 168 
rect 468 168 471 171 
rect 468 171 471 174 
rect 468 174 471 177 
rect 468 177 471 180 
rect 468 180 471 183 
rect 468 183 471 186 
rect 468 186 471 189 
rect 468 189 471 192 
rect 468 192 471 195 
rect 468 195 471 198 
rect 468 198 471 201 
rect 468 201 471 204 
rect 468 204 471 207 
rect 468 207 471 210 
rect 468 210 471 213 
rect 468 213 471 216 
rect 468 216 471 219 
rect 468 219 471 222 
rect 468 222 471 225 
rect 468 225 471 228 
rect 468 228 471 231 
rect 468 231 471 234 
rect 468 234 471 237 
rect 468 237 471 240 
rect 468 240 471 243 
rect 468 243 471 246 
rect 468 246 471 249 
rect 468 249 471 252 
rect 468 252 471 255 
rect 468 255 471 258 
rect 468 258 471 261 
rect 468 261 471 264 
rect 468 264 471 267 
rect 468 267 471 270 
rect 468 270 471 273 
rect 468 273 471 276 
rect 468 276 471 279 
rect 468 279 471 282 
rect 468 282 471 285 
rect 468 285 471 288 
rect 468 288 471 291 
rect 468 291 471 294 
rect 468 294 471 297 
rect 468 297 471 300 
rect 468 300 471 303 
rect 468 303 471 306 
rect 468 306 471 309 
rect 468 309 471 312 
rect 468 312 471 315 
rect 468 315 471 318 
rect 468 318 471 321 
rect 468 321 471 324 
rect 468 324 471 327 
rect 468 327 471 330 
rect 468 330 471 333 
rect 468 333 471 336 
rect 468 336 471 339 
rect 468 339 471 342 
rect 468 342 471 345 
rect 468 345 471 348 
rect 468 348 471 351 
rect 468 351 471 354 
rect 468 354 471 357 
rect 468 357 471 360 
rect 468 360 471 363 
rect 468 363 471 366 
rect 468 366 471 369 
rect 468 369 471 372 
rect 468 372 471 375 
rect 468 375 471 378 
rect 468 378 471 381 
rect 468 381 471 384 
rect 468 384 471 387 
rect 468 387 471 390 
rect 468 390 471 393 
rect 468 393 471 396 
rect 468 396 471 399 
rect 468 399 471 402 
rect 468 402 471 405 
rect 468 405 471 408 
rect 468 408 471 411 
rect 468 411 471 414 
rect 468 414 471 417 
rect 468 417 471 420 
rect 468 420 471 423 
rect 468 423 471 426 
rect 468 426 471 429 
rect 468 429 471 432 
rect 468 432 471 435 
rect 468 435 471 438 
rect 468 438 471 441 
rect 468 441 471 444 
rect 468 444 471 447 
rect 468 447 471 450 
rect 468 450 471 453 
rect 468 453 471 456 
rect 468 456 471 459 
rect 468 459 471 462 
rect 468 462 471 465 
rect 468 465 471 468 
rect 468 468 471 471 
rect 468 471 471 474 
rect 468 474 471 477 
rect 468 477 471 480 
rect 468 480 471 483 
rect 468 483 471 486 
rect 468 486 471 489 
rect 468 489 471 492 
rect 468 492 471 495 
rect 468 495 471 498 
rect 468 498 471 501 
rect 468 501 471 504 
rect 468 504 471 507 
rect 468 507 471 510 
rect 471 0 474 3 
rect 471 3 474 6 
rect 471 6 474 9 
rect 471 9 474 12 
rect 471 12 474 15 
rect 471 15 474 18 
rect 471 18 474 21 
rect 471 21 474 24 
rect 471 24 474 27 
rect 471 27 474 30 
rect 471 30 474 33 
rect 471 33 474 36 
rect 471 36 474 39 
rect 471 39 474 42 
rect 471 42 474 45 
rect 471 45 474 48 
rect 471 48 474 51 
rect 471 51 474 54 
rect 471 54 474 57 
rect 471 57 474 60 
rect 471 60 474 63 
rect 471 63 474 66 
rect 471 66 474 69 
rect 471 69 474 72 
rect 471 72 474 75 
rect 471 75 474 78 
rect 471 78 474 81 
rect 471 81 474 84 
rect 471 84 474 87 
rect 471 87 474 90 
rect 471 90 474 93 
rect 471 93 474 96 
rect 471 96 474 99 
rect 471 99 474 102 
rect 471 102 474 105 
rect 471 105 474 108 
rect 471 108 474 111 
rect 471 111 474 114 
rect 471 114 474 117 
rect 471 117 474 120 
rect 471 120 474 123 
rect 471 123 474 126 
rect 471 126 474 129 
rect 471 129 474 132 
rect 471 132 474 135 
rect 471 135 474 138 
rect 471 138 474 141 
rect 471 141 474 144 
rect 471 144 474 147 
rect 471 147 474 150 
rect 471 150 474 153 
rect 471 153 474 156 
rect 471 156 474 159 
rect 471 159 474 162 
rect 471 162 474 165 
rect 471 165 474 168 
rect 471 168 474 171 
rect 471 171 474 174 
rect 471 174 474 177 
rect 471 177 474 180 
rect 471 180 474 183 
rect 471 183 474 186 
rect 471 186 474 189 
rect 471 189 474 192 
rect 471 192 474 195 
rect 471 195 474 198 
rect 471 198 474 201 
rect 471 201 474 204 
rect 471 204 474 207 
rect 471 207 474 210 
rect 471 210 474 213 
rect 471 213 474 216 
rect 471 216 474 219 
rect 471 219 474 222 
rect 471 222 474 225 
rect 471 225 474 228 
rect 471 228 474 231 
rect 471 231 474 234 
rect 471 234 474 237 
rect 471 237 474 240 
rect 471 240 474 243 
rect 471 243 474 246 
rect 471 246 474 249 
rect 471 249 474 252 
rect 471 252 474 255 
rect 471 255 474 258 
rect 471 258 474 261 
rect 471 261 474 264 
rect 471 264 474 267 
rect 471 267 474 270 
rect 471 270 474 273 
rect 471 273 474 276 
rect 471 276 474 279 
rect 471 279 474 282 
rect 471 282 474 285 
rect 471 285 474 288 
rect 471 288 474 291 
rect 471 291 474 294 
rect 471 294 474 297 
rect 471 297 474 300 
rect 471 300 474 303 
rect 471 303 474 306 
rect 471 306 474 309 
rect 471 309 474 312 
rect 471 312 474 315 
rect 471 315 474 318 
rect 471 318 474 321 
rect 471 321 474 324 
rect 471 324 474 327 
rect 471 327 474 330 
rect 471 330 474 333 
rect 471 333 474 336 
rect 471 336 474 339 
rect 471 339 474 342 
rect 471 342 474 345 
rect 471 345 474 348 
rect 471 348 474 351 
rect 471 351 474 354 
rect 471 354 474 357 
rect 471 357 474 360 
rect 471 360 474 363 
rect 471 363 474 366 
rect 471 366 474 369 
rect 471 369 474 372 
rect 471 372 474 375 
rect 471 375 474 378 
rect 471 378 474 381 
rect 471 381 474 384 
rect 471 384 474 387 
rect 471 387 474 390 
rect 471 390 474 393 
rect 471 393 474 396 
rect 471 396 474 399 
rect 471 399 474 402 
rect 471 402 474 405 
rect 471 405 474 408 
rect 471 408 474 411 
rect 471 411 474 414 
rect 471 414 474 417 
rect 471 417 474 420 
rect 471 420 474 423 
rect 471 423 474 426 
rect 471 426 474 429 
rect 471 429 474 432 
rect 471 432 474 435 
rect 471 435 474 438 
rect 471 438 474 441 
rect 471 441 474 444 
rect 471 444 474 447 
rect 471 447 474 450 
rect 471 450 474 453 
rect 471 453 474 456 
rect 471 456 474 459 
rect 471 459 474 462 
rect 471 462 474 465 
rect 471 465 474 468 
rect 471 468 474 471 
rect 471 471 474 474 
rect 471 474 474 477 
rect 471 477 474 480 
rect 471 480 474 483 
rect 471 483 474 486 
rect 471 486 474 489 
rect 471 489 474 492 
rect 471 492 474 495 
rect 471 495 474 498 
rect 471 498 474 501 
rect 471 501 474 504 
rect 471 504 474 507 
rect 471 507 474 510 
rect 474 0 477 3 
rect 474 3 477 6 
rect 474 6 477 9 
rect 474 9 477 12 
rect 474 12 477 15 
rect 474 15 477 18 
rect 474 18 477 21 
rect 474 21 477 24 
rect 474 24 477 27 
rect 474 27 477 30 
rect 474 30 477 33 
rect 474 33 477 36 
rect 474 36 477 39 
rect 474 39 477 42 
rect 474 42 477 45 
rect 474 45 477 48 
rect 474 48 477 51 
rect 474 51 477 54 
rect 474 54 477 57 
rect 474 57 477 60 
rect 474 60 477 63 
rect 474 63 477 66 
rect 474 66 477 69 
rect 474 69 477 72 
rect 474 72 477 75 
rect 474 75 477 78 
rect 474 78 477 81 
rect 474 81 477 84 
rect 474 84 477 87 
rect 474 87 477 90 
rect 474 90 477 93 
rect 474 93 477 96 
rect 474 96 477 99 
rect 474 99 477 102 
rect 474 102 477 105 
rect 474 105 477 108 
rect 474 108 477 111 
rect 474 111 477 114 
rect 474 114 477 117 
rect 474 117 477 120 
rect 474 120 477 123 
rect 474 123 477 126 
rect 474 126 477 129 
rect 474 129 477 132 
rect 474 132 477 135 
rect 474 135 477 138 
rect 474 138 477 141 
rect 474 141 477 144 
rect 474 144 477 147 
rect 474 147 477 150 
rect 474 150 477 153 
rect 474 153 477 156 
rect 474 156 477 159 
rect 474 159 477 162 
rect 474 162 477 165 
rect 474 165 477 168 
rect 474 168 477 171 
rect 474 171 477 174 
rect 474 174 477 177 
rect 474 177 477 180 
rect 474 180 477 183 
rect 474 183 477 186 
rect 474 186 477 189 
rect 474 189 477 192 
rect 474 192 477 195 
rect 474 195 477 198 
rect 474 198 477 201 
rect 474 201 477 204 
rect 474 204 477 207 
rect 474 207 477 210 
rect 474 210 477 213 
rect 474 213 477 216 
rect 474 216 477 219 
rect 474 219 477 222 
rect 474 222 477 225 
rect 474 225 477 228 
rect 474 228 477 231 
rect 474 231 477 234 
rect 474 234 477 237 
rect 474 237 477 240 
rect 474 240 477 243 
rect 474 243 477 246 
rect 474 246 477 249 
rect 474 249 477 252 
rect 474 252 477 255 
rect 474 255 477 258 
rect 474 258 477 261 
rect 474 261 477 264 
rect 474 264 477 267 
rect 474 267 477 270 
rect 474 270 477 273 
rect 474 273 477 276 
rect 474 276 477 279 
rect 474 279 477 282 
rect 474 282 477 285 
rect 474 285 477 288 
rect 474 288 477 291 
rect 474 291 477 294 
rect 474 294 477 297 
rect 474 297 477 300 
rect 474 300 477 303 
rect 474 303 477 306 
rect 474 306 477 309 
rect 474 309 477 312 
rect 474 312 477 315 
rect 474 315 477 318 
rect 474 318 477 321 
rect 474 321 477 324 
rect 474 324 477 327 
rect 474 327 477 330 
rect 474 330 477 333 
rect 474 333 477 336 
rect 474 336 477 339 
rect 474 339 477 342 
rect 474 342 477 345 
rect 474 345 477 348 
rect 474 348 477 351 
rect 474 351 477 354 
rect 474 354 477 357 
rect 474 357 477 360 
rect 474 360 477 363 
rect 474 363 477 366 
rect 474 366 477 369 
rect 474 369 477 372 
rect 474 372 477 375 
rect 474 375 477 378 
rect 474 378 477 381 
rect 474 381 477 384 
rect 474 384 477 387 
rect 474 387 477 390 
rect 474 390 477 393 
rect 474 393 477 396 
rect 474 396 477 399 
rect 474 399 477 402 
rect 474 402 477 405 
rect 474 405 477 408 
rect 474 408 477 411 
rect 474 411 477 414 
rect 474 414 477 417 
rect 474 417 477 420 
rect 474 420 477 423 
rect 474 423 477 426 
rect 474 426 477 429 
rect 474 429 477 432 
rect 474 432 477 435 
rect 474 435 477 438 
rect 474 438 477 441 
rect 474 441 477 444 
rect 474 444 477 447 
rect 474 447 477 450 
rect 474 450 477 453 
rect 474 453 477 456 
rect 474 456 477 459 
rect 474 459 477 462 
rect 474 462 477 465 
rect 474 465 477 468 
rect 474 468 477 471 
rect 474 471 477 474 
rect 474 474 477 477 
rect 474 477 477 480 
rect 474 480 477 483 
rect 474 483 477 486 
rect 474 486 477 489 
rect 474 489 477 492 
rect 474 492 477 495 
rect 474 495 477 498 
rect 474 498 477 501 
rect 474 501 477 504 
rect 474 504 477 507 
rect 474 507 477 510 
rect 477 0 480 3 
rect 477 3 480 6 
rect 477 6 480 9 
rect 477 9 480 12 
rect 477 12 480 15 
rect 477 15 480 18 
rect 477 18 480 21 
rect 477 21 480 24 
rect 477 24 480 27 
rect 477 27 480 30 
rect 477 30 480 33 
rect 477 33 480 36 
rect 477 36 480 39 
rect 477 39 480 42 
rect 477 42 480 45 
rect 477 45 480 48 
rect 477 48 480 51 
rect 477 51 480 54 
rect 477 54 480 57 
rect 477 57 480 60 
rect 477 60 480 63 
rect 477 63 480 66 
rect 477 66 480 69 
rect 477 69 480 72 
rect 477 72 480 75 
rect 477 75 480 78 
rect 477 78 480 81 
rect 477 81 480 84 
rect 477 84 480 87 
rect 477 87 480 90 
rect 477 90 480 93 
rect 477 93 480 96 
rect 477 96 480 99 
rect 477 99 480 102 
rect 477 102 480 105 
rect 477 105 480 108 
rect 477 108 480 111 
rect 477 111 480 114 
rect 477 114 480 117 
rect 477 117 480 120 
rect 477 120 480 123 
rect 477 123 480 126 
rect 477 126 480 129 
rect 477 129 480 132 
rect 477 132 480 135 
rect 477 135 480 138 
rect 477 138 480 141 
rect 477 141 480 144 
rect 477 144 480 147 
rect 477 147 480 150 
rect 477 150 480 153 
rect 477 153 480 156 
rect 477 156 480 159 
rect 477 159 480 162 
rect 477 162 480 165 
rect 477 165 480 168 
rect 477 168 480 171 
rect 477 171 480 174 
rect 477 174 480 177 
rect 477 177 480 180 
rect 477 180 480 183 
rect 477 183 480 186 
rect 477 186 480 189 
rect 477 189 480 192 
rect 477 192 480 195 
rect 477 195 480 198 
rect 477 198 480 201 
rect 477 201 480 204 
rect 477 204 480 207 
rect 477 207 480 210 
rect 477 210 480 213 
rect 477 213 480 216 
rect 477 216 480 219 
rect 477 219 480 222 
rect 477 222 480 225 
rect 477 225 480 228 
rect 477 228 480 231 
rect 477 231 480 234 
rect 477 234 480 237 
rect 477 237 480 240 
rect 477 240 480 243 
rect 477 243 480 246 
rect 477 246 480 249 
rect 477 249 480 252 
rect 477 252 480 255 
rect 477 255 480 258 
rect 477 258 480 261 
rect 477 261 480 264 
rect 477 264 480 267 
rect 477 267 480 270 
rect 477 270 480 273 
rect 477 273 480 276 
rect 477 276 480 279 
rect 477 279 480 282 
rect 477 282 480 285 
rect 477 285 480 288 
rect 477 288 480 291 
rect 477 291 480 294 
rect 477 294 480 297 
rect 477 297 480 300 
rect 477 300 480 303 
rect 477 303 480 306 
rect 477 306 480 309 
rect 477 309 480 312 
rect 477 312 480 315 
rect 477 315 480 318 
rect 477 318 480 321 
rect 477 321 480 324 
rect 477 324 480 327 
rect 477 327 480 330 
rect 477 330 480 333 
rect 477 333 480 336 
rect 477 336 480 339 
rect 477 339 480 342 
rect 477 342 480 345 
rect 477 345 480 348 
rect 477 348 480 351 
rect 477 351 480 354 
rect 477 354 480 357 
rect 477 357 480 360 
rect 477 360 480 363 
rect 477 363 480 366 
rect 477 366 480 369 
rect 477 369 480 372 
rect 477 372 480 375 
rect 477 375 480 378 
rect 477 378 480 381 
rect 477 381 480 384 
rect 477 384 480 387 
rect 477 387 480 390 
rect 477 390 480 393 
rect 477 393 480 396 
rect 477 396 480 399 
rect 477 399 480 402 
rect 477 402 480 405 
rect 477 405 480 408 
rect 477 408 480 411 
rect 477 411 480 414 
rect 477 414 480 417 
rect 477 417 480 420 
rect 477 420 480 423 
rect 477 423 480 426 
rect 477 426 480 429 
rect 477 429 480 432 
rect 477 432 480 435 
rect 477 435 480 438 
rect 477 438 480 441 
rect 477 441 480 444 
rect 477 444 480 447 
rect 477 447 480 450 
rect 477 450 480 453 
rect 477 453 480 456 
rect 477 456 480 459 
rect 477 459 480 462 
rect 477 462 480 465 
rect 477 465 480 468 
rect 477 468 480 471 
rect 477 471 480 474 
rect 477 474 480 477 
rect 477 477 480 480 
rect 477 480 480 483 
rect 477 483 480 486 
rect 477 486 480 489 
rect 477 489 480 492 
rect 477 492 480 495 
rect 477 495 480 498 
rect 477 498 480 501 
rect 477 501 480 504 
rect 477 504 480 507 
rect 477 507 480 510 
rect 480 0 483 3 
rect 480 3 483 6 
rect 480 6 483 9 
rect 480 9 483 12 
rect 480 12 483 15 
rect 480 15 483 18 
rect 480 18 483 21 
rect 480 21 483 24 
rect 480 24 483 27 
rect 480 27 483 30 
rect 480 30 483 33 
rect 480 33 483 36 
rect 480 36 483 39 
rect 480 39 483 42 
rect 480 42 483 45 
rect 480 45 483 48 
rect 480 48 483 51 
rect 480 51 483 54 
rect 480 54 483 57 
rect 480 57 483 60 
rect 480 60 483 63 
rect 480 63 483 66 
rect 480 66 483 69 
rect 480 69 483 72 
rect 480 72 483 75 
rect 480 75 483 78 
rect 480 78 483 81 
rect 480 81 483 84 
rect 480 84 483 87 
rect 480 87 483 90 
rect 480 90 483 93 
rect 480 93 483 96 
rect 480 96 483 99 
rect 480 99 483 102 
rect 480 102 483 105 
rect 480 105 483 108 
rect 480 108 483 111 
rect 480 111 483 114 
rect 480 114 483 117 
rect 480 117 483 120 
rect 480 120 483 123 
rect 480 123 483 126 
rect 480 126 483 129 
rect 480 129 483 132 
rect 480 132 483 135 
rect 480 135 483 138 
rect 480 138 483 141 
rect 480 141 483 144 
rect 480 144 483 147 
rect 480 147 483 150 
rect 480 150 483 153 
rect 480 153 483 156 
rect 480 156 483 159 
rect 480 159 483 162 
rect 480 162 483 165 
rect 480 165 483 168 
rect 480 168 483 171 
rect 480 171 483 174 
rect 480 174 483 177 
rect 480 177 483 180 
rect 480 180 483 183 
rect 480 183 483 186 
rect 480 186 483 189 
rect 480 189 483 192 
rect 480 192 483 195 
rect 480 195 483 198 
rect 480 198 483 201 
rect 480 201 483 204 
rect 480 204 483 207 
rect 480 207 483 210 
rect 480 210 483 213 
rect 480 213 483 216 
rect 480 216 483 219 
rect 480 219 483 222 
rect 480 222 483 225 
rect 480 225 483 228 
rect 480 228 483 231 
rect 480 231 483 234 
rect 480 234 483 237 
rect 480 237 483 240 
rect 480 240 483 243 
rect 480 243 483 246 
rect 480 246 483 249 
rect 480 249 483 252 
rect 480 252 483 255 
rect 480 255 483 258 
rect 480 258 483 261 
rect 480 261 483 264 
rect 480 264 483 267 
rect 480 267 483 270 
rect 480 270 483 273 
rect 480 273 483 276 
rect 480 276 483 279 
rect 480 279 483 282 
rect 480 282 483 285 
rect 480 285 483 288 
rect 480 288 483 291 
rect 480 291 483 294 
rect 480 294 483 297 
rect 480 297 483 300 
rect 480 300 483 303 
rect 480 303 483 306 
rect 480 306 483 309 
rect 480 309 483 312 
rect 480 312 483 315 
rect 480 315 483 318 
rect 480 318 483 321 
rect 480 321 483 324 
rect 480 324 483 327 
rect 480 327 483 330 
rect 480 330 483 333 
rect 480 333 483 336 
rect 480 336 483 339 
rect 480 339 483 342 
rect 480 342 483 345 
rect 480 345 483 348 
rect 480 348 483 351 
rect 480 351 483 354 
rect 480 354 483 357 
rect 480 357 483 360 
rect 480 360 483 363 
rect 480 363 483 366 
rect 480 366 483 369 
rect 480 369 483 372 
rect 480 372 483 375 
rect 480 375 483 378 
rect 480 378 483 381 
rect 480 381 483 384 
rect 480 384 483 387 
rect 480 387 483 390 
rect 480 390 483 393 
rect 480 393 483 396 
rect 480 396 483 399 
rect 480 399 483 402 
rect 480 402 483 405 
rect 480 405 483 408 
rect 480 408 483 411 
rect 480 411 483 414 
rect 480 414 483 417 
rect 480 417 483 420 
rect 480 420 483 423 
rect 480 423 483 426 
rect 480 426 483 429 
rect 480 429 483 432 
rect 480 432 483 435 
rect 480 435 483 438 
rect 480 438 483 441 
rect 480 441 483 444 
rect 480 444 483 447 
rect 480 447 483 450 
rect 480 450 483 453 
rect 480 453 483 456 
rect 480 456 483 459 
rect 480 459 483 462 
rect 480 462 483 465 
rect 480 465 483 468 
rect 480 468 483 471 
rect 480 471 483 474 
rect 480 474 483 477 
rect 480 477 483 480 
rect 480 480 483 483 
rect 480 483 483 486 
rect 480 486 483 489 
rect 480 489 483 492 
rect 480 492 483 495 
rect 480 495 483 498 
rect 480 498 483 501 
rect 480 501 483 504 
rect 480 504 483 507 
rect 480 507 483 510 
rect 483 0 486 3 
rect 483 3 486 6 
rect 483 6 486 9 
rect 483 9 486 12 
rect 483 12 486 15 
rect 483 15 486 18 
rect 483 18 486 21 
rect 483 21 486 24 
rect 483 24 486 27 
rect 483 27 486 30 
rect 483 30 486 33 
rect 483 33 486 36 
rect 483 36 486 39 
rect 483 39 486 42 
rect 483 42 486 45 
rect 483 45 486 48 
rect 483 48 486 51 
rect 483 51 486 54 
rect 483 54 486 57 
rect 483 57 486 60 
rect 483 60 486 63 
rect 483 63 486 66 
rect 483 66 486 69 
rect 483 69 486 72 
rect 483 72 486 75 
rect 483 75 486 78 
rect 483 78 486 81 
rect 483 81 486 84 
rect 483 84 486 87 
rect 483 87 486 90 
rect 483 90 486 93 
rect 483 93 486 96 
rect 483 96 486 99 
rect 483 99 486 102 
rect 483 102 486 105 
rect 483 105 486 108 
rect 483 108 486 111 
rect 483 111 486 114 
rect 483 114 486 117 
rect 483 117 486 120 
rect 483 120 486 123 
rect 483 123 486 126 
rect 483 126 486 129 
rect 483 129 486 132 
rect 483 132 486 135 
rect 483 135 486 138 
rect 483 138 486 141 
rect 483 141 486 144 
rect 483 144 486 147 
rect 483 147 486 150 
rect 483 150 486 153 
rect 483 153 486 156 
rect 483 156 486 159 
rect 483 159 486 162 
rect 483 162 486 165 
rect 483 165 486 168 
rect 483 168 486 171 
rect 483 171 486 174 
rect 483 174 486 177 
rect 483 177 486 180 
rect 483 180 486 183 
rect 483 183 486 186 
rect 483 186 486 189 
rect 483 189 486 192 
rect 483 192 486 195 
rect 483 195 486 198 
rect 483 198 486 201 
rect 483 201 486 204 
rect 483 204 486 207 
rect 483 207 486 210 
rect 483 210 486 213 
rect 483 213 486 216 
rect 483 216 486 219 
rect 483 219 486 222 
rect 483 222 486 225 
rect 483 225 486 228 
rect 483 228 486 231 
rect 483 231 486 234 
rect 483 234 486 237 
rect 483 237 486 240 
rect 483 240 486 243 
rect 483 243 486 246 
rect 483 246 486 249 
rect 483 249 486 252 
rect 483 252 486 255 
rect 483 255 486 258 
rect 483 258 486 261 
rect 483 261 486 264 
rect 483 264 486 267 
rect 483 267 486 270 
rect 483 270 486 273 
rect 483 273 486 276 
rect 483 276 486 279 
rect 483 279 486 282 
rect 483 282 486 285 
rect 483 285 486 288 
rect 483 288 486 291 
rect 483 291 486 294 
rect 483 294 486 297 
rect 483 297 486 300 
rect 483 300 486 303 
rect 483 303 486 306 
rect 483 306 486 309 
rect 483 309 486 312 
rect 483 312 486 315 
rect 483 315 486 318 
rect 483 318 486 321 
rect 483 321 486 324 
rect 483 324 486 327 
rect 483 327 486 330 
rect 483 330 486 333 
rect 483 333 486 336 
rect 483 336 486 339 
rect 483 339 486 342 
rect 483 342 486 345 
rect 483 345 486 348 
rect 483 348 486 351 
rect 483 351 486 354 
rect 483 354 486 357 
rect 483 357 486 360 
rect 483 360 486 363 
rect 483 363 486 366 
rect 483 366 486 369 
rect 483 369 486 372 
rect 483 372 486 375 
rect 483 375 486 378 
rect 483 378 486 381 
rect 483 381 486 384 
rect 483 384 486 387 
rect 483 387 486 390 
rect 483 390 486 393 
rect 483 393 486 396 
rect 483 396 486 399 
rect 483 399 486 402 
rect 483 402 486 405 
rect 483 405 486 408 
rect 483 408 486 411 
rect 483 411 486 414 
rect 483 414 486 417 
rect 483 417 486 420 
rect 483 420 486 423 
rect 483 423 486 426 
rect 483 426 486 429 
rect 483 429 486 432 
rect 483 432 486 435 
rect 483 435 486 438 
rect 483 438 486 441 
rect 483 441 486 444 
rect 483 444 486 447 
rect 483 447 486 450 
rect 483 450 486 453 
rect 483 453 486 456 
rect 483 456 486 459 
rect 483 459 486 462 
rect 483 462 486 465 
rect 483 465 486 468 
rect 483 468 486 471 
rect 483 471 486 474 
rect 483 474 486 477 
rect 483 477 486 480 
rect 483 480 486 483 
rect 483 483 486 486 
rect 483 486 486 489 
rect 483 489 486 492 
rect 483 492 486 495 
rect 483 495 486 498 
rect 483 498 486 501 
rect 483 501 486 504 
rect 483 504 486 507 
rect 483 507 486 510 
rect 486 0 489 3 
rect 486 3 489 6 
rect 486 6 489 9 
rect 486 9 489 12 
rect 486 12 489 15 
rect 486 15 489 18 
rect 486 18 489 21 
rect 486 21 489 24 
rect 486 24 489 27 
rect 486 27 489 30 
rect 486 30 489 33 
rect 486 33 489 36 
rect 486 36 489 39 
rect 486 39 489 42 
rect 486 42 489 45 
rect 486 45 489 48 
rect 486 48 489 51 
rect 486 51 489 54 
rect 486 54 489 57 
rect 486 57 489 60 
rect 486 60 489 63 
rect 486 63 489 66 
rect 486 66 489 69 
rect 486 69 489 72 
rect 486 72 489 75 
rect 486 75 489 78 
rect 486 78 489 81 
rect 486 81 489 84 
rect 486 84 489 87 
rect 486 87 489 90 
rect 486 90 489 93 
rect 486 93 489 96 
rect 486 96 489 99 
rect 486 99 489 102 
rect 486 102 489 105 
rect 486 105 489 108 
rect 486 108 489 111 
rect 486 111 489 114 
rect 486 114 489 117 
rect 486 117 489 120 
rect 486 120 489 123 
rect 486 123 489 126 
rect 486 126 489 129 
rect 486 129 489 132 
rect 486 132 489 135 
rect 486 135 489 138 
rect 486 138 489 141 
rect 486 141 489 144 
rect 486 144 489 147 
rect 486 147 489 150 
rect 486 150 489 153 
rect 486 153 489 156 
rect 486 156 489 159 
rect 486 159 489 162 
rect 486 162 489 165 
rect 486 165 489 168 
rect 486 168 489 171 
rect 486 171 489 174 
rect 486 174 489 177 
rect 486 177 489 180 
rect 486 180 489 183 
rect 486 183 489 186 
rect 486 186 489 189 
rect 486 189 489 192 
rect 486 192 489 195 
rect 486 195 489 198 
rect 486 198 489 201 
rect 486 201 489 204 
rect 486 204 489 207 
rect 486 207 489 210 
rect 486 210 489 213 
rect 486 213 489 216 
rect 486 216 489 219 
rect 486 219 489 222 
rect 486 222 489 225 
rect 486 225 489 228 
rect 486 228 489 231 
rect 486 231 489 234 
rect 486 234 489 237 
rect 486 237 489 240 
rect 486 240 489 243 
rect 486 243 489 246 
rect 486 246 489 249 
rect 486 249 489 252 
rect 486 252 489 255 
rect 486 255 489 258 
rect 486 258 489 261 
rect 486 261 489 264 
rect 486 264 489 267 
rect 486 267 489 270 
rect 486 270 489 273 
rect 486 273 489 276 
rect 486 276 489 279 
rect 486 279 489 282 
rect 486 282 489 285 
rect 486 285 489 288 
rect 486 288 489 291 
rect 486 291 489 294 
rect 486 294 489 297 
rect 486 297 489 300 
rect 486 300 489 303 
rect 486 303 489 306 
rect 486 306 489 309 
rect 486 309 489 312 
rect 486 312 489 315 
rect 486 315 489 318 
rect 486 318 489 321 
rect 486 321 489 324 
rect 486 324 489 327 
rect 486 327 489 330 
rect 486 330 489 333 
rect 486 333 489 336 
rect 486 336 489 339 
rect 486 339 489 342 
rect 486 342 489 345 
rect 486 345 489 348 
rect 486 348 489 351 
rect 486 351 489 354 
rect 486 354 489 357 
rect 486 357 489 360 
rect 486 360 489 363 
rect 486 363 489 366 
rect 486 366 489 369 
rect 486 369 489 372 
rect 486 372 489 375 
rect 486 375 489 378 
rect 486 378 489 381 
rect 486 381 489 384 
rect 486 384 489 387 
rect 486 387 489 390 
rect 486 390 489 393 
rect 486 393 489 396 
rect 486 396 489 399 
rect 486 399 489 402 
rect 486 402 489 405 
rect 486 405 489 408 
rect 486 408 489 411 
rect 486 411 489 414 
rect 486 414 489 417 
rect 486 417 489 420 
rect 486 420 489 423 
rect 486 423 489 426 
rect 486 426 489 429 
rect 486 429 489 432 
rect 486 432 489 435 
rect 486 435 489 438 
rect 486 438 489 441 
rect 486 441 489 444 
rect 486 444 489 447 
rect 486 447 489 450 
rect 486 450 489 453 
rect 486 453 489 456 
rect 486 456 489 459 
rect 486 459 489 462 
rect 486 462 489 465 
rect 486 465 489 468 
rect 486 468 489 471 
rect 486 471 489 474 
rect 486 474 489 477 
rect 486 477 489 480 
rect 486 480 489 483 
rect 486 483 489 486 
rect 486 486 489 489 
rect 486 489 489 492 
rect 486 492 489 495 
rect 486 495 489 498 
rect 486 498 489 501 
rect 486 501 489 504 
rect 486 504 489 507 
rect 486 507 489 510 
rect 489 0 492 3 
rect 489 3 492 6 
rect 489 6 492 9 
rect 489 9 492 12 
rect 489 12 492 15 
rect 489 15 492 18 
rect 489 18 492 21 
rect 489 21 492 24 
rect 489 24 492 27 
rect 489 27 492 30 
rect 489 30 492 33 
rect 489 33 492 36 
rect 489 36 492 39 
rect 489 39 492 42 
rect 489 42 492 45 
rect 489 45 492 48 
rect 489 48 492 51 
rect 489 51 492 54 
rect 489 54 492 57 
rect 489 57 492 60 
rect 489 60 492 63 
rect 489 63 492 66 
rect 489 66 492 69 
rect 489 69 492 72 
rect 489 72 492 75 
rect 489 75 492 78 
rect 489 78 492 81 
rect 489 81 492 84 
rect 489 84 492 87 
rect 489 87 492 90 
rect 489 90 492 93 
rect 489 93 492 96 
rect 489 96 492 99 
rect 489 99 492 102 
rect 489 102 492 105 
rect 489 105 492 108 
rect 489 108 492 111 
rect 489 111 492 114 
rect 489 114 492 117 
rect 489 117 492 120 
rect 489 120 492 123 
rect 489 123 492 126 
rect 489 126 492 129 
rect 489 129 492 132 
rect 489 132 492 135 
rect 489 135 492 138 
rect 489 138 492 141 
rect 489 141 492 144 
rect 489 144 492 147 
rect 489 147 492 150 
rect 489 150 492 153 
rect 489 153 492 156 
rect 489 156 492 159 
rect 489 159 492 162 
rect 489 162 492 165 
rect 489 165 492 168 
rect 489 168 492 171 
rect 489 171 492 174 
rect 489 174 492 177 
rect 489 177 492 180 
rect 489 180 492 183 
rect 489 183 492 186 
rect 489 186 492 189 
rect 489 189 492 192 
rect 489 192 492 195 
rect 489 195 492 198 
rect 489 198 492 201 
rect 489 201 492 204 
rect 489 204 492 207 
rect 489 207 492 210 
rect 489 210 492 213 
rect 489 213 492 216 
rect 489 216 492 219 
rect 489 219 492 222 
rect 489 222 492 225 
rect 489 225 492 228 
rect 489 228 492 231 
rect 489 231 492 234 
rect 489 234 492 237 
rect 489 237 492 240 
rect 489 240 492 243 
rect 489 243 492 246 
rect 489 246 492 249 
rect 489 249 492 252 
rect 489 252 492 255 
rect 489 255 492 258 
rect 489 258 492 261 
rect 489 261 492 264 
rect 489 264 492 267 
rect 489 267 492 270 
rect 489 270 492 273 
rect 489 273 492 276 
rect 489 276 492 279 
rect 489 279 492 282 
rect 489 282 492 285 
rect 489 285 492 288 
rect 489 288 492 291 
rect 489 291 492 294 
rect 489 294 492 297 
rect 489 297 492 300 
rect 489 300 492 303 
rect 489 303 492 306 
rect 489 306 492 309 
rect 489 309 492 312 
rect 489 312 492 315 
rect 489 315 492 318 
rect 489 318 492 321 
rect 489 321 492 324 
rect 489 324 492 327 
rect 489 327 492 330 
rect 489 330 492 333 
rect 489 333 492 336 
rect 489 336 492 339 
rect 489 339 492 342 
rect 489 342 492 345 
rect 489 345 492 348 
rect 489 348 492 351 
rect 489 351 492 354 
rect 489 354 492 357 
rect 489 357 492 360 
rect 489 360 492 363 
rect 489 363 492 366 
rect 489 366 492 369 
rect 489 369 492 372 
rect 489 372 492 375 
rect 489 375 492 378 
rect 489 378 492 381 
rect 489 381 492 384 
rect 489 384 492 387 
rect 489 387 492 390 
rect 489 390 492 393 
rect 489 393 492 396 
rect 489 396 492 399 
rect 489 399 492 402 
rect 489 402 492 405 
rect 489 405 492 408 
rect 489 408 492 411 
rect 489 411 492 414 
rect 489 414 492 417 
rect 489 417 492 420 
rect 489 420 492 423 
rect 489 423 492 426 
rect 489 426 492 429 
rect 489 429 492 432 
rect 489 432 492 435 
rect 489 435 492 438 
rect 489 438 492 441 
rect 489 441 492 444 
rect 489 444 492 447 
rect 489 447 492 450 
rect 489 450 492 453 
rect 489 453 492 456 
rect 489 456 492 459 
rect 489 459 492 462 
rect 489 462 492 465 
rect 489 465 492 468 
rect 489 468 492 471 
rect 489 471 492 474 
rect 489 474 492 477 
rect 489 477 492 480 
rect 489 480 492 483 
rect 489 483 492 486 
rect 489 486 492 489 
rect 489 489 492 492 
rect 489 492 492 495 
rect 489 495 492 498 
rect 489 498 492 501 
rect 489 501 492 504 
rect 489 504 492 507 
rect 489 507 492 510 
rect 492 0 495 3 
rect 492 3 495 6 
rect 492 6 495 9 
rect 492 9 495 12 
rect 492 12 495 15 
rect 492 15 495 18 
rect 492 18 495 21 
rect 492 21 495 24 
rect 492 24 495 27 
rect 492 27 495 30 
rect 492 30 495 33 
rect 492 33 495 36 
rect 492 36 495 39 
rect 492 39 495 42 
rect 492 42 495 45 
rect 492 45 495 48 
rect 492 48 495 51 
rect 492 51 495 54 
rect 492 54 495 57 
rect 492 57 495 60 
rect 492 60 495 63 
rect 492 63 495 66 
rect 492 66 495 69 
rect 492 69 495 72 
rect 492 72 495 75 
rect 492 75 495 78 
rect 492 78 495 81 
rect 492 81 495 84 
rect 492 84 495 87 
rect 492 87 495 90 
rect 492 90 495 93 
rect 492 93 495 96 
rect 492 96 495 99 
rect 492 99 495 102 
rect 492 102 495 105 
rect 492 105 495 108 
rect 492 108 495 111 
rect 492 111 495 114 
rect 492 114 495 117 
rect 492 117 495 120 
rect 492 120 495 123 
rect 492 123 495 126 
rect 492 126 495 129 
rect 492 129 495 132 
rect 492 132 495 135 
rect 492 135 495 138 
rect 492 138 495 141 
rect 492 141 495 144 
rect 492 144 495 147 
rect 492 147 495 150 
rect 492 150 495 153 
rect 492 153 495 156 
rect 492 156 495 159 
rect 492 159 495 162 
rect 492 162 495 165 
rect 492 165 495 168 
rect 492 168 495 171 
rect 492 171 495 174 
rect 492 174 495 177 
rect 492 177 495 180 
rect 492 180 495 183 
rect 492 183 495 186 
rect 492 186 495 189 
rect 492 189 495 192 
rect 492 192 495 195 
rect 492 195 495 198 
rect 492 198 495 201 
rect 492 201 495 204 
rect 492 204 495 207 
rect 492 207 495 210 
rect 492 210 495 213 
rect 492 213 495 216 
rect 492 216 495 219 
rect 492 219 495 222 
rect 492 222 495 225 
rect 492 225 495 228 
rect 492 228 495 231 
rect 492 231 495 234 
rect 492 234 495 237 
rect 492 237 495 240 
rect 492 240 495 243 
rect 492 243 495 246 
rect 492 246 495 249 
rect 492 249 495 252 
rect 492 252 495 255 
rect 492 255 495 258 
rect 492 258 495 261 
rect 492 261 495 264 
rect 492 264 495 267 
rect 492 267 495 270 
rect 492 270 495 273 
rect 492 273 495 276 
rect 492 276 495 279 
rect 492 279 495 282 
rect 492 282 495 285 
rect 492 285 495 288 
rect 492 288 495 291 
rect 492 291 495 294 
rect 492 294 495 297 
rect 492 297 495 300 
rect 492 300 495 303 
rect 492 303 495 306 
rect 492 306 495 309 
rect 492 309 495 312 
rect 492 312 495 315 
rect 492 315 495 318 
rect 492 318 495 321 
rect 492 321 495 324 
rect 492 324 495 327 
rect 492 327 495 330 
rect 492 330 495 333 
rect 492 333 495 336 
rect 492 336 495 339 
rect 492 339 495 342 
rect 492 342 495 345 
rect 492 345 495 348 
rect 492 348 495 351 
rect 492 351 495 354 
rect 492 354 495 357 
rect 492 357 495 360 
rect 492 360 495 363 
rect 492 363 495 366 
rect 492 366 495 369 
rect 492 369 495 372 
rect 492 372 495 375 
rect 492 375 495 378 
rect 492 378 495 381 
rect 492 381 495 384 
rect 492 384 495 387 
rect 492 387 495 390 
rect 492 390 495 393 
rect 492 393 495 396 
rect 492 396 495 399 
rect 492 399 495 402 
rect 492 402 495 405 
rect 492 405 495 408 
rect 492 408 495 411 
rect 492 411 495 414 
rect 492 414 495 417 
rect 492 417 495 420 
rect 492 420 495 423 
rect 492 423 495 426 
rect 492 426 495 429 
rect 492 429 495 432 
rect 492 432 495 435 
rect 492 435 495 438 
rect 492 438 495 441 
rect 492 441 495 444 
rect 492 444 495 447 
rect 492 447 495 450 
rect 492 450 495 453 
rect 492 453 495 456 
rect 492 456 495 459 
rect 492 459 495 462 
rect 492 462 495 465 
rect 492 465 495 468 
rect 492 468 495 471 
rect 492 471 495 474 
rect 492 474 495 477 
rect 492 477 495 480 
rect 492 480 495 483 
rect 492 483 495 486 
rect 492 486 495 489 
rect 492 489 495 492 
rect 492 492 495 495 
rect 492 495 495 498 
rect 492 498 495 501 
rect 492 501 495 504 
rect 492 504 495 507 
rect 492 507 495 510 
rect 495 0 498 3 
rect 495 3 498 6 
rect 495 6 498 9 
rect 495 9 498 12 
rect 495 12 498 15 
rect 495 15 498 18 
rect 495 18 498 21 
rect 495 21 498 24 
rect 495 24 498 27 
rect 495 27 498 30 
rect 495 30 498 33 
rect 495 33 498 36 
rect 495 36 498 39 
rect 495 39 498 42 
rect 495 42 498 45 
rect 495 45 498 48 
rect 495 48 498 51 
rect 495 51 498 54 
rect 495 54 498 57 
rect 495 57 498 60 
rect 495 60 498 63 
rect 495 63 498 66 
rect 495 66 498 69 
rect 495 69 498 72 
rect 495 72 498 75 
rect 495 75 498 78 
rect 495 78 498 81 
rect 495 81 498 84 
rect 495 84 498 87 
rect 495 87 498 90 
rect 495 90 498 93 
rect 495 93 498 96 
rect 495 96 498 99 
rect 495 99 498 102 
rect 495 102 498 105 
rect 495 105 498 108 
rect 495 108 498 111 
rect 495 111 498 114 
rect 495 114 498 117 
rect 495 117 498 120 
rect 495 120 498 123 
rect 495 123 498 126 
rect 495 126 498 129 
rect 495 129 498 132 
rect 495 132 498 135 
rect 495 135 498 138 
rect 495 138 498 141 
rect 495 141 498 144 
rect 495 144 498 147 
rect 495 147 498 150 
rect 495 150 498 153 
rect 495 153 498 156 
rect 495 156 498 159 
rect 495 159 498 162 
rect 495 162 498 165 
rect 495 165 498 168 
rect 495 168 498 171 
rect 495 171 498 174 
rect 495 174 498 177 
rect 495 177 498 180 
rect 495 180 498 183 
rect 495 183 498 186 
rect 495 186 498 189 
rect 495 189 498 192 
rect 495 192 498 195 
rect 495 195 498 198 
rect 495 198 498 201 
rect 495 201 498 204 
rect 495 204 498 207 
rect 495 207 498 210 
rect 495 210 498 213 
rect 495 213 498 216 
rect 495 216 498 219 
rect 495 219 498 222 
rect 495 222 498 225 
rect 495 225 498 228 
rect 495 228 498 231 
rect 495 231 498 234 
rect 495 234 498 237 
rect 495 237 498 240 
rect 495 240 498 243 
rect 495 243 498 246 
rect 495 246 498 249 
rect 495 249 498 252 
rect 495 252 498 255 
rect 495 255 498 258 
rect 495 258 498 261 
rect 495 261 498 264 
rect 495 264 498 267 
rect 495 267 498 270 
rect 495 270 498 273 
rect 495 273 498 276 
rect 495 276 498 279 
rect 495 279 498 282 
rect 495 282 498 285 
rect 495 285 498 288 
rect 495 288 498 291 
rect 495 291 498 294 
rect 495 294 498 297 
rect 495 297 498 300 
rect 495 300 498 303 
rect 495 303 498 306 
rect 495 306 498 309 
rect 495 309 498 312 
rect 495 312 498 315 
rect 495 315 498 318 
rect 495 318 498 321 
rect 495 321 498 324 
rect 495 324 498 327 
rect 495 327 498 330 
rect 495 330 498 333 
rect 495 333 498 336 
rect 495 336 498 339 
rect 495 339 498 342 
rect 495 342 498 345 
rect 495 345 498 348 
rect 495 348 498 351 
rect 495 351 498 354 
rect 495 354 498 357 
rect 495 357 498 360 
rect 495 360 498 363 
rect 495 363 498 366 
rect 495 366 498 369 
rect 495 369 498 372 
rect 495 372 498 375 
rect 495 375 498 378 
rect 495 378 498 381 
rect 495 381 498 384 
rect 495 384 498 387 
rect 495 387 498 390 
rect 495 390 498 393 
rect 495 393 498 396 
rect 495 396 498 399 
rect 495 399 498 402 
rect 495 402 498 405 
rect 495 405 498 408 
rect 495 408 498 411 
rect 495 411 498 414 
rect 495 414 498 417 
rect 495 417 498 420 
rect 495 420 498 423 
rect 495 423 498 426 
rect 495 426 498 429 
rect 495 429 498 432 
rect 495 432 498 435 
rect 495 435 498 438 
rect 495 438 498 441 
rect 495 441 498 444 
rect 495 444 498 447 
rect 495 447 498 450 
rect 495 450 498 453 
rect 495 453 498 456 
rect 495 456 498 459 
rect 495 459 498 462 
rect 495 462 498 465 
rect 495 465 498 468 
rect 495 468 498 471 
rect 495 471 498 474 
rect 495 474 498 477 
rect 495 477 498 480 
rect 495 480 498 483 
rect 495 483 498 486 
rect 495 486 498 489 
rect 495 489 498 492 
rect 495 492 498 495 
rect 495 495 498 498 
rect 495 498 498 501 
rect 495 501 498 504 
rect 495 504 498 507 
rect 495 507 498 510 
rect 498 0 501 3 
rect 498 3 501 6 
rect 498 6 501 9 
rect 498 9 501 12 
rect 498 12 501 15 
rect 498 15 501 18 
rect 498 18 501 21 
rect 498 21 501 24 
rect 498 24 501 27 
rect 498 27 501 30 
rect 498 30 501 33 
rect 498 33 501 36 
rect 498 36 501 39 
rect 498 39 501 42 
rect 498 42 501 45 
rect 498 45 501 48 
rect 498 48 501 51 
rect 498 51 501 54 
rect 498 54 501 57 
rect 498 57 501 60 
rect 498 60 501 63 
rect 498 63 501 66 
rect 498 66 501 69 
rect 498 69 501 72 
rect 498 72 501 75 
rect 498 75 501 78 
rect 498 78 501 81 
rect 498 81 501 84 
rect 498 84 501 87 
rect 498 87 501 90 
rect 498 90 501 93 
rect 498 93 501 96 
rect 498 96 501 99 
rect 498 99 501 102 
rect 498 102 501 105 
rect 498 105 501 108 
rect 498 108 501 111 
rect 498 111 501 114 
rect 498 114 501 117 
rect 498 117 501 120 
rect 498 120 501 123 
rect 498 123 501 126 
rect 498 126 501 129 
rect 498 129 501 132 
rect 498 132 501 135 
rect 498 135 501 138 
rect 498 138 501 141 
rect 498 141 501 144 
rect 498 144 501 147 
rect 498 147 501 150 
rect 498 150 501 153 
rect 498 153 501 156 
rect 498 156 501 159 
rect 498 159 501 162 
rect 498 162 501 165 
rect 498 165 501 168 
rect 498 168 501 171 
rect 498 171 501 174 
rect 498 174 501 177 
rect 498 177 501 180 
rect 498 180 501 183 
rect 498 183 501 186 
rect 498 186 501 189 
rect 498 189 501 192 
rect 498 192 501 195 
rect 498 195 501 198 
rect 498 198 501 201 
rect 498 201 501 204 
rect 498 204 501 207 
rect 498 207 501 210 
rect 498 210 501 213 
rect 498 213 501 216 
rect 498 216 501 219 
rect 498 219 501 222 
rect 498 222 501 225 
rect 498 225 501 228 
rect 498 228 501 231 
rect 498 231 501 234 
rect 498 234 501 237 
rect 498 237 501 240 
rect 498 240 501 243 
rect 498 243 501 246 
rect 498 246 501 249 
rect 498 249 501 252 
rect 498 252 501 255 
rect 498 255 501 258 
rect 498 258 501 261 
rect 498 261 501 264 
rect 498 264 501 267 
rect 498 267 501 270 
rect 498 270 501 273 
rect 498 273 501 276 
rect 498 276 501 279 
rect 498 279 501 282 
rect 498 282 501 285 
rect 498 285 501 288 
rect 498 288 501 291 
rect 498 291 501 294 
rect 498 294 501 297 
rect 498 297 501 300 
rect 498 300 501 303 
rect 498 303 501 306 
rect 498 306 501 309 
rect 498 309 501 312 
rect 498 312 501 315 
rect 498 315 501 318 
rect 498 318 501 321 
rect 498 321 501 324 
rect 498 324 501 327 
rect 498 327 501 330 
rect 498 330 501 333 
rect 498 333 501 336 
rect 498 336 501 339 
rect 498 339 501 342 
rect 498 342 501 345 
rect 498 345 501 348 
rect 498 348 501 351 
rect 498 351 501 354 
rect 498 354 501 357 
rect 498 357 501 360 
rect 498 360 501 363 
rect 498 363 501 366 
rect 498 366 501 369 
rect 498 369 501 372 
rect 498 372 501 375 
rect 498 375 501 378 
rect 498 378 501 381 
rect 498 381 501 384 
rect 498 384 501 387 
rect 498 387 501 390 
rect 498 390 501 393 
rect 498 393 501 396 
rect 498 396 501 399 
rect 498 399 501 402 
rect 498 402 501 405 
rect 498 405 501 408 
rect 498 408 501 411 
rect 498 411 501 414 
rect 498 414 501 417 
rect 498 417 501 420 
rect 498 420 501 423 
rect 498 423 501 426 
rect 498 426 501 429 
rect 498 429 501 432 
rect 498 432 501 435 
rect 498 435 501 438 
rect 498 438 501 441 
rect 498 441 501 444 
rect 498 444 501 447 
rect 498 447 501 450 
rect 498 450 501 453 
rect 498 453 501 456 
rect 498 456 501 459 
rect 498 459 501 462 
rect 498 462 501 465 
rect 498 465 501 468 
rect 498 468 501 471 
rect 498 471 501 474 
rect 498 474 501 477 
rect 498 477 501 480 
rect 498 480 501 483 
rect 498 483 501 486 
rect 498 486 501 489 
rect 498 489 501 492 
rect 498 492 501 495 
rect 498 495 501 498 
rect 498 498 501 501 
rect 498 501 501 504 
rect 498 504 501 507 
rect 498 507 501 510 
rect 501 0 504 3 
rect 501 3 504 6 
rect 501 6 504 9 
rect 501 9 504 12 
rect 501 12 504 15 
rect 501 15 504 18 
rect 501 18 504 21 
rect 501 21 504 24 
rect 501 24 504 27 
rect 501 27 504 30 
rect 501 30 504 33 
rect 501 33 504 36 
rect 501 36 504 39 
rect 501 39 504 42 
rect 501 42 504 45 
rect 501 45 504 48 
rect 501 48 504 51 
rect 501 51 504 54 
rect 501 54 504 57 
rect 501 57 504 60 
rect 501 60 504 63 
rect 501 63 504 66 
rect 501 66 504 69 
rect 501 69 504 72 
rect 501 72 504 75 
rect 501 75 504 78 
rect 501 78 504 81 
rect 501 81 504 84 
rect 501 84 504 87 
rect 501 87 504 90 
rect 501 90 504 93 
rect 501 93 504 96 
rect 501 96 504 99 
rect 501 99 504 102 
rect 501 102 504 105 
rect 501 105 504 108 
rect 501 108 504 111 
rect 501 111 504 114 
rect 501 114 504 117 
rect 501 117 504 120 
rect 501 120 504 123 
rect 501 123 504 126 
rect 501 126 504 129 
rect 501 129 504 132 
rect 501 132 504 135 
rect 501 135 504 138 
rect 501 138 504 141 
rect 501 141 504 144 
rect 501 144 504 147 
rect 501 147 504 150 
rect 501 150 504 153 
rect 501 153 504 156 
rect 501 156 504 159 
rect 501 159 504 162 
rect 501 162 504 165 
rect 501 165 504 168 
rect 501 168 504 171 
rect 501 171 504 174 
rect 501 174 504 177 
rect 501 177 504 180 
rect 501 180 504 183 
rect 501 183 504 186 
rect 501 186 504 189 
rect 501 189 504 192 
rect 501 192 504 195 
rect 501 195 504 198 
rect 501 198 504 201 
rect 501 201 504 204 
rect 501 204 504 207 
rect 501 207 504 210 
rect 501 210 504 213 
rect 501 213 504 216 
rect 501 216 504 219 
rect 501 219 504 222 
rect 501 222 504 225 
rect 501 225 504 228 
rect 501 228 504 231 
rect 501 231 504 234 
rect 501 234 504 237 
rect 501 237 504 240 
rect 501 240 504 243 
rect 501 243 504 246 
rect 501 246 504 249 
rect 501 249 504 252 
rect 501 252 504 255 
rect 501 255 504 258 
rect 501 258 504 261 
rect 501 261 504 264 
rect 501 264 504 267 
rect 501 267 504 270 
rect 501 270 504 273 
rect 501 273 504 276 
rect 501 276 504 279 
rect 501 279 504 282 
rect 501 282 504 285 
rect 501 285 504 288 
rect 501 288 504 291 
rect 501 291 504 294 
rect 501 294 504 297 
rect 501 297 504 300 
rect 501 300 504 303 
rect 501 303 504 306 
rect 501 306 504 309 
rect 501 309 504 312 
rect 501 312 504 315 
rect 501 315 504 318 
rect 501 318 504 321 
rect 501 321 504 324 
rect 501 324 504 327 
rect 501 327 504 330 
rect 501 330 504 333 
rect 501 333 504 336 
rect 501 336 504 339 
rect 501 339 504 342 
rect 501 342 504 345 
rect 501 345 504 348 
rect 501 348 504 351 
rect 501 351 504 354 
rect 501 354 504 357 
rect 501 357 504 360 
rect 501 360 504 363 
rect 501 363 504 366 
rect 501 366 504 369 
rect 501 369 504 372 
rect 501 372 504 375 
rect 501 375 504 378 
rect 501 378 504 381 
rect 501 381 504 384 
rect 501 384 504 387 
rect 501 387 504 390 
rect 501 390 504 393 
rect 501 393 504 396 
rect 501 396 504 399 
rect 501 399 504 402 
rect 501 402 504 405 
rect 501 405 504 408 
rect 501 408 504 411 
rect 501 411 504 414 
rect 501 414 504 417 
rect 501 417 504 420 
rect 501 420 504 423 
rect 501 423 504 426 
rect 501 426 504 429 
rect 501 429 504 432 
rect 501 432 504 435 
rect 501 435 504 438 
rect 501 438 504 441 
rect 501 441 504 444 
rect 501 444 504 447 
rect 501 447 504 450 
rect 501 450 504 453 
rect 501 453 504 456 
rect 501 456 504 459 
rect 501 459 504 462 
rect 501 462 504 465 
rect 501 465 504 468 
rect 501 468 504 471 
rect 501 471 504 474 
rect 501 474 504 477 
rect 501 477 504 480 
rect 501 480 504 483 
rect 501 483 504 486 
rect 501 486 504 489 
rect 501 489 504 492 
rect 501 492 504 495 
rect 501 495 504 498 
rect 501 498 504 501 
rect 501 501 504 504 
rect 501 504 504 507 
rect 501 507 504 510 
rect 504 0 507 3 
rect 504 3 507 6 
rect 504 6 507 9 
rect 504 9 507 12 
rect 504 12 507 15 
rect 504 15 507 18 
rect 504 18 507 21 
rect 504 21 507 24 
rect 504 24 507 27 
rect 504 27 507 30 
rect 504 30 507 33 
rect 504 33 507 36 
rect 504 36 507 39 
rect 504 39 507 42 
rect 504 42 507 45 
rect 504 45 507 48 
rect 504 48 507 51 
rect 504 51 507 54 
rect 504 54 507 57 
rect 504 57 507 60 
rect 504 60 507 63 
rect 504 63 507 66 
rect 504 66 507 69 
rect 504 69 507 72 
rect 504 72 507 75 
rect 504 75 507 78 
rect 504 78 507 81 
rect 504 81 507 84 
rect 504 84 507 87 
rect 504 87 507 90 
rect 504 90 507 93 
rect 504 93 507 96 
rect 504 96 507 99 
rect 504 99 507 102 
rect 504 102 507 105 
rect 504 105 507 108 
rect 504 108 507 111 
rect 504 111 507 114 
rect 504 114 507 117 
rect 504 117 507 120 
rect 504 120 507 123 
rect 504 123 507 126 
rect 504 126 507 129 
rect 504 129 507 132 
rect 504 132 507 135 
rect 504 135 507 138 
rect 504 138 507 141 
rect 504 141 507 144 
rect 504 144 507 147 
rect 504 147 507 150 
rect 504 150 507 153 
rect 504 153 507 156 
rect 504 156 507 159 
rect 504 159 507 162 
rect 504 162 507 165 
rect 504 165 507 168 
rect 504 168 507 171 
rect 504 171 507 174 
rect 504 174 507 177 
rect 504 177 507 180 
rect 504 180 507 183 
rect 504 183 507 186 
rect 504 186 507 189 
rect 504 189 507 192 
rect 504 192 507 195 
rect 504 195 507 198 
rect 504 198 507 201 
rect 504 201 507 204 
rect 504 204 507 207 
rect 504 207 507 210 
rect 504 210 507 213 
rect 504 213 507 216 
rect 504 216 507 219 
rect 504 219 507 222 
rect 504 222 507 225 
rect 504 225 507 228 
rect 504 228 507 231 
rect 504 231 507 234 
rect 504 234 507 237 
rect 504 237 507 240 
rect 504 240 507 243 
rect 504 243 507 246 
rect 504 246 507 249 
rect 504 249 507 252 
rect 504 252 507 255 
rect 504 255 507 258 
rect 504 258 507 261 
rect 504 261 507 264 
rect 504 264 507 267 
rect 504 267 507 270 
rect 504 270 507 273 
rect 504 273 507 276 
rect 504 276 507 279 
rect 504 279 507 282 
rect 504 282 507 285 
rect 504 285 507 288 
rect 504 288 507 291 
rect 504 291 507 294 
rect 504 294 507 297 
rect 504 297 507 300 
rect 504 300 507 303 
rect 504 303 507 306 
rect 504 306 507 309 
rect 504 309 507 312 
rect 504 312 507 315 
rect 504 315 507 318 
rect 504 318 507 321 
rect 504 321 507 324 
rect 504 324 507 327 
rect 504 327 507 330 
rect 504 330 507 333 
rect 504 333 507 336 
rect 504 336 507 339 
rect 504 339 507 342 
rect 504 342 507 345 
rect 504 345 507 348 
rect 504 348 507 351 
rect 504 351 507 354 
rect 504 354 507 357 
rect 504 357 507 360 
rect 504 360 507 363 
rect 504 363 507 366 
rect 504 366 507 369 
rect 504 369 507 372 
rect 504 372 507 375 
rect 504 375 507 378 
rect 504 378 507 381 
rect 504 381 507 384 
rect 504 384 507 387 
rect 504 387 507 390 
rect 504 390 507 393 
rect 504 393 507 396 
rect 504 396 507 399 
rect 504 399 507 402 
rect 504 402 507 405 
rect 504 405 507 408 
rect 504 408 507 411 
rect 504 411 507 414 
rect 504 414 507 417 
rect 504 417 507 420 
rect 504 420 507 423 
rect 504 423 507 426 
rect 504 426 507 429 
rect 504 429 507 432 
rect 504 432 507 435 
rect 504 435 507 438 
rect 504 438 507 441 
rect 504 441 507 444 
rect 504 444 507 447 
rect 504 447 507 450 
rect 504 450 507 453 
rect 504 453 507 456 
rect 504 456 507 459 
rect 504 459 507 462 
rect 504 462 507 465 
rect 504 465 507 468 
rect 504 468 507 471 
rect 504 471 507 474 
rect 504 474 507 477 
rect 504 477 507 480 
rect 504 480 507 483 
rect 504 483 507 486 
rect 504 486 507 489 
rect 504 489 507 492 
rect 504 492 507 495 
rect 504 495 507 498 
rect 504 498 507 501 
rect 504 501 507 504 
rect 504 504 507 507 
rect 504 507 507 510 
rect 507 0 510 3 
rect 507 3 510 6 
rect 507 6 510 9 
rect 507 9 510 12 
rect 507 12 510 15 
rect 507 15 510 18 
rect 507 18 510 21 
rect 507 21 510 24 
rect 507 24 510 27 
rect 507 27 510 30 
rect 507 30 510 33 
rect 507 33 510 36 
rect 507 36 510 39 
rect 507 39 510 42 
rect 507 42 510 45 
rect 507 45 510 48 
rect 507 48 510 51 
rect 507 51 510 54 
rect 507 54 510 57 
rect 507 57 510 60 
rect 507 60 510 63 
rect 507 63 510 66 
rect 507 66 510 69 
rect 507 69 510 72 
rect 507 72 510 75 
rect 507 75 510 78 
rect 507 78 510 81 
rect 507 81 510 84 
rect 507 84 510 87 
rect 507 87 510 90 
rect 507 90 510 93 
rect 507 93 510 96 
rect 507 96 510 99 
rect 507 99 510 102 
rect 507 102 510 105 
rect 507 105 510 108 
rect 507 108 510 111 
rect 507 111 510 114 
rect 507 114 510 117 
rect 507 117 510 120 
rect 507 120 510 123 
rect 507 123 510 126 
rect 507 126 510 129 
rect 507 129 510 132 
rect 507 132 510 135 
rect 507 135 510 138 
rect 507 138 510 141 
rect 507 141 510 144 
rect 507 144 510 147 
rect 507 147 510 150 
rect 507 150 510 153 
rect 507 153 510 156 
rect 507 156 510 159 
rect 507 159 510 162 
rect 507 162 510 165 
rect 507 165 510 168 
rect 507 168 510 171 
rect 507 171 510 174 
rect 507 174 510 177 
rect 507 177 510 180 
rect 507 180 510 183 
rect 507 183 510 186 
rect 507 186 510 189 
rect 507 189 510 192 
rect 507 192 510 195 
rect 507 195 510 198 
rect 507 198 510 201 
rect 507 201 510 204 
rect 507 204 510 207 
rect 507 207 510 210 
rect 507 210 510 213 
rect 507 213 510 216 
rect 507 216 510 219 
rect 507 219 510 222 
rect 507 222 510 225 
rect 507 225 510 228 
rect 507 228 510 231 
rect 507 231 510 234 
rect 507 234 510 237 
rect 507 237 510 240 
rect 507 240 510 243 
rect 507 243 510 246 
rect 507 246 510 249 
rect 507 249 510 252 
rect 507 252 510 255 
rect 507 255 510 258 
rect 507 258 510 261 
rect 507 261 510 264 
rect 507 264 510 267 
rect 507 267 510 270 
rect 507 270 510 273 
rect 507 273 510 276 
rect 507 276 510 279 
rect 507 279 510 282 
rect 507 282 510 285 
rect 507 285 510 288 
rect 507 288 510 291 
rect 507 291 510 294 
rect 507 294 510 297 
rect 507 297 510 300 
rect 507 300 510 303 
rect 507 303 510 306 
rect 507 306 510 309 
rect 507 309 510 312 
rect 507 312 510 315 
rect 507 315 510 318 
rect 507 318 510 321 
rect 507 321 510 324 
rect 507 324 510 327 
rect 507 327 510 330 
rect 507 330 510 333 
rect 507 333 510 336 
rect 507 336 510 339 
rect 507 339 510 342 
rect 507 342 510 345 
rect 507 345 510 348 
rect 507 348 510 351 
rect 507 351 510 354 
rect 507 354 510 357 
rect 507 357 510 360 
rect 507 360 510 363 
rect 507 363 510 366 
rect 507 366 510 369 
rect 507 369 510 372 
rect 507 372 510 375 
rect 507 375 510 378 
rect 507 378 510 381 
rect 507 381 510 384 
rect 507 384 510 387 
rect 507 387 510 390 
rect 507 390 510 393 
rect 507 393 510 396 
rect 507 396 510 399 
rect 507 399 510 402 
rect 507 402 510 405 
rect 507 405 510 408 
rect 507 408 510 411 
rect 507 411 510 414 
rect 507 414 510 417 
rect 507 417 510 420 
rect 507 420 510 423 
rect 507 423 510 426 
rect 507 426 510 429 
rect 507 429 510 432 
rect 507 432 510 435 
rect 507 435 510 438 
rect 507 438 510 441 
rect 507 441 510 444 
rect 507 444 510 447 
rect 507 447 510 450 
rect 507 450 510 453 
rect 507 453 510 456 
rect 507 456 510 459 
rect 507 459 510 462 
rect 507 462 510 465 
rect 507 465 510 468 
rect 507 468 510 471 
rect 507 471 510 474 
rect 507 474 510 477 
rect 507 477 510 480 
rect 507 480 510 483 
rect 507 483 510 486 
rect 507 486 510 489 
rect 507 489 510 492 
rect 507 492 510 495 
rect 507 495 510 498 
rect 507 498 510 501 
rect 507 501 510 504 
rect 507 504 510 507 
rect 507 507 510 510 
<< end >>
3.99seconds.
